
module rx_DW01_add_10_1 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;
  assign \carry[1]  = A[0];

  FA1A U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(\carry[3] )
         );
  FA1A U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(\carry[4] )
         );
  FA1A U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(\carry[5] )
         );
  FA1A U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(\carry[6] )
         );
  FA1A U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(\carry[7] )
         );
  FA1A U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(\carry[8] )
         );
  FA1A U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(\carry[9] )
         );
  FA1A U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(\carry[2] )
         );
  EO3P U1_9 ( .A(A[9]), .B(B[9]), .C(\carry[9] ), .Z(SUM[9]) );
endmodule


module rx_DW01_add_10_0 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  FA1A U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(\carry[2] )
         );
  FA1A U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(\carry[3] )
         );
  FA1A U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(\carry[4] )
         );
  FA1A U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(\carry[5] )
         );
  FA1A U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(\carry[6] )
         );
  FA1A U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(\carry[7] )
         );
  FA1A U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(\carry[8] )
         );
  FA1A U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(\carry[9] )
         );
  EO3P U1_9 ( .A(A[9]), .B(B[9]), .C(\carry[9] ), .Z(SUM[9]) );
  AN2 U4 ( .A(B[0]), .B(A[0]), .Z(\carry[1] ) );
  EO U5 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
endmodule


module rx ( sum_0, dec_tap_1, sum_1 );
  input [9:0] sum_0;
  input [9:0] dec_tap_1;
  output [9:0] sum_1;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sum_1[0] = 1'b0;

  rx_DW01_add_10_1 add_0_root_add_10_3 ( .A({N9, N8, N7, N6, N5, N4, N3, N2, 
        N1, N0}), .B({N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), .CI(1'b0), 
        .SUM({sum_1[9:1], SYNOPSYS_UNCONNECTED__0}) );
  rx_DW01_add_10_0 r260 ( .A(sum_0), .B(dec_tap_1), .CI(1'b0), .SUM({N9, N8, 
        N7, N6, N5, N4, N3, N2, N1, N0}) );
endmodule


module tx_DW_mult_uns_1 ( a, b, product );
  input [63:0] a;
  input [63:0] b;
  output [127:0] product;
  wire   n1, n2, n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n50, n60, n70, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n877, n878, n879, n880,
         n882, n883, n884, n885, n886, n888, n889, n890, n891, n892, n894,
         n895, n896, n897, n898, n900, n901, n902, n903, n904, n906, n907,
         n908, n909, n910, n912, n913, n914, n915, n916, n918, n919, n920,
         n921, n922, n924, n925, n926, n927, n928, n930, n931, n932, n933,
         n934, n936, n937, n938, n939, n940, n942, n943, n944, n945, n946,
         n948, n949, n950, n951, n952, n954, n955, n956, n957, n958, n960,
         n961, n962, n963, n964, n966, n967, n968, n969, n970, n972, n973,
         n974, n975, n976, n978, n979, n980, n981, n982, n984, n985, n986,
         n987, n988, n990, n991, n992, n993, n994, n996, n997, n998, n999,
         n1000, n1002, n1003, n1004, n1005, n1006, n1008, n1009, n1010, n1011,
         n1012, n1014, n1015, n1016, n1017, n1018, n1020, n1021, n1022, n1023,
         n1024, n1026, n1027, n1028, n1029, n1030, n1032, n1033, n1034, n1035,
         n1036, n1038, n1039, n1040, n1041, n1042, n1044, n1045, n1046, n1047,
         n1048, n1050, n1051, n1052, n1053, n1054, n1056, n1057, n1058, n1059,
         n1060, n1062, n1063, n1064, n1065, n1066, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897;

  IV U1 ( .A(n10251), .Z(n1068) );
  ND2 OR_NOTi ( .A(n1068), .B(n10733), .Z(n1519) );
  IV U11 ( .A(n10573), .Z(n1066) );
  IV U3 ( .A(n1390), .Z(n1065) );
  IV U21 ( .A(n10573), .Z(n1064) );
  IV U12 ( .A(n10409), .Z(n1063) );
  AO7 AO21i ( .A(n1063), .B(n1064), .C(n1065), .Z(n3727) );
  IV U13 ( .A(n10251), .Z(n1062) );
  ND2 OR_NOTi1 ( .A(n1062), .B(n10728), .Z(n1584) );
  IV U14 ( .A(n10568), .Z(n1060) );
  IV U31 ( .A(n1391), .Z(n1059) );
  IV U23 ( .A(n10568), .Z(n1058) );
  IV U15 ( .A(n10404), .Z(n1057) );
  AO7 AO21i1 ( .A(n1057), .B(n1058), .C(n1059), .Z(n3793) );
  IV U16 ( .A(n10251), .Z(n1056) );
  ND2 OR_NOTi2 ( .A(n1056), .B(n10723), .Z(n1649) );
  IV U17 ( .A(n10563), .Z(n1054) );
  IV U32 ( .A(n1392), .Z(n1053) );
  IV U25 ( .A(n10563), .Z(n1052) );
  IV U18 ( .A(n10399), .Z(n1051) );
  AO7 AO21i2 ( .A(n1051), .B(n1052), .C(n1053), .Z(n3859) );
  IV U19 ( .A(n10251), .Z(n1050) );
  ND2 OR_NOTi3 ( .A(n1050), .B(n10718), .Z(n1714) );
  IV U110 ( .A(n10558), .Z(n1048) );
  IV U33 ( .A(n1393), .Z(n1047) );
  IV U27 ( .A(n10558), .Z(n1046) );
  IV U111 ( .A(n10394), .Z(n1045) );
  AO7 AO21i3 ( .A(n1045), .B(n1046), .C(n1047), .Z(n3925) );
  IV U112 ( .A(n10251), .Z(n1044) );
  ND2 OR_NOTi4 ( .A(n1044), .B(n10713), .Z(n1779) );
  IV U113 ( .A(n10553), .Z(n1042) );
  IV U34 ( .A(n1394), .Z(n1041) );
  IV U29 ( .A(n10553), .Z(n1040) );
  IV U114 ( .A(n10389), .Z(n1039) );
  AO7 AO21i4 ( .A(n1039), .B(n1040), .C(n1041), .Z(n3991) );
  IV U115 ( .A(n10250), .Z(n1038) );
  ND2 OR_NOTi5 ( .A(n1038), .B(n10708), .Z(n1844) );
  IV U116 ( .A(n10548), .Z(n1036) );
  IV U35 ( .A(n1395), .Z(n1035) );
  IV U211 ( .A(n10548), .Z(n1034) );
  IV U117 ( .A(n10384), .Z(n1033) );
  AO7 AO21i5 ( .A(n1033), .B(n1034), .C(n1035), .Z(n4057) );
  IV U118 ( .A(n10250), .Z(n1032) );
  ND2 OR_NOTi6 ( .A(n1032), .B(n10703), .Z(n1909) );
  IV U119 ( .A(n10543), .Z(n1030) );
  IV U36 ( .A(n1396), .Z(n1029) );
  IV U213 ( .A(n10543), .Z(n1028) );
  IV U120 ( .A(n10379), .Z(n1027) );
  AO7 AO21i6 ( .A(n1027), .B(n1028), .C(n1029), .Z(n4123) );
  IV U121 ( .A(n10250), .Z(n1026) );
  ND2 OR_NOTi7 ( .A(n1026), .B(n10698), .Z(n1974) );
  IV U122 ( .A(n10538), .Z(n1024) );
  IV U37 ( .A(n1397), .Z(n1023) );
  IV U215 ( .A(n10538), .Z(n1022) );
  IV U123 ( .A(n10374), .Z(n1021) );
  AO7 AO21i7 ( .A(n1021), .B(n1022), .C(n1023), .Z(n4189) );
  IV U124 ( .A(n10250), .Z(n1020) );
  ND2 OR_NOTi8 ( .A(n1020), .B(n10693), .Z(n2039) );
  IV U125 ( .A(n10533), .Z(n1018) );
  IV U38 ( .A(n1398), .Z(n1017) );
  IV U217 ( .A(n10533), .Z(n1016) );
  IV U126 ( .A(n10369), .Z(n1015) );
  AO7 AO21i8 ( .A(n1015), .B(n1016), .C(n1017), .Z(n4255) );
  IV U127 ( .A(n10250), .Z(n1014) );
  ND2 OR_NOTi9 ( .A(n1014), .B(n10688), .Z(n2104) );
  IV U128 ( .A(n10528), .Z(n1012) );
  IV U39 ( .A(n1399), .Z(n1011) );
  IV U219 ( .A(n10528), .Z(n1010) );
  IV U129 ( .A(n10364), .Z(n1009) );
  AO7 AO21i9 ( .A(n1009), .B(n1010), .C(n1011), .Z(n4321) );
  IV U130 ( .A(n10250), .Z(n1008) );
  ND2 OR_NOTi10 ( .A(n1008), .B(n10683), .Z(n2169) );
  IV U131 ( .A(n10523), .Z(n1006) );
  IV U310 ( .A(n1400), .Z(n1005) );
  IV U221 ( .A(n10523), .Z(n1004) );
  IV U132 ( .A(n10359), .Z(n1003) );
  AO7 AO21i10 ( .A(n1003), .B(n1004), .C(n1005), .Z(n4387) );
  IV U133 ( .A(n10250), .Z(n1002) );
  ND2 OR_NOTi11 ( .A(n1002), .B(n10678), .Z(n2234) );
  IV U134 ( .A(n10518), .Z(n1000) );
  IV U311 ( .A(n1401), .Z(n999) );
  IV U223 ( .A(n10518), .Z(n998) );
  IV U135 ( .A(n10354), .Z(n997) );
  AO7 AO21i11 ( .A(n997), .B(n998), .C(n999), .Z(n4453) );
  IV U136 ( .A(n10249), .Z(n996) );
  ND2 OR_NOTi12 ( .A(n996), .B(n10673), .Z(n2299) );
  IV U137 ( .A(n10513), .Z(n994) );
  IV U312 ( .A(n1402), .Z(n993) );
  IV U225 ( .A(n10513), .Z(n992) );
  IV U138 ( .A(n10349), .Z(n991) );
  AO7 AO21i12 ( .A(n991), .B(n992), .C(n993), .Z(n4519) );
  IV U139 ( .A(n10249), .Z(n990) );
  ND2 OR_NOTi13 ( .A(n990), .B(n10668), .Z(n2364) );
  IV U140 ( .A(n10508), .Z(n988) );
  IV U313 ( .A(n1403), .Z(n987) );
  IV U227 ( .A(n10508), .Z(n986) );
  IV U141 ( .A(n10344), .Z(n985) );
  AO7 AO21i13 ( .A(n985), .B(n986), .C(n987), .Z(n4585) );
  IV U142 ( .A(n10249), .Z(n984) );
  ND2 OR_NOTi14 ( .A(n984), .B(n10663), .Z(n2429) );
  IV U143 ( .A(n10503), .Z(n982) );
  IV U314 ( .A(n1404), .Z(n981) );
  IV U229 ( .A(n10503), .Z(n980) );
  IV U144 ( .A(n10339), .Z(n979) );
  AO7 AO21i14 ( .A(n979), .B(n980), .C(n981), .Z(n4651) );
  IV U145 ( .A(n10249), .Z(n978) );
  ND2 OR_NOTi15 ( .A(n978), .B(n10658), .Z(n2494) );
  IV U146 ( .A(n10498), .Z(n976) );
  IV U315 ( .A(n1405), .Z(n975) );
  IV U231 ( .A(n10498), .Z(n974) );
  IV U147 ( .A(n10334), .Z(n973) );
  AO7 AO21i15 ( .A(n973), .B(n974), .C(n975), .Z(n4717) );
  IV U148 ( .A(n10249), .Z(n972) );
  ND2 OR_NOTi16 ( .A(n972), .B(n10653), .Z(n2559) );
  IV U149 ( .A(n10493), .Z(n970) );
  IV U316 ( .A(n1406), .Z(n969) );
  IV U233 ( .A(n10493), .Z(n968) );
  IV U150 ( .A(n10329), .Z(n967) );
  AO7 AO21i16 ( .A(n967), .B(n968), .C(n969), .Z(n4783) );
  IV U151 ( .A(n10249), .Z(n966) );
  ND2 OR_NOTi17 ( .A(n966), .B(n10648), .Z(n2624) );
  IV U152 ( .A(n10488), .Z(n964) );
  IV U317 ( .A(n1407), .Z(n963) );
  IV U235 ( .A(n10488), .Z(n962) );
  IV U153 ( .A(n10324), .Z(n961) );
  AO7 AO21i17 ( .A(n961), .B(n962), .C(n963), .Z(n4849) );
  IV U154 ( .A(n10249), .Z(n960) );
  ND2 OR_NOTi18 ( .A(n960), .B(n10643), .Z(n2689) );
  IV U155 ( .A(n10483), .Z(n958) );
  IV U318 ( .A(n1408), .Z(n957) );
  IV U237 ( .A(n10483), .Z(n956) );
  IV U156 ( .A(n10319), .Z(n955) );
  AO7 AO21i18 ( .A(n955), .B(n956), .C(n957), .Z(n4915) );
  IV U157 ( .A(n10248), .Z(n954) );
  ND2 OR_NOTi19 ( .A(n954), .B(n10638), .Z(n2754) );
  IV U158 ( .A(n10478), .Z(n952) );
  IV U319 ( .A(n1409), .Z(n951) );
  IV U239 ( .A(n10478), .Z(n950) );
  IV U159 ( .A(n10314), .Z(n949) );
  AO7 AO21i19 ( .A(n949), .B(n950), .C(n951), .Z(n4981) );
  IV U160 ( .A(n10248), .Z(n948) );
  ND2 OR_NOTi20 ( .A(n948), .B(n10633), .Z(n2819) );
  IV U161 ( .A(n10473), .Z(n946) );
  IV U320 ( .A(n1410), .Z(n945) );
  IV U241 ( .A(n10473), .Z(n944) );
  IV U162 ( .A(n10309), .Z(n943) );
  AO7 AO21i20 ( .A(n943), .B(n944), .C(n945), .Z(n5047) );
  IV U163 ( .A(n10248), .Z(n942) );
  ND2 OR_NOTi21 ( .A(n942), .B(n10628), .Z(n2884) );
  IV U164 ( .A(n10468), .Z(n940) );
  IV U321 ( .A(n1411), .Z(n939) );
  IV U243 ( .A(n10468), .Z(n938) );
  IV U165 ( .A(n10304), .Z(n937) );
  AO7 AO21i21 ( .A(n937), .B(n938), .C(n939), .Z(n5113) );
  IV U166 ( .A(n10248), .Z(n936) );
  ND2 OR_NOTi22 ( .A(n936), .B(n10623), .Z(n2949) );
  IV U167 ( .A(n10463), .Z(n934) );
  IV U322 ( .A(n1412), .Z(n933) );
  IV U245 ( .A(n10463), .Z(n932) );
  IV U168 ( .A(n10299), .Z(n931) );
  AO7 AO21i22 ( .A(n931), .B(n932), .C(n933), .Z(n5179) );
  IV U169 ( .A(n10248), .Z(n930) );
  ND2 OR_NOTi23 ( .A(n930), .B(n10618), .Z(n3014) );
  IV U170 ( .A(n10458), .Z(n928) );
  IV U323 ( .A(n1413), .Z(n927) );
  IV U247 ( .A(n10458), .Z(n926) );
  IV U171 ( .A(n10294), .Z(n925) );
  AO7 AO21i23 ( .A(n925), .B(n926), .C(n927), .Z(n5245) );
  IV U172 ( .A(n10248), .Z(n924) );
  ND2 OR_NOTi24 ( .A(n924), .B(n10613), .Z(n3079) );
  IV U173 ( .A(n10453), .Z(n922) );
  IV U324 ( .A(n1414), .Z(n921) );
  IV U249 ( .A(n10453), .Z(n920) );
  IV U174 ( .A(n10289), .Z(n919) );
  AO7 AO21i24 ( .A(n919), .B(n920), .C(n921), .Z(n5311) );
  IV U175 ( .A(n10248), .Z(n918) );
  ND2 OR_NOTi25 ( .A(n918), .B(n10608), .Z(n3144) );
  IV U176 ( .A(n10448), .Z(n916) );
  IV U325 ( .A(n1415), .Z(n915) );
  IV U251 ( .A(n10448), .Z(n914) );
  IV U177 ( .A(n10284), .Z(n913) );
  AO7 AO21i25 ( .A(n913), .B(n914), .C(n915), .Z(n5377) );
  IV U178 ( .A(n10247), .Z(n912) );
  ND2 OR_NOTi26 ( .A(n912), .B(n10603), .Z(n3209) );
  IV U179 ( .A(n10443), .Z(n910) );
  IV U326 ( .A(n1416), .Z(n909) );
  IV U253 ( .A(n10443), .Z(n908) );
  IV U180 ( .A(n10279), .Z(n907) );
  AO7 AO21i26 ( .A(n907), .B(n908), .C(n909), .Z(n5443) );
  IV U181 ( .A(n10247), .Z(n906) );
  ND2 OR_NOTi27 ( .A(n906), .B(n10598), .Z(n3274) );
  IV U182 ( .A(n10438), .Z(n904) );
  IV U327 ( .A(n1417), .Z(n903) );
  IV U255 ( .A(n10438), .Z(n902) );
  IV U183 ( .A(n10274), .Z(n901) );
  AO7 AO21i27 ( .A(n901), .B(n902), .C(n903), .Z(n5509) );
  IV U184 ( .A(n10247), .Z(n900) );
  ND2 OR_NOTi28 ( .A(n900), .B(n10593), .Z(n3339) );
  IV U185 ( .A(n10433), .Z(n898) );
  IV U328 ( .A(n1418), .Z(n897) );
  IV U257 ( .A(n10433), .Z(n896) );
  IV U186 ( .A(n10269), .Z(n895) );
  AO7 AO21i28 ( .A(n895), .B(n896), .C(n897), .Z(n5575) );
  IV U187 ( .A(n10247), .Z(n894) );
  ND2 OR_NOTi29 ( .A(n894), .B(n10588), .Z(n3404) );
  IV U188 ( .A(n10428), .Z(n892) );
  IV U329 ( .A(n1419), .Z(n891) );
  IV U259 ( .A(n10428), .Z(n890) );
  IV U189 ( .A(n10264), .Z(n889) );
  AO7 AO21i29 ( .A(n889), .B(n890), .C(n891), .Z(n5641) );
  IV U190 ( .A(n10247), .Z(n888) );
  ND2 OR_NOTi30 ( .A(n888), .B(n10583), .Z(n3469) );
  IV U191 ( .A(n10423), .Z(n886) );
  IV U330 ( .A(n1420), .Z(n885) );
  IV U261 ( .A(n10423), .Z(n884) );
  IV U192 ( .A(n10259), .Z(n883) );
  AO7 AO21i30 ( .A(n883), .B(n884), .C(n885), .Z(n5707) );
  IV U193 ( .A(n10247), .Z(n882) );
  ND2 OR_NOTi31 ( .A(n882), .B(n10578), .Z(n3534) );
  IV U194 ( .A(n10418), .Z(n880) );
  IV U331 ( .A(n1421), .Z(n879) );
  IV U263 ( .A(n10418), .Z(n878) );
  IV U195 ( .A(n10254), .Z(n877) );
  AO7 AO21i31 ( .A(n877), .B(n878), .C(n879), .Z(n5773) );
  IV U196 ( .A(n10414), .Z(n875) );
  IVP U4 ( .A(n1358), .Z(n1) );
  IVP U6 ( .A(n1358), .Z(n2) );
  IVP U8 ( .A(n1358), .Z(n3) );
  IVP U10 ( .A(n1358), .Z(n8) );
  IVP U30 ( .A(n1358), .Z(n9) );
  IVP U41 ( .A(n1359), .Z(n10) );
  IVP U43 ( .A(n1359), .Z(n11) );
  IVP U45 ( .A(n1359), .Z(n12) );
  IVP U47 ( .A(n1359), .Z(n13) );
  IVP U49 ( .A(n1359), .Z(n14) );
  IVP U51 ( .A(n1360), .Z(n15) );
  IVP U53 ( .A(n1360), .Z(n16) );
  IVP U55 ( .A(n1360), .Z(n17) );
  IVP U57 ( .A(n1360), .Z(n18) );
  IVP U59 ( .A(n1360), .Z(n19) );
  IVP U61 ( .A(n1361), .Z(n20) );
  IVP U63 ( .A(n1361), .Z(n21) );
  IVP U65 ( .A(n1361), .Z(n22) );
  IVP U67 ( .A(n1361), .Z(n23) );
  IVP U69 ( .A(n1361), .Z(n24) );
  IVP U71 ( .A(n1362), .Z(n25) );
  IVP U73 ( .A(n1362), .Z(n26) );
  IVP U75 ( .A(n1362), .Z(n27) );
  IVP U77 ( .A(n1362), .Z(n28) );
  IVP U79 ( .A(n1362), .Z(n29) );
  IVP U81 ( .A(n1363), .Z(n30) );
  IVP U83 ( .A(n1363), .Z(n31) );
  IVP U85 ( .A(n1363), .Z(n32) );
  IVP U87 ( .A(n1363), .Z(n33) );
  IVP U89 ( .A(n1363), .Z(n34) );
  IVP U91 ( .A(n1364), .Z(n35) );
  IVP U93 ( .A(n1364), .Z(n36) );
  IVP U95 ( .A(n1364), .Z(n37) );
  IVP U97 ( .A(n1364), .Z(n38) );
  IVP U99 ( .A(n1364), .Z(n39) );
  IVP U101 ( .A(n1365), .Z(n40) );
  IVP U103 ( .A(n1365), .Z(n50) );
  IVP U105 ( .A(n1365), .Z(n60) );
  IVP U107 ( .A(n1365), .Z(n70) );
  IVP U109 ( .A(n1365), .Z(n80) );
  IVP U198 ( .A(n1366), .Z(n81) );
  IVP U200 ( .A(n1366), .Z(n82) );
  IVP U202 ( .A(n1366), .Z(n83) );
  IVP U204 ( .A(n1366), .Z(n84) );
  IVP U206 ( .A(n1366), .Z(n85) );
  IVP U208 ( .A(n1367), .Z(n86) );
  IVP U265 ( .A(n1367), .Z(n87) );
  IVP U267 ( .A(n1367), .Z(n88) );
  IVP U269 ( .A(n1367), .Z(n89) );
  IVP U271 ( .A(n1367), .Z(n90) );
  IVP U273 ( .A(n1368), .Z(n91) );
  IVP U275 ( .A(n1368), .Z(n92) );
  IVP U277 ( .A(n1368), .Z(n93) );
  IVP U279 ( .A(n1368), .Z(n94) );
  IVP U281 ( .A(n1368), .Z(n95) );
  IVP U283 ( .A(n1369), .Z(n96) );
  IVP U285 ( .A(n1369), .Z(n97) );
  IVP U287 ( .A(n1369), .Z(n98) );
  IVP U289 ( .A(n1369), .Z(n99) );
  IVP U291 ( .A(n1369), .Z(n100) );
  IVP U293 ( .A(n1370), .Z(n101) );
  IVP U295 ( .A(n1370), .Z(n102) );
  IVP U297 ( .A(n1370), .Z(n103) );
  IVP U299 ( .A(n1370), .Z(n104) );
  IVP U301 ( .A(n1370), .Z(n105) );
  IVP U303 ( .A(n1371), .Z(n106) );
  IVP U305 ( .A(n1371), .Z(n107) );
  IVP U307 ( .A(n1371), .Z(n108) );
  IVP U309 ( .A(n1371), .Z(n109) );
  IVP U333 ( .A(n1371), .Z(n110) );
  IVP U335 ( .A(n1372), .Z(n111) );
  IVP U337 ( .A(n1372), .Z(n112) );
  IVP U339 ( .A(n1372), .Z(n113) );
  IVP U341 ( .A(n1372), .Z(n114) );
  IVP U343 ( .A(n1372), .Z(n115) );
  IVP U345 ( .A(n1373), .Z(n116) );
  IVP U347 ( .A(n1373), .Z(n117) );
  IVP U349 ( .A(n1373), .Z(n118) );
  IVP U351 ( .A(n1373), .Z(n119) );
  IVP U353 ( .A(n1373), .Z(n120) );
  IVP U355 ( .A(n1374), .Z(n121) );
  IVP U357 ( .A(n1374), .Z(n122) );
  IVP U359 ( .A(n1374), .Z(n123) );
  IVP U361 ( .A(n1374), .Z(n124) );
  IVP U363 ( .A(n1374), .Z(n125) );
  IVP U365 ( .A(n1375), .Z(n126) );
  IVP U367 ( .A(n1375), .Z(n127) );
  IVP U369 ( .A(n1375), .Z(n128) );
  IVP U371 ( .A(n1375), .Z(n129) );
  IVP U373 ( .A(n1375), .Z(n130) );
  IVP U375 ( .A(n1376), .Z(n131) );
  IVP U377 ( .A(n1376), .Z(n132) );
  IVP U379 ( .A(n1376), .Z(n133) );
  IVP U381 ( .A(n1376), .Z(n134) );
  IVP U383 ( .A(n1376), .Z(n135) );
  IVP U385 ( .A(n1377), .Z(n136) );
  IVP U387 ( .A(n1377), .Z(n137) );
  IVP U389 ( .A(n1377), .Z(n138) );
  IVP U391 ( .A(n1377), .Z(n139) );
  IVP U393 ( .A(n1377), .Z(n140) );
  IVP U395 ( .A(n1378), .Z(n141) );
  IVP U397 ( .A(n1378), .Z(n142) );
  IVP U399 ( .A(n1378), .Z(n143) );
  IVP U401 ( .A(n1378), .Z(n144) );
  IVP U403 ( .A(n1378), .Z(n145) );
  IVP U405 ( .A(n1379), .Z(n146) );
  IVP U407 ( .A(n1379), .Z(n147) );
  IVP U409 ( .A(n1379), .Z(n148) );
  IVP U411 ( .A(n1379), .Z(n149) );
  IVP U413 ( .A(n1379), .Z(n150) );
  IVP U415 ( .A(n1380), .Z(n151) );
  IVP U417 ( .A(n1380), .Z(n152) );
  IVP U419 ( .A(n1380), .Z(n153) );
  IVP U421 ( .A(n1380), .Z(n154) );
  IVP U423 ( .A(n1380), .Z(n155) );
  IVP U425 ( .A(n1381), .Z(n156) );
  IVP U427 ( .A(n1381), .Z(n157) );
  IVP U429 ( .A(n1381), .Z(n158) );
  IVP U431 ( .A(n1381), .Z(n159) );
  IVP U433 ( .A(n1381), .Z(n160) );
  IVP U435 ( .A(n1382), .Z(n161) );
  IVP U437 ( .A(n1382), .Z(n162) );
  IVP U439 ( .A(n1382), .Z(n163) );
  IVP U441 ( .A(n1382), .Z(n164) );
  IVP U443 ( .A(n1382), .Z(n165) );
  IVP U445 ( .A(n1383), .Z(n166) );
  IVP U447 ( .A(n1383), .Z(n167) );
  IVP U449 ( .A(n1383), .Z(n168) );
  IVP U451 ( .A(n1383), .Z(n169) );
  IVP U453 ( .A(n1383), .Z(n170) );
  IVP U455 ( .A(n1384), .Z(n171) );
  IVP U457 ( .A(n1384), .Z(n172) );
  IVP U459 ( .A(n1384), .Z(n173) );
  IVP U461 ( .A(n1384), .Z(n174) );
  IVP U463 ( .A(n1384), .Z(n175) );
  IVP U465 ( .A(n1385), .Z(n176) );
  IVP U467 ( .A(n1385), .Z(n177) );
  IVP U469 ( .A(n1385), .Z(n178) );
  IVP U471 ( .A(n1385), .Z(n179) );
  IVP U473 ( .A(n1385), .Z(n180) );
  IVP U475 ( .A(n1386), .Z(n181) );
  IVP U477 ( .A(n1386), .Z(n182) );
  IVP U479 ( .A(n1386), .Z(n183) );
  IVP U481 ( .A(n1386), .Z(n184) );
  IVP U483 ( .A(n1386), .Z(n185) );
  IVP U485 ( .A(n1387), .Z(n186) );
  IVP U487 ( .A(n1387), .Z(n187) );
  IVP U489 ( .A(n1387), .Z(n188) );
  IVP U491 ( .A(n1387), .Z(n189) );
  IVP U493 ( .A(n1387), .Z(n190) );
  IVP U495 ( .A(n1388), .Z(n191) );
  IVP U497 ( .A(n1388), .Z(n192) );
  IVP U499 ( .A(n1388), .Z(n193) );
  IVP U501 ( .A(n1388), .Z(n194) );
  IVP U503 ( .A(n1388), .Z(n195) );
  IVP U505 ( .A(n1389), .Z(n196) );
  IVP U507 ( .A(n1389), .Z(n197) );
  IVP U509 ( .A(n1389), .Z(n198) );
  IVP U511 ( .A(n1389), .Z(n199) );
  IVP U513 ( .A(n1389), .Z(n200) );
  IVP U515 ( .A(n1422), .Z(n201) );
  IVP U517 ( .A(n1422), .Z(n202) );
  IVP U519 ( .A(n1422), .Z(n203) );
  IVP U521 ( .A(n1422), .Z(n204) );
  IVP U523 ( .A(n1422), .Z(n205) );
  IVP U525 ( .A(n1423), .Z(n206) );
  IVP U527 ( .A(n1423), .Z(n207) );
  IVP U529 ( .A(n1423), .Z(n208) );
  IVP U531 ( .A(n1423), .Z(n209) );
  IVP U533 ( .A(n1423), .Z(n210) );
  IVP U535 ( .A(n1424), .Z(n211) );
  IVP U537 ( .A(n1424), .Z(n212) );
  IVP U539 ( .A(n1424), .Z(n213) );
  IVP U541 ( .A(n1424), .Z(n214) );
  IVP U543 ( .A(n1424), .Z(n215) );
  IVP U545 ( .A(n1425), .Z(n216) );
  IVP U547 ( .A(n1425), .Z(n217) );
  IVP U549 ( .A(n1425), .Z(n218) );
  IVP U551 ( .A(n1425), .Z(n219) );
  IVP U553 ( .A(n1425), .Z(n220) );
  IVP U555 ( .A(n1426), .Z(n221) );
  IVP U557 ( .A(n1426), .Z(n222) );
  IVP U559 ( .A(n1426), .Z(n223) );
  IVP U561 ( .A(n1426), .Z(n224) );
  IVP U563 ( .A(n1426), .Z(n225) );
  IVP U565 ( .A(n1427), .Z(n226) );
  IVP U567 ( .A(n1427), .Z(n227) );
  IVP U569 ( .A(n1427), .Z(n228) );
  IVP U571 ( .A(n1427), .Z(n229) );
  IVP U573 ( .A(n1427), .Z(n230) );
  IVP U575 ( .A(n1428), .Z(n231) );
  IVP U577 ( .A(n1428), .Z(n232) );
  IVP U579 ( .A(n1428), .Z(n233) );
  IVP U581 ( .A(n1428), .Z(n234) );
  IVP U583 ( .A(n1428), .Z(n235) );
  IVP U585 ( .A(n1429), .Z(n236) );
  IVP U587 ( .A(n1429), .Z(n237) );
  IVP U589 ( .A(n1429), .Z(n238) );
  IVP U591 ( .A(n1429), .Z(n239) );
  IVP U593 ( .A(n1429), .Z(n240) );
  IVP U595 ( .A(n1430), .Z(n241) );
  IVP U597 ( .A(n1430), .Z(n242) );
  IVP U599 ( .A(n1430), .Z(n243) );
  IVP U601 ( .A(n1430), .Z(n244) );
  IVP U603 ( .A(n1430), .Z(n245) );
  IVP U605 ( .A(n1431), .Z(n246) );
  IVP U607 ( .A(n1431), .Z(n247) );
  IVP U609 ( .A(n1431), .Z(n248) );
  IVP U611 ( .A(n1431), .Z(n249) );
  IVP U613 ( .A(n1431), .Z(n250) );
  IVP U615 ( .A(n1432), .Z(n251) );
  IVP U617 ( .A(n1432), .Z(n252) );
  IVP U619 ( .A(n1432), .Z(n253) );
  IVP U621 ( .A(n1432), .Z(n254) );
  IVP U623 ( .A(n1432), .Z(n255) );
  IVP U625 ( .A(n1433), .Z(n256) );
  IVP U627 ( .A(n1433), .Z(n257) );
  IVP U629 ( .A(n1433), .Z(n258) );
  IVP U631 ( .A(n1433), .Z(n259) );
  IVP U633 ( .A(n1433), .Z(n260) );
  IVP U635 ( .A(n1434), .Z(n261) );
  IVP U637 ( .A(n1434), .Z(n262) );
  IVP U639 ( .A(n1434), .Z(n263) );
  IVP U641 ( .A(n1434), .Z(n264) );
  IVP U643 ( .A(n1434), .Z(n265) );
  IVP U645 ( .A(n1435), .Z(n266) );
  IVP U647 ( .A(n1435), .Z(n267) );
  IVP U649 ( .A(n1435), .Z(n268) );
  IVP U651 ( .A(n1435), .Z(n269) );
  IVP U653 ( .A(n1435), .Z(n270) );
  IVP U655 ( .A(n1436), .Z(n271) );
  IVP U657 ( .A(n1436), .Z(n272) );
  IVP U659 ( .A(n1436), .Z(n273) );
  IVP U661 ( .A(n1436), .Z(n274) );
  IVP U663 ( .A(n1436), .Z(n275) );
  IVP U665 ( .A(n1437), .Z(n276) );
  IVP U667 ( .A(n1437), .Z(n277) );
  IVP U669 ( .A(n1437), .Z(n278) );
  IVP U671 ( .A(n1437), .Z(n279) );
  IVP U673 ( .A(n1437), .Z(n280) );
  IVP U675 ( .A(n1438), .Z(n281) );
  IVP U677 ( .A(n1438), .Z(n282) );
  IVP U679 ( .A(n1438), .Z(n283) );
  IVP U681 ( .A(n1438), .Z(n284) );
  IVP U683 ( .A(n1438), .Z(n285) );
  IVP U685 ( .A(n1439), .Z(n286) );
  IVP U687 ( .A(n1439), .Z(n287) );
  IVP U689 ( .A(n1439), .Z(n288) );
  IVP U691 ( .A(n1439), .Z(n289) );
  IVP U693 ( .A(n1439), .Z(n290) );
  IVP U695 ( .A(n1440), .Z(n291) );
  IVP U697 ( .A(n1440), .Z(n292) );
  IVP U699 ( .A(n1440), .Z(n293) );
  IVP U701 ( .A(n1440), .Z(n294) );
  IVP U703 ( .A(n1440), .Z(n295) );
  IVP U705 ( .A(n1441), .Z(n296) );
  IVP U707 ( .A(n1441), .Z(n297) );
  IVP U709 ( .A(n1441), .Z(n298) );
  IVP U711 ( .A(n1441), .Z(n299) );
  IVP U713 ( .A(n1441), .Z(n300) );
  IVP U715 ( .A(n1442), .Z(n301) );
  IVP U717 ( .A(n1442), .Z(n302) );
  IVP U719 ( .A(n1442), .Z(n303) );
  IVP U721 ( .A(n1442), .Z(n304) );
  IVP U723 ( .A(n1442), .Z(n305) );
  IVP U725 ( .A(n1443), .Z(n306) );
  IVP U727 ( .A(n1443), .Z(n307) );
  IVP U729 ( .A(n1443), .Z(n308) );
  IVP U731 ( .A(n1443), .Z(n309) );
  IVP U733 ( .A(n1443), .Z(n310) );
  IVP U735 ( .A(n1444), .Z(n311) );
  IVP U737 ( .A(n1444), .Z(n312) );
  IVP U739 ( .A(n1444), .Z(n313) );
  IVP U741 ( .A(n1444), .Z(n314) );
  IVP U743 ( .A(n1444), .Z(n315) );
  IVP U745 ( .A(n1445), .Z(n316) );
  IVP U747 ( .A(n1445), .Z(n317) );
  IVP U749 ( .A(n1445), .Z(n318) );
  IVP U751 ( .A(n1445), .Z(n319) );
  IVP U753 ( .A(n1445), .Z(n320) );
  IVP U755 ( .A(n1446), .Z(n321) );
  IVP U757 ( .A(n1446), .Z(n322) );
  IVP U759 ( .A(n1446), .Z(n323) );
  IVP U761 ( .A(n1446), .Z(n324) );
  IVP U763 ( .A(n1446), .Z(n325) );
  IVP U765 ( .A(n1447), .Z(n326) );
  IVP U767 ( .A(n1447), .Z(n327) );
  IVP U769 ( .A(n1447), .Z(n328) );
  IVP U771 ( .A(n1447), .Z(n329) );
  IVP U773 ( .A(n1447), .Z(n330) );
  IVP U775 ( .A(n1448), .Z(n331) );
  IVP U777 ( .A(n1448), .Z(n332) );
  IVP U779 ( .A(n1448), .Z(n333) );
  IVP U781 ( .A(n1448), .Z(n334) );
  IVP U783 ( .A(n1448), .Z(n335) );
  IVP U785 ( .A(n1449), .Z(n336) );
  IVP U787 ( .A(n1449), .Z(n337) );
  IVP U789 ( .A(n1449), .Z(n338) );
  IVP U791 ( .A(n1449), .Z(n339) );
  IVP U793 ( .A(n1449), .Z(n340) );
  IVP U795 ( .A(n1450), .Z(n341) );
  IVP U797 ( .A(n1450), .Z(n342) );
  IVP U799 ( .A(n1450), .Z(n343) );
  IVP U801 ( .A(n1450), .Z(n344) );
  IVP U803 ( .A(n1450), .Z(n345) );
  IVP U805 ( .A(n1451), .Z(n346) );
  IVP U807 ( .A(n1451), .Z(n347) );
  IVP U809 ( .A(n1451), .Z(n348) );
  IVP U811 ( .A(n1451), .Z(n349) );
  IVP U813 ( .A(n1451), .Z(n350) );
  IVP U815 ( .A(n1452), .Z(n351) );
  IVP U817 ( .A(n1452), .Z(n352) );
  IVP U819 ( .A(n1452), .Z(n353) );
  IVP U821 ( .A(n1452), .Z(n354) );
  IVP U823 ( .A(n1452), .Z(n355) );
  IVP U825 ( .A(n1453), .Z(n356) );
  IVP U827 ( .A(n1453), .Z(n357) );
  IVP U829 ( .A(n1453), .Z(n358) );
  IVP U831 ( .A(n1453), .Z(n359) );
  IVP U833 ( .A(n1453), .Z(n360) );
  IVP U835 ( .A(n199), .Z(n361) );
  IVP U837 ( .A(n196), .Z(n362) );
  IVP U839 ( .A(n197), .Z(n363) );
  IVP U841 ( .A(n198), .Z(n364) );
  IVP U843 ( .A(n1454), .Z(n365) );
  IVP U845 ( .A(n1454), .Z(n366) );
  IVP U847 ( .A(n1454), .Z(n367) );
  IVP U849 ( .A(n1454), .Z(n368) );
  IVP U851 ( .A(n1454), .Z(n369) );
  IVP U853 ( .A(n1455), .Z(n370) );
  IVP U855 ( .A(n1455), .Z(n371) );
  IVP U857 ( .A(n1455), .Z(n372) );
  IVP U859 ( .A(n1455), .Z(n373) );
  IVP U861 ( .A(n1455), .Z(n374) );
  IVP U863 ( .A(n1456), .Z(n375) );
  IVP U865 ( .A(n1456), .Z(n376) );
  IVP U867 ( .A(n1456), .Z(n377) );
  IVP U869 ( .A(n1456), .Z(n378) );
  IVP U871 ( .A(n1456), .Z(n379) );
  IVP U873 ( .A(n1457), .Z(n380) );
  IVP U875 ( .A(n1457), .Z(n381) );
  IVP U877 ( .A(n1457), .Z(n382) );
  IVP U879 ( .A(n1457), .Z(n383) );
  IVP U881 ( .A(n1457), .Z(n384) );
  IVP U883 ( .A(n1458), .Z(n385) );
  IVP U885 ( .A(n1458), .Z(n386) );
  IVP U887 ( .A(n1458), .Z(n387) );
  IVP U889 ( .A(n1458), .Z(n388) );
  IVP U891 ( .A(n1458), .Z(n389) );
  IVP U893 ( .A(n1459), .Z(n390) );
  IVP U895 ( .A(n1459), .Z(n391) );
  IVP U897 ( .A(n1459), .Z(n392) );
  IVP U899 ( .A(n1459), .Z(n393) );
  IVP U901 ( .A(n1459), .Z(n394) );
  IVP U903 ( .A(n1460), .Z(n395) );
  IVP U905 ( .A(n1460), .Z(n396) );
  IVP U907 ( .A(n1460), .Z(n397) );
  IVP U909 ( .A(n1460), .Z(n398) );
  IVP U911 ( .A(n1460), .Z(n399) );
  IVP U913 ( .A(n1461), .Z(n400) );
  IVP U915 ( .A(n1461), .Z(n401) );
  IVP U917 ( .A(n1461), .Z(n402) );
  IVP U919 ( .A(n1461), .Z(n403) );
  IVP U921 ( .A(n1461), .Z(n404) );
  IVP U923 ( .A(n1462), .Z(n405) );
  IVP U925 ( .A(n1462), .Z(n406) );
  IVP U927 ( .A(n1462), .Z(n407) );
  IVP U929 ( .A(n1462), .Z(n408) );
  IVP U931 ( .A(n1462), .Z(n409) );
  IVP U933 ( .A(n1463), .Z(n465) );
  IVP U935 ( .A(n1463), .Z(n466) );
  IVP U937 ( .A(n1463), .Z(n467) );
  IVP U939 ( .A(n1463), .Z(n468) );
  IVP U941 ( .A(n1463), .Z(n469) );
  IVP U943 ( .A(n1464), .Z(n470) );
  IVP U945 ( .A(n1464), .Z(n471) );
  IVP U947 ( .A(n1464), .Z(n472) );
  IVP U949 ( .A(n1464), .Z(n473) );
  IVP U951 ( .A(n1464), .Z(n474) );
  IVP U953 ( .A(n1465), .Z(n475) );
  IVP U955 ( .A(n1465), .Z(n476) );
  IVP U957 ( .A(n1465), .Z(n477) );
  IVP U959 ( .A(n1465), .Z(n478) );
  IVP U961 ( .A(n1465), .Z(n479) );
  IVP U963 ( .A(n1466), .Z(n480) );
  IVP U965 ( .A(n1466), .Z(n481) );
  IVP U967 ( .A(n1466), .Z(n482) );
  IVP U969 ( .A(n1466), .Z(n483) );
  IVP U971 ( .A(n1466), .Z(n484) );
  IVP U973 ( .A(n1467), .Z(n485) );
  IVP U975 ( .A(n1467), .Z(n486) );
  IVP U977 ( .A(n1467), .Z(n487) );
  IVP U979 ( .A(n1467), .Z(n488) );
  IVP U981 ( .A(n1467), .Z(n489) );
  IVP U983 ( .A(n1468), .Z(n490) );
  IVP U985 ( .A(n1468), .Z(n491) );
  IVP U987 ( .A(n1468), .Z(n492) );
  IVP U989 ( .A(n1468), .Z(n493) );
  IVP U991 ( .A(n1468), .Z(n494) );
  IVP U993 ( .A(n1469), .Z(n495) );
  IVP U995 ( .A(n1469), .Z(n496) );
  IVP U997 ( .A(n1469), .Z(n497) );
  IVP U999 ( .A(n1469), .Z(n498) );
  IVP U1001 ( .A(n1469), .Z(n499) );
  IVP U1003 ( .A(n1470), .Z(n500) );
  IVP U1005 ( .A(n1470), .Z(n501) );
  IVP U1007 ( .A(n1470), .Z(n502) );
  IVP U1009 ( .A(n1470), .Z(n503) );
  IVP U1011 ( .A(n1470), .Z(n504) );
  IVP U1013 ( .A(n1471), .Z(n505) );
  IVP U1015 ( .A(n1471), .Z(n506) );
  IVP U1017 ( .A(n1471), .Z(n507) );
  IVP U1019 ( .A(n1471), .Z(n508) );
  IVP U1021 ( .A(n1471), .Z(n509) );
  IVP U1023 ( .A(n1472), .Z(n565) );
  IVP U1025 ( .A(n1472), .Z(n566) );
  IVP U1027 ( .A(n1472), .Z(n567) );
  IVP U1029 ( .A(n1472), .Z(n568) );
  IVP U1031 ( .A(n1472), .Z(n569) );
  IVP U1033 ( .A(n1473), .Z(n570) );
  IVP U1035 ( .A(n1473), .Z(n571) );
  IVP U1037 ( .A(n1473), .Z(n572) );
  IVP U1039 ( .A(n1473), .Z(n573) );
  IVP U1041 ( .A(n1473), .Z(n574) );
  IVP U1043 ( .A(n1474), .Z(n575) );
  IVP U1045 ( .A(n1474), .Z(n576) );
  IVP U1047 ( .A(n1474), .Z(n577) );
  IVP U1049 ( .A(n1474), .Z(n578) );
  IVP U1051 ( .A(n1474), .Z(n579) );
  IVP U1053 ( .A(n1475), .Z(n580) );
  IVP U1055 ( .A(n1475), .Z(n581) );
  IVP U1057 ( .A(n1475), .Z(n582) );
  IVP U1059 ( .A(n1475), .Z(n583) );
  IVP U1061 ( .A(n1475), .Z(n584) );
  IVP U1063 ( .A(n1476), .Z(n585) );
  IVP U1065 ( .A(n1476), .Z(n586) );
  IVP U1067 ( .A(n1476), .Z(n587) );
  IVP U1069 ( .A(n1476), .Z(n588) );
  IVP U1071 ( .A(n1476), .Z(n589) );
  IVP U1073 ( .A(n1477), .Z(n590) );
  IVP U1075 ( .A(n1477), .Z(n591) );
  IVP U1077 ( .A(n1477), .Z(n592) );
  IVP U1079 ( .A(n1477), .Z(n593) );
  IVP U1081 ( .A(n1477), .Z(n594) );
  IVP U1083 ( .A(n1478), .Z(n595) );
  IVP U1085 ( .A(n1478), .Z(n596) );
  IVP U1087 ( .A(n1478), .Z(n597) );
  IVP U1089 ( .A(n1478), .Z(n598) );
  IVP U1091 ( .A(n1478), .Z(n599) );
  IVP U1093 ( .A(n1479), .Z(n600) );
  IVP U1095 ( .A(n1479), .Z(n601) );
  IVP U1097 ( .A(n1479), .Z(n602) );
  IVP U1099 ( .A(n1479), .Z(n603) );
  IVP U1101 ( .A(n1479), .Z(n604) );
  IVP U1103 ( .A(n1480), .Z(n605) );
  IVP U1105 ( .A(n1480), .Z(n606) );
  IVP U1107 ( .A(n1480), .Z(n607) );
  IVP U1109 ( .A(n1480), .Z(n608) );
  IVP U1111 ( .A(n1480), .Z(n609) );
  IVP U1113 ( .A(n1481), .Z(n632) );
  IVP U1115 ( .A(n1481), .Z(n633) );
  IVP U1117 ( .A(n1481), .Z(n634) );
  IVP U1119 ( .A(n1481), .Z(n635) );
  IVP U1121 ( .A(n1481), .Z(n636) );
  IVP U1123 ( .A(n1482), .Z(n637) );
  IVP U1125 ( .A(n1482), .Z(n638) );
  IVP U1127 ( .A(n1482), .Z(n639) );
  IVP U1129 ( .A(n1482), .Z(n640) );
  IVP U1131 ( .A(n1482), .Z(n641) );
  IVP U1133 ( .A(n1483), .Z(n642) );
  IVP U1135 ( .A(n1483), .Z(n643) );
  IVP U1137 ( .A(n1483), .Z(n644) );
  IVP U1139 ( .A(n1483), .Z(n645) );
  IVP U1141 ( .A(n1483), .Z(n646) );
  IVP U1143 ( .A(n1484), .Z(n647) );
  IVP U1145 ( .A(n1484), .Z(n648) );
  IVP U1147 ( .A(n1484), .Z(n649) );
  IVP U1149 ( .A(n1484), .Z(n650) );
  IVP U1151 ( .A(n1484), .Z(n651) );
  IVP U1153 ( .A(n1485), .Z(n652) );
  IVP U1155 ( .A(n1485), .Z(n653) );
  IVP U1157 ( .A(n1485), .Z(n654) );
  IVP U1159 ( .A(n1485), .Z(n655) );
  IVP U1161 ( .A(n1485), .Z(n656) );
  IVP U1163 ( .A(n1518), .Z(n657) );
  IVP U1165 ( .A(n1518), .Z(n658) );
  IVP U1167 ( .A(n1518), .Z(n659) );
  IVP U1169 ( .A(n1518), .Z(n660) );
  IVP U1171 ( .A(n1518), .Z(n661) );
  IVP U1173 ( .A(n1518), .Z(n662) );
  IVP U1175 ( .A(n1518), .Z(n663) );
  IVP U1177 ( .A(b[1]), .Z(n664) );
  IVP U1179 ( .A(b[1]), .Z(n665) );
  IVP U1181 ( .A(b[1]), .Z(n666) );
  IVP U1183 ( .A(b[2]), .Z(n667) );
  IVP U1185 ( .A(b[2]), .Z(n668) );
  IVP U1187 ( .A(b[2]), .Z(n669) );
  IVP U1189 ( .A(b[3]), .Z(n670) );
  IVP U1191 ( .A(b[3]), .Z(n671) );
  IVP U1193 ( .A(b[3]), .Z(n672) );
  IVP U1195 ( .A(b[4]), .Z(n673) );
  IVP U1197 ( .A(b[4]), .Z(n674) );
  IVP U1199 ( .A(b[4]), .Z(n675) );
  IVP U1201 ( .A(b[5]), .Z(n676) );
  IVP U1203 ( .A(b[5]), .Z(n677) );
  IVP U1205 ( .A(b[5]), .Z(n678) );
  IVP U1207 ( .A(b[6]), .Z(n679) );
  IVP U1209 ( .A(b[6]), .Z(n680) );
  IVP U1211 ( .A(b[6]), .Z(n681) );
  IVP U1213 ( .A(b[7]), .Z(n682) );
  IVP U1215 ( .A(b[7]), .Z(n683) );
  IVP U1217 ( .A(b[7]), .Z(n684) );
  IVP U1219 ( .A(b[8]), .Z(n685) );
  IVP U1221 ( .A(b[8]), .Z(n686) );
  IVP U1223 ( .A(b[8]), .Z(n687) );
  IVP U1225 ( .A(b[9]), .Z(n688) );
  IVP U1227 ( .A(b[9]), .Z(n689) );
  IVP U1229 ( .A(b[9]), .Z(n690) );
  IVP U1231 ( .A(b[10]), .Z(n691) );
  IVP U1233 ( .A(b[10]), .Z(n692) );
  IVP U1235 ( .A(b[10]), .Z(n693) );
  IVP U1237 ( .A(b[11]), .Z(n694) );
  IVP U1239 ( .A(b[11]), .Z(n695) );
  IVP U1241 ( .A(b[11]), .Z(n696) );
  IVP U1243 ( .A(b[12]), .Z(n697) );
  IVP U1245 ( .A(b[12]), .Z(n698) );
  IVP U1247 ( .A(b[12]), .Z(n699) );
  IVP U1249 ( .A(b[13]), .Z(n700) );
  IVP U1251 ( .A(b[13]), .Z(n701) );
  IVP U1253 ( .A(b[13]), .Z(n702) );
  IVP U1255 ( .A(b[14]), .Z(n703) );
  IVP U1257 ( .A(b[14]), .Z(n704) );
  IVP U1259 ( .A(b[14]), .Z(n705) );
  IVP U1261 ( .A(b[15]), .Z(n706) );
  IVP U1263 ( .A(b[15]), .Z(n707) );
  IVP U1265 ( .A(b[15]), .Z(n708) );
  IVP U1267 ( .A(b[16]), .Z(n709) );
  IVP U1269 ( .A(b[16]), .Z(n732) );
  IVP U1271 ( .A(b[16]), .Z(n733) );
  IVP U1273 ( .A(b[17]), .Z(n734) );
  IVP U1275 ( .A(b[17]), .Z(n735) );
  IVP U1277 ( .A(b[17]), .Z(n736) );
  IVP U1279 ( .A(b[18]), .Z(n737) );
  IVP U1281 ( .A(b[18]), .Z(n738) );
  IVP U1283 ( .A(b[18]), .Z(n739) );
  IVP U1285 ( .A(b[19]), .Z(n740) );
  IVP U1287 ( .A(b[19]), .Z(n741) );
  IVP U1289 ( .A(b[19]), .Z(n742) );
  IVP U1291 ( .A(b[20]), .Z(n743) );
  IVP U1293 ( .A(b[20]), .Z(n744) );
  IVP U1295 ( .A(b[20]), .Z(n745) );
  IVP U1297 ( .A(b[21]), .Z(n746) );
  IVP U1299 ( .A(b[21]), .Z(n747) );
  IVP U1301 ( .A(b[21]), .Z(n748) );
  IVP U1303 ( .A(b[22]), .Z(n749) );
  IVP U1305 ( .A(b[22]), .Z(n750) );
  IVP U1307 ( .A(b[22]), .Z(n751) );
  IVP U1309 ( .A(b[23]), .Z(n752) );
  IVP U1311 ( .A(b[23]), .Z(n753) );
  IVP U1313 ( .A(b[23]), .Z(n754) );
  IVP U1315 ( .A(b[24]), .Z(n755) );
  IVP U1317 ( .A(b[24]), .Z(n756) );
  IVP U1319 ( .A(b[24]), .Z(n757) );
  IVP U1321 ( .A(b[25]), .Z(n758) );
  IVP U1323 ( .A(b[25]), .Z(n759) );
  IVP U1325 ( .A(b[25]), .Z(n760) );
  IVP U1327 ( .A(b[26]), .Z(n761) );
  IVP U1329 ( .A(b[26]), .Z(n762) );
  IVP U1331 ( .A(b[26]), .Z(n763) );
  IVP U1333 ( .A(b[27]), .Z(n764) );
  IVP U1335 ( .A(b[27]), .Z(n765) );
  IVP U1337 ( .A(b[27]), .Z(n766) );
  IVP U1339 ( .A(b[28]), .Z(n767) );
  IVP U1341 ( .A(b[28]), .Z(n768) );
  IVP U1343 ( .A(b[28]), .Z(n769) );
  IVP U1345 ( .A(b[29]), .Z(n770) );
  IVP U1347 ( .A(b[29]), .Z(n771) );
  IVP U1349 ( .A(b[29]), .Z(n772) );
  IVP U1351 ( .A(b[30]), .Z(n773) );
  IVP U1353 ( .A(b[30]), .Z(n774) );
  IVP U1355 ( .A(b[30]), .Z(n775) );
  IVP U1357 ( .A(b[31]), .Z(n776) );
  IVP U1359 ( .A(b[31]), .Z(n777) );
  IVP U1361 ( .A(b[31]), .Z(n778) );
  IVP U1363 ( .A(b[32]), .Z(n779) );
  IVP U1365 ( .A(b[32]), .Z(n780) );
  IVP U1367 ( .A(b[32]), .Z(n781) );
  IVP U1369 ( .A(b[33]), .Z(n782) );
  IVP U1371 ( .A(b[33]), .Z(n783) );
  IVP U1373 ( .A(b[33]), .Z(n784) );
  IVP U1375 ( .A(b[34]), .Z(n785) );
  IVP U1377 ( .A(b[34]), .Z(n786) );
  IVP U1379 ( .A(b[34]), .Z(n787) );
  IVP U1381 ( .A(b[35]), .Z(n788) );
  IVP U1383 ( .A(b[35]), .Z(n789) );
  IVP U1385 ( .A(b[35]), .Z(n790) );
  IVP U1387 ( .A(b[36]), .Z(n791) );
  IVP U1389 ( .A(b[36]), .Z(n792) );
  IVP U1391 ( .A(b[36]), .Z(n793) );
  IVP U1393 ( .A(b[37]), .Z(n794) );
  IVP U1395 ( .A(b[37]), .Z(n795) );
  IVP U1397 ( .A(b[37]), .Z(n796) );
  IVP U1399 ( .A(b[38]), .Z(n797) );
  IVP U1401 ( .A(b[38]), .Z(n798) );
  IVP U1403 ( .A(b[38]), .Z(n799) );
  IVP U1405 ( .A(b[39]), .Z(n800) );
  IVP U1407 ( .A(b[39]), .Z(n801) );
  IVP U1409 ( .A(b[39]), .Z(n802) );
  IVP U1411 ( .A(b[40]), .Z(n803) );
  IVP U1413 ( .A(b[40]), .Z(n804) );
  IVP U1415 ( .A(b[40]), .Z(n805) );
  IVP U1417 ( .A(b[41]), .Z(n806) );
  IVP U1419 ( .A(b[41]), .Z(n807) );
  IVP U1421 ( .A(b[41]), .Z(n808) );
  IVP U1423 ( .A(b[42]), .Z(n809) );
  IVP U1425 ( .A(b[42]), .Z(n810) );
  IVP U1427 ( .A(b[42]), .Z(n811) );
  IVP U1429 ( .A(b[43]), .Z(n812) );
  IVP U1431 ( .A(b[43]), .Z(n813) );
  IVP U1433 ( .A(b[43]), .Z(n814) );
  IVP U1435 ( .A(b[44]), .Z(n815) );
  IVP U1437 ( .A(b[44]), .Z(n816) );
  IVP U1439 ( .A(b[44]), .Z(n817) );
  IVP U1441 ( .A(b[45]), .Z(n818) );
  IVP U1443 ( .A(b[45]), .Z(n819) );
  IVP U1445 ( .A(b[45]), .Z(n820) );
  IVP U1447 ( .A(b[46]), .Z(n821) );
  IVP U1449 ( .A(b[46]), .Z(n822) );
  IVP U1451 ( .A(b[46]), .Z(n823) );
  IVP U1453 ( .A(b[47]), .Z(n824) );
  IVP U1455 ( .A(b[47]), .Z(n825) );
  IVP U1457 ( .A(b[47]), .Z(n826) );
  IVP U1459 ( .A(b[48]), .Z(n827) );
  IVP U1461 ( .A(b[48]), .Z(n828) );
  IVP U1463 ( .A(b[48]), .Z(n829) );
  IVP U1465 ( .A(b[49]), .Z(n830) );
  IVP U1467 ( .A(b[49]), .Z(n831) );
  IVP U1469 ( .A(b[49]), .Z(n832) );
  IVP U1471 ( .A(b[50]), .Z(n833) );
  IVP U1473 ( .A(b[50]), .Z(n834) );
  IVP U1475 ( .A(b[50]), .Z(n835) );
  IVP U1477 ( .A(b[51]), .Z(n836) );
  IVP U1479 ( .A(b[51]), .Z(n837) );
  IVP U1481 ( .A(b[51]), .Z(n838) );
  IVP U1483 ( .A(b[52]), .Z(n839) );
  IVP U1485 ( .A(b[52]), .Z(n840) );
  IVP U1487 ( .A(b[52]), .Z(n841) );
  IVP U1489 ( .A(b[53]), .Z(n842) );
  IVP U1491 ( .A(b[53]), .Z(n843) );
  IVP U1493 ( .A(b[53]), .Z(n844) );
  IVP U1495 ( .A(b[54]), .Z(n845) );
  IVP U1497 ( .A(b[54]), .Z(n846) );
  IVP U1499 ( .A(b[54]), .Z(n847) );
  IVP U1501 ( .A(b[55]), .Z(n848) );
  IVP U1503 ( .A(b[55]), .Z(n849) );
  IVP U1505 ( .A(b[55]), .Z(n850) );
  IVP U1507 ( .A(b[56]), .Z(n851) );
  IVP U1509 ( .A(b[56]), .Z(n852) );
  IVP U1511 ( .A(b[56]), .Z(n853) );
  IVP U1513 ( .A(b[57]), .Z(n854) );
  IVP U1515 ( .A(b[57]), .Z(n855) );
  IVP U1517 ( .A(b[57]), .Z(n856) );
  IVP U1519 ( .A(b[58]), .Z(n857) );
  IVP U1521 ( .A(b[58]), .Z(n858) );
  IVP U1523 ( .A(b[58]), .Z(n859) );
  IVP U1525 ( .A(b[59]), .Z(n860) );
  IVP U1527 ( .A(b[59]), .Z(n861) );
  IVP U1529 ( .A(b[59]), .Z(n862) );
  IVP U1531 ( .A(b[60]), .Z(n863) );
  IVP U1533 ( .A(b[60]), .Z(n864) );
  IVP U1535 ( .A(b[60]), .Z(n865) );
  IVP U1537 ( .A(b[61]), .Z(n866) );
  IVP U1539 ( .A(b[61]), .Z(n867) );
  IVP U1541 ( .A(b[61]), .Z(n868) );
  IVP U1543 ( .A(b[62]), .Z(n869) );
  IVP U1545 ( .A(b[62]), .Z(n870) );
  IVP U1547 ( .A(b[62]), .Z(n871) );
  IVP U1549 ( .A(b[63]), .Z(n872) );
  IVP U1551 ( .A(b[63]), .Z(n873) );
  IVP U1553 ( .A(b[63]), .Z(n874) );
  IVP U1555 ( .A(b[0]), .Z(n1069) );
  IVP U1557 ( .A(n1357), .Z(n1070) );
  IVP U1559 ( .A(n1324), .Z(n1071) );
  IVP U1561 ( .A(a[63]), .Z(n1072) );
  IVP U1563 ( .A(n1356), .Z(n1073) );
  IVP U1565 ( .A(n1323), .Z(n1074) );
  IVP U1567 ( .A(a[61]), .Z(n1075) );
  IVP U1569 ( .A(n1355), .Z(n1076) );
  IVP U1571 ( .A(n1322), .Z(n1077) );
  IVP U1573 ( .A(a[59]), .Z(n1078) );
  IVP U1575 ( .A(n1354), .Z(n1079) );
  IVP U1577 ( .A(n1321), .Z(n1080) );
  IVP U1579 ( .A(a[57]), .Z(n1081) );
  IVP U1581 ( .A(n1353), .Z(n1082) );
  IVP U1583 ( .A(n1320), .Z(n1083) );
  IVP U1585 ( .A(a[55]), .Z(n1084) );
  IVP U1587 ( .A(n1352), .Z(n1085) );
  IVP U1589 ( .A(n1319), .Z(n1086) );
  IVP U1591 ( .A(a[53]), .Z(n1087) );
  IVP U1593 ( .A(n1351), .Z(n1088) );
  IVP U1595 ( .A(n1318), .Z(n1089) );
  IVP U1597 ( .A(a[51]), .Z(n1090) );
  IVP U1599 ( .A(n1350), .Z(n1091) );
  IVP U1601 ( .A(n1317), .Z(n1092) );
  IVP U1603 ( .A(a[49]), .Z(n1093) );
  IVP U1605 ( .A(n1349), .Z(n1094) );
  IVP U1607 ( .A(n1316), .Z(n1095) );
  IVP U1609 ( .A(a[47]), .Z(n1096) );
  IVP U1611 ( .A(n1348), .Z(n1097) );
  IVP U1613 ( .A(n1315), .Z(n1098) );
  IVP U1615 ( .A(a[45]), .Z(n1099) );
  IVP U1617 ( .A(n1347), .Z(n1100) );
  IVP U1619 ( .A(n1314), .Z(n1101) );
  IVP U1621 ( .A(a[43]), .Z(n1102) );
  IVP U1623 ( .A(n1346), .Z(n1103) );
  IVP U1625 ( .A(n1313), .Z(n1104) );
  IVP U1627 ( .A(a[41]), .Z(n1105) );
  IVP U1629 ( .A(n1345), .Z(n1106) );
  IVP U1631 ( .A(n1312), .Z(n1107) );
  IVP U1633 ( .A(a[39]), .Z(n1108) );
  IVP U1635 ( .A(n1344), .Z(n1109) );
  IVP U1637 ( .A(n1311), .Z(n1110) );
  IVP U1639 ( .A(a[37]), .Z(n1111) );
  IVP U1641 ( .A(n1343), .Z(n1112) );
  IVP U1643 ( .A(n1310), .Z(n1113) );
  IVP U1645 ( .A(a[35]), .Z(n1114) );
  IVP U1647 ( .A(n1342), .Z(n1115) );
  IVP U1649 ( .A(n1309), .Z(n1116) );
  IVP U1651 ( .A(a[33]), .Z(n1117) );
  IVP U1653 ( .A(n1341), .Z(n1118) );
  IVP U1655 ( .A(n1308), .Z(n1119) );
  IVP U1657 ( .A(a[31]), .Z(n1120) );
  IVP U1659 ( .A(n1340), .Z(n1121) );
  IVP U1661 ( .A(n1307), .Z(n1122) );
  IVP U1663 ( .A(a[29]), .Z(n1123) );
  IVP U1665 ( .A(n1339), .Z(n1124) );
  IVP U1667 ( .A(n1306), .Z(n1125) );
  IVP U1669 ( .A(a[27]), .Z(n1126) );
  IVP U1671 ( .A(n1338), .Z(n1127) );
  IVP U1673 ( .A(n1305), .Z(n1128) );
  IVP U1675 ( .A(a[25]), .Z(n1129) );
  IVP U1677 ( .A(n1337), .Z(n1130) );
  IVP U1679 ( .A(n1304), .Z(n1131) );
  IVP U1681 ( .A(a[23]), .Z(n1132) );
  IVP U1683 ( .A(n1336), .Z(n1133) );
  IVP U1685 ( .A(n1303), .Z(n1134) );
  IVP U1687 ( .A(a[21]), .Z(n1135) );
  IVP U1689 ( .A(n1335), .Z(n1136) );
  IVP U1691 ( .A(n1302), .Z(n1137) );
  IVP U1693 ( .A(a[19]), .Z(n1138) );
  IVP U1695 ( .A(n1334), .Z(n1139) );
  IVP U1697 ( .A(n1301), .Z(n1140) );
  IVP U1699 ( .A(a[17]), .Z(n1141) );
  IVP U1701 ( .A(n1333), .Z(n1142) );
  IVP U1703 ( .A(n1300), .Z(n1143) );
  IVP U1705 ( .A(a[15]), .Z(n1144) );
  IVP U1707 ( .A(n1332), .Z(n1145) );
  IVP U1709 ( .A(n1299), .Z(n1146) );
  IVP U1711 ( .A(a[13]), .Z(n1147) );
  IVP U1713 ( .A(n1331), .Z(n1148) );
  IVP U1715 ( .A(n1298), .Z(n1149) );
  IVP U1717 ( .A(a[11]), .Z(n1150) );
  IVP U1719 ( .A(n1330), .Z(n1151) );
  IVP U1721 ( .A(n1297), .Z(n1152) );
  IVP U1723 ( .A(a[9]), .Z(n1153) );
  IVP U1725 ( .A(n1329), .Z(n1154) );
  IVP U1727 ( .A(n1296), .Z(n1155) );
  IVP U1729 ( .A(a[7]), .Z(n1156) );
  IVP U1731 ( .A(n1328), .Z(n1157) );
  IVP U1733 ( .A(n1295), .Z(n1158) );
  IVP U1735 ( .A(a[5]), .Z(n1159) );
  IVP U1737 ( .A(n1327), .Z(n1160) );
  IVP U1739 ( .A(n1294), .Z(n1161) );
  IVP U1741 ( .A(a[3]), .Z(n1162) );
  IVP U1743 ( .A(n1326), .Z(n1163) );
  IVP U1745 ( .A(n1293), .Z(n1164) );
  IVP U1747 ( .A(a[1]), .Z(n1165) );
  IVP U1749 ( .A(a[0]), .Z(n1293) );
  EO U1750 ( .A(a[0]), .B(a[1]), .Z(n1486) );
  ND2 U1751 ( .A(n1486), .B(n1293), .Z(n1326) );
  EN U1752 ( .A(a[2]), .B(a[1]), .Z(n1294) );
  EO U1753 ( .A(a[2]), .B(a[3]), .Z(n1487) );
  ND2 U1754 ( .A(n1294), .B(n1487), .Z(n1327) );
  EN U1755 ( .A(a[4]), .B(a[3]), .Z(n1295) );
  EO U1756 ( .A(a[4]), .B(a[5]), .Z(n1488) );
  ND2 U1757 ( .A(n1295), .B(n1488), .Z(n1328) );
  EN U1758 ( .A(a[6]), .B(a[5]), .Z(n1296) );
  EO U1759 ( .A(a[6]), .B(a[7]), .Z(n1489) );
  ND2 U1760 ( .A(n1296), .B(n1489), .Z(n1329) );
  EN U1761 ( .A(a[8]), .B(a[7]), .Z(n1297) );
  EO U1762 ( .A(a[8]), .B(a[9]), .Z(n1490) );
  ND2 U1763 ( .A(n1297), .B(n1490), .Z(n1330) );
  EN U1764 ( .A(a[10]), .B(a[9]), .Z(n1298) );
  EO U1765 ( .A(a[10]), .B(a[11]), .Z(n1491) );
  ND2 U1766 ( .A(n1298), .B(n1491), .Z(n1331) );
  EN U1767 ( .A(a[12]), .B(a[11]), .Z(n1299) );
  EO U1768 ( .A(a[12]), .B(a[13]), .Z(n1492) );
  ND2 U1769 ( .A(n1299), .B(n1492), .Z(n1332) );
  EN U1770 ( .A(a[14]), .B(a[13]), .Z(n1300) );
  EO U1771 ( .A(a[14]), .B(a[15]), .Z(n1493) );
  ND2 U1772 ( .A(n1300), .B(n1493), .Z(n1333) );
  EN U1773 ( .A(a[16]), .B(a[15]), .Z(n1301) );
  EO U1774 ( .A(a[16]), .B(a[17]), .Z(n1494) );
  ND2 U1775 ( .A(n1301), .B(n1494), .Z(n1334) );
  EN U1776 ( .A(a[18]), .B(a[17]), .Z(n1302) );
  EO U1777 ( .A(a[18]), .B(a[19]), .Z(n1495) );
  ND2 U1778 ( .A(n1302), .B(n1495), .Z(n1335) );
  EN U1779 ( .A(a[20]), .B(a[19]), .Z(n1303) );
  EO U1780 ( .A(a[20]), .B(a[21]), .Z(n1496) );
  ND2 U1781 ( .A(n1303), .B(n1496), .Z(n1336) );
  EN U1782 ( .A(a[22]), .B(a[21]), .Z(n1304) );
  EO U1783 ( .A(a[22]), .B(a[23]), .Z(n1497) );
  ND2 U1784 ( .A(n1304), .B(n1497), .Z(n1337) );
  EN U1785 ( .A(a[24]), .B(a[23]), .Z(n1305) );
  EO U1786 ( .A(a[24]), .B(a[25]), .Z(n1498) );
  ND2 U1787 ( .A(n1305), .B(n1498), .Z(n1338) );
  EN U1788 ( .A(a[26]), .B(a[25]), .Z(n1306) );
  EO U1789 ( .A(a[26]), .B(a[27]), .Z(n1499) );
  ND2 U1790 ( .A(n1306), .B(n1499), .Z(n1339) );
  EN U1791 ( .A(a[28]), .B(a[27]), .Z(n1307) );
  EO U1792 ( .A(a[28]), .B(a[29]), .Z(n1500) );
  ND2 U1793 ( .A(n1307), .B(n1500), .Z(n1340) );
  EN U1794 ( .A(a[30]), .B(a[29]), .Z(n1308) );
  EO U1795 ( .A(a[30]), .B(a[31]), .Z(n1501) );
  ND2 U1796 ( .A(n1308), .B(n1501), .Z(n1341) );
  EN U1797 ( .A(a[32]), .B(a[31]), .Z(n1309) );
  EO U1798 ( .A(a[32]), .B(a[33]), .Z(n1502) );
  ND2 U1799 ( .A(n1309), .B(n1502), .Z(n1342) );
  EN U1800 ( .A(a[34]), .B(a[33]), .Z(n1310) );
  EO U1801 ( .A(a[34]), .B(a[35]), .Z(n1503) );
  ND2 U1802 ( .A(n1310), .B(n1503), .Z(n1343) );
  EN U1803 ( .A(a[36]), .B(a[35]), .Z(n1311) );
  EO U1804 ( .A(a[36]), .B(a[37]), .Z(n1504) );
  ND2 U1805 ( .A(n1311), .B(n1504), .Z(n1344) );
  EN U1806 ( .A(a[38]), .B(a[37]), .Z(n1312) );
  EO U1807 ( .A(a[38]), .B(a[39]), .Z(n1505) );
  ND2 U1808 ( .A(n1312), .B(n1505), .Z(n1345) );
  EN U1809 ( .A(a[40]), .B(a[39]), .Z(n1313) );
  EO U1810 ( .A(a[40]), .B(a[41]), .Z(n1506) );
  ND2 U1811 ( .A(n1313), .B(n1506), .Z(n1346) );
  EN U1812 ( .A(a[42]), .B(a[41]), .Z(n1314) );
  EO U1813 ( .A(a[42]), .B(a[43]), .Z(n1507) );
  ND2 U1814 ( .A(n1314), .B(n1507), .Z(n1347) );
  EN U1815 ( .A(a[44]), .B(a[43]), .Z(n1315) );
  EO U1816 ( .A(a[44]), .B(a[45]), .Z(n1508) );
  ND2 U1817 ( .A(n1315), .B(n1508), .Z(n1348) );
  EN U1818 ( .A(a[46]), .B(a[45]), .Z(n1316) );
  EO U1819 ( .A(a[46]), .B(a[47]), .Z(n1509) );
  ND2 U1820 ( .A(n1316), .B(n1509), .Z(n1349) );
  EN U1821 ( .A(a[48]), .B(a[47]), .Z(n1317) );
  EO U1822 ( .A(a[48]), .B(a[49]), .Z(n1510) );
  ND2 U1823 ( .A(n1317), .B(n1510), .Z(n1350) );
  EN U1824 ( .A(a[50]), .B(a[49]), .Z(n1318) );
  EO U1825 ( .A(a[50]), .B(a[51]), .Z(n1511) );
  ND2 U1826 ( .A(n1318), .B(n1511), .Z(n1351) );
  EN U1827 ( .A(a[52]), .B(a[51]), .Z(n1319) );
  EO U1828 ( .A(a[52]), .B(a[53]), .Z(n1512) );
  ND2 U1829 ( .A(n1319), .B(n1512), .Z(n1352) );
  EN U1830 ( .A(a[54]), .B(a[53]), .Z(n1320) );
  EO U1831 ( .A(a[54]), .B(a[55]), .Z(n1513) );
  ND2 U1832 ( .A(n1320), .B(n1513), .Z(n1353) );
  EN U1833 ( .A(a[56]), .B(a[55]), .Z(n1321) );
  EO U1834 ( .A(a[56]), .B(a[57]), .Z(n1514) );
  ND2 U1835 ( .A(n1321), .B(n1514), .Z(n1354) );
  EN U1836 ( .A(a[58]), .B(a[57]), .Z(n1322) );
  EO U1837 ( .A(a[58]), .B(a[59]), .Z(n1515) );
  ND2 U1838 ( .A(n1322), .B(n1515), .Z(n1355) );
  EN U1839 ( .A(a[60]), .B(a[59]), .Z(n1323) );
  EO U1840 ( .A(a[60]), .B(a[61]), .Z(n1516) );
  ND2 U1841 ( .A(n1323), .B(n1516), .Z(n1356) );
  EN U1842 ( .A(a[62]), .B(a[61]), .Z(n1324) );
  EO U1843 ( .A(a[62]), .B(a[63]), .Z(n1517) );
  ND2 U1844 ( .A(n1324), .B(n1517), .Z(n1357) );
  IVP U1846 ( .A(n10737), .Z(n1390) );
  IVP U1847 ( .A(n10732), .Z(n1391) );
  IVP U1848 ( .A(n10727), .Z(n1392) );
  IVP U1849 ( .A(n10722), .Z(n1393) );
  IVP U1850 ( .A(n10717), .Z(n1394) );
  IVP U1851 ( .A(n10712), .Z(n1395) );
  IVP U1852 ( .A(n10707), .Z(n1396) );
  IVP U1853 ( .A(n10702), .Z(n1397) );
  IVP U1854 ( .A(n10697), .Z(n1398) );
  IVP U1855 ( .A(n10692), .Z(n1399) );
  IVP U1856 ( .A(n10687), .Z(n1400) );
  IVP U1857 ( .A(n10682), .Z(n1401) );
  IVP U1858 ( .A(n10677), .Z(n1402) );
  IVP U1859 ( .A(n10672), .Z(n1403) );
  IVP U1860 ( .A(n10667), .Z(n1404) );
  IVP U1861 ( .A(n10662), .Z(n1405) );
  IVP U1862 ( .A(n10657), .Z(n1406) );
  IVP U1863 ( .A(n10652), .Z(n1407) );
  IVP U1864 ( .A(n10647), .Z(n1408) );
  IVP U1865 ( .A(n10642), .Z(n1409) );
  IVP U1866 ( .A(n10637), .Z(n1410) );
  IVP U1867 ( .A(n10632), .Z(n1411) );
  IVP U1868 ( .A(n10627), .Z(n1412) );
  IVP U1869 ( .A(n10622), .Z(n1413) );
  IVP U1870 ( .A(n10617), .Z(n1414) );
  IVP U1871 ( .A(n10612), .Z(n1415) );
  IVP U1872 ( .A(n10607), .Z(n1416) );
  IVP U1873 ( .A(n10602), .Z(n1417) );
  IVP U1874 ( .A(n10597), .Z(n1418) );
  IVP U1875 ( .A(n10592), .Z(n1419) );
  IVP U1876 ( .A(n10587), .Z(n1420) );
  IVP U1877 ( .A(n10582), .Z(n1421) );
  EN U1878 ( .A(n10253), .B(n10737), .Z(n1520) );
  EN U1879 ( .A(n10246), .B(n10737), .Z(n1521) );
  EN U1880 ( .A(n10243), .B(n10737), .Z(n1522) );
  EN U1881 ( .A(n10240), .B(n10737), .Z(n1523) );
  EN U1882 ( .A(n10237), .B(n10737), .Z(n1524) );
  EN U1883 ( .A(n10234), .B(n10737), .Z(n1525) );
  EN U1884 ( .A(n10231), .B(n10737), .Z(n1526) );
  EN U1885 ( .A(n10228), .B(n10737), .Z(n1527) );
  EN U1886 ( .A(n10225), .B(n10737), .Z(n1528) );
  EN U1887 ( .A(n10222), .B(n10736), .Z(n1529) );
  EN U1888 ( .A(n10219), .B(n10736), .Z(n1530) );
  EN U1889 ( .A(n10216), .B(n10736), .Z(n1531) );
  EN U1890 ( .A(n10213), .B(n10736), .Z(n1532) );
  EN U1891 ( .A(n10210), .B(n10736), .Z(n1533) );
  EN U1892 ( .A(n10207), .B(n10736), .Z(n1534) );
  EN U1893 ( .A(n10204), .B(n10736), .Z(n1535) );
  EN U1894 ( .A(n10201), .B(n10736), .Z(n1536) );
  EN U1895 ( .A(n10198), .B(n10736), .Z(n1537) );
  EN U1896 ( .A(n10195), .B(n10736), .Z(n1538) );
  EN U1897 ( .A(n10192), .B(n10736), .Z(n1539) );
  EN U1898 ( .A(n10189), .B(n10736), .Z(n1540) );
  EN U1899 ( .A(n10186), .B(n10736), .Z(n1541) );
  EN U1900 ( .A(n10183), .B(n10736), .Z(n1542) );
  EN U1901 ( .A(n10180), .B(n10735), .Z(n1543) );
  EN U1902 ( .A(n10177), .B(n10735), .Z(n1544) );
  EN U1903 ( .A(n10174), .B(n10735), .Z(n1545) );
  EN U1904 ( .A(n10171), .B(n10735), .Z(n1546) );
  EN U1905 ( .A(n10168), .B(n10735), .Z(n1547) );
  EN U1906 ( .A(n10165), .B(n10735), .Z(n1548) );
  EN U1907 ( .A(n10162), .B(n10735), .Z(n1549) );
  EN U1908 ( .A(n10159), .B(n10735), .Z(n1550) );
  EN U1909 ( .A(n10156), .B(n10735), .Z(n1551) );
  EN U1910 ( .A(n10153), .B(n10735), .Z(n1552) );
  EN U1911 ( .A(n10150), .B(n10735), .Z(n1553) );
  EN U1912 ( .A(n10147), .B(n10735), .Z(n1554) );
  EN U1913 ( .A(n10144), .B(n10735), .Z(n1555) );
  EN U1914 ( .A(n10141), .B(n10735), .Z(n1556) );
  EN U1915 ( .A(n10138), .B(n10734), .Z(n1557) );
  EN U1916 ( .A(n10135), .B(n10734), .Z(n1558) );
  EN U1917 ( .A(n10132), .B(n10734), .Z(n1559) );
  EN U1918 ( .A(n10129), .B(n10734), .Z(n1560) );
  EN U1919 ( .A(n10126), .B(n10734), .Z(n1561) );
  EN U1920 ( .A(n10123), .B(n10734), .Z(n1562) );
  EN U1921 ( .A(n10120), .B(n10734), .Z(n1563) );
  EN U1922 ( .A(n10117), .B(n10734), .Z(n1564) );
  EN U1923 ( .A(n10114), .B(n10734), .Z(n1565) );
  EN U1924 ( .A(n10111), .B(n10734), .Z(n1566) );
  EN U1925 ( .A(n10108), .B(n10734), .Z(n1567) );
  EN U1926 ( .A(n10105), .B(n10734), .Z(n1568) );
  EN U1927 ( .A(n10102), .B(n10734), .Z(n1569) );
  EN U1928 ( .A(n10099), .B(n10734), .Z(n1570) );
  EN U1929 ( .A(n10096), .B(n10733), .Z(n1571) );
  EN U1930 ( .A(n10093), .B(n10733), .Z(n1572) );
  EN U1931 ( .A(n10090), .B(n10733), .Z(n1573) );
  EN U1932 ( .A(n10087), .B(n10733), .Z(n1574) );
  EN U1933 ( .A(n10084), .B(n10733), .Z(n1575) );
  EN U1934 ( .A(n10081), .B(n10733), .Z(n1576) );
  EN U1935 ( .A(n10078), .B(n10733), .Z(n1577) );
  EN U1936 ( .A(n10075), .B(n10733), .Z(n1578) );
  EN U1937 ( .A(n10072), .B(n10733), .Z(n1579) );
  EN U1938 ( .A(n10069), .B(n10733), .Z(n1580) );
  EN U1939 ( .A(n10066), .B(n10733), .Z(n1581) );
  EN U1940 ( .A(n10063), .B(n10733), .Z(n1582) );
  EN U1941 ( .A(n10060), .B(n10733), .Z(n1583) );
  AO4 U1942 ( .A(n10413), .B(n1520), .C(n1521), .D(n10577), .Z(n3663) );
  AO4 U1943 ( .A(n10413), .B(n1521), .C(n1522), .D(n10577), .Z(n3664) );
  AO4 U1944 ( .A(n10413), .B(n1522), .C(n1523), .D(n10577), .Z(n3665) );
  AO4 U1945 ( .A(n10413), .B(n1523), .C(n1524), .D(n10577), .Z(n3666) );
  AO4 U1946 ( .A(n10413), .B(n1524), .C(n1525), .D(n10577), .Z(n3667) );
  AO4 U1947 ( .A(n10413), .B(n1525), .C(n1526), .D(n10577), .Z(n3668) );
  AO4 U1948 ( .A(n10413), .B(n1526), .C(n1527), .D(n10577), .Z(n3669) );
  AO4 U1949 ( .A(n10413), .B(n1527), .C(n1528), .D(n10577), .Z(n3670) );
  AO4 U1950 ( .A(n10413), .B(n1528), .C(n1529), .D(n10577), .Z(n3671) );
  AO4 U1951 ( .A(n10413), .B(n1529), .C(n1530), .D(n10577), .Z(n3672) );
  AO4 U1952 ( .A(n10412), .B(n1530), .C(n1531), .D(n10577), .Z(n3673) );
  AO4 U1953 ( .A(n10412), .B(n1531), .C(n1532), .D(n10576), .Z(n3674) );
  AO4 U1954 ( .A(n10412), .B(n1532), .C(n1533), .D(n10576), .Z(n3675) );
  AO4 U1955 ( .A(n10412), .B(n1533), .C(n1534), .D(n10576), .Z(n3676) );
  AO4 U1956 ( .A(n10412), .B(n1534), .C(n1535), .D(n10576), .Z(n3677) );
  AO4 U1957 ( .A(n10412), .B(n1535), .C(n1536), .D(n10576), .Z(n3678) );
  AO4 U1958 ( .A(n10412), .B(n1536), .C(n1537), .D(n10576), .Z(n3679) );
  AO4 U1959 ( .A(n10412), .B(n1537), .C(n1538), .D(n10576), .Z(n3680) );
  AO4 U1960 ( .A(n10412), .B(n1538), .C(n1539), .D(n10576), .Z(n3681) );
  AO4 U1961 ( .A(n10412), .B(n1539), .C(n1540), .D(n10576), .Z(n3682) );
  AO4 U1962 ( .A(n10412), .B(n1540), .C(n1541), .D(n10576), .Z(n3683) );
  AO4 U1963 ( .A(n10412), .B(n1541), .C(n1542), .D(n10576), .Z(n3684) );
  AO4 U1964 ( .A(n10412), .B(n1542), .C(n1543), .D(n10576), .Z(n3685) );
  AO4 U1965 ( .A(n10412), .B(n1543), .C(n1544), .D(n10576), .Z(n3686) );
  AO4 U1966 ( .A(n10411), .B(n1544), .C(n1545), .D(n10576), .Z(n3687) );
  AO4 U1967 ( .A(n10411), .B(n1545), .C(n1546), .D(n10575), .Z(n3688) );
  AO4 U1968 ( .A(n10411), .B(n1546), .C(n1547), .D(n10575), .Z(n3689) );
  AO4 U1969 ( .A(n10411), .B(n1547), .C(n1548), .D(n10575), .Z(n3690) );
  AO4 U1970 ( .A(n10411), .B(n1548), .C(n1549), .D(n10575), .Z(n3691) );
  AO4 U1971 ( .A(n10411), .B(n1549), .C(n1550), .D(n10575), .Z(n3692) );
  AO4 U1972 ( .A(n10411), .B(n1550), .C(n1551), .D(n10575), .Z(n3693) );
  AO4 U1973 ( .A(n10411), .B(n1551), .C(n1552), .D(n10575), .Z(n3694) );
  AO4 U1974 ( .A(n10411), .B(n1552), .C(n1553), .D(n10575), .Z(n3695) );
  AO4 U1975 ( .A(n10411), .B(n1553), .C(n1554), .D(n10575), .Z(n3696) );
  AO4 U1976 ( .A(n10411), .B(n1554), .C(n1555), .D(n10575), .Z(n3697) );
  AO4 U1977 ( .A(n10411), .B(n1555), .C(n1556), .D(n10575), .Z(n3698) );
  AO4 U1978 ( .A(n10411), .B(n1556), .C(n1557), .D(n10575), .Z(n3699) );
  AO4 U1979 ( .A(n10411), .B(n1557), .C(n1558), .D(n10575), .Z(n3700) );
  AO4 U1980 ( .A(n10410), .B(n1558), .C(n1559), .D(n10575), .Z(n3701) );
  AO4 U1981 ( .A(n10410), .B(n1559), .C(n1560), .D(n10574), .Z(n3702) );
  AO4 U1982 ( .A(n10410), .B(n1560), .C(n1561), .D(n10574), .Z(n3703) );
  AO4 U1983 ( .A(n10410), .B(n1561), .C(n1562), .D(n10574), .Z(n3704) );
  AO4 U1984 ( .A(n10410), .B(n1562), .C(n1563), .D(n10574), .Z(n3705) );
  AO4 U1985 ( .A(n10410), .B(n1563), .C(n1564), .D(n10574), .Z(n3706) );
  AO4 U1986 ( .A(n10410), .B(n1564), .C(n1565), .D(n10574), .Z(n3707) );
  AO4 U1987 ( .A(n10410), .B(n1565), .C(n1566), .D(n10574), .Z(n3708) );
  AO4 U1988 ( .A(n10410), .B(n1566), .C(n1567), .D(n10574), .Z(n3709) );
  AO4 U1989 ( .A(n10410), .B(n1567), .C(n1568), .D(n10574), .Z(n3710) );
  AO4 U1990 ( .A(n10410), .B(n1568), .C(n1569), .D(n10574), .Z(n3711) );
  AO4 U1991 ( .A(n10410), .B(n1569), .C(n1570), .D(n10574), .Z(n3712) );
  AO4 U1992 ( .A(n10410), .B(n1570), .C(n1571), .D(n10574), .Z(n3713) );
  AO4 U1993 ( .A(n10410), .B(n1571), .C(n1572), .D(n10574), .Z(n3714) );
  AO4 U1994 ( .A(n10409), .B(n1572), .C(n1573), .D(n10574), .Z(n3715) );
  AO4 U1995 ( .A(n10409), .B(n1573), .C(n1574), .D(n10573), .Z(n3716) );
  AO4 U1996 ( .A(n10409), .B(n1574), .C(n1575), .D(n10573), .Z(n3717) );
  AO4 U1997 ( .A(n10409), .B(n1575), .C(n1576), .D(n10573), .Z(n3718) );
  AO4 U1998 ( .A(n10409), .B(n1576), .C(n1577), .D(n10573), .Z(n3719) );
  AO4 U1999 ( .A(n10409), .B(n1577), .C(n1578), .D(n10573), .Z(n3720) );
  AO4 U2000 ( .A(n10409), .B(n1578), .C(n1579), .D(n10573), .Z(n3721) );
  AO4 U2001 ( .A(n10409), .B(n1579), .C(n1580), .D(n10573), .Z(n3722) );
  AO4 U2002 ( .A(n10409), .B(n1580), .C(n1581), .D(n10573), .Z(n3723) );
  AO4 U2003 ( .A(n10409), .B(n1581), .C(n1582), .D(n10573), .Z(n3724) );
  AO4 U2004 ( .A(n10409), .B(n1582), .C(n1583), .D(n10573), .Z(n3725) );
  AO4 U2005 ( .A(n10409), .B(n1583), .C(n1390), .D(n10573), .Z(n3726) );
  AO4 U2006 ( .A(n1519), .B(n10573), .C(n10409), .D(n1390), .Z(n5838) );
  EN U2007 ( .A(n10253), .B(n10732), .Z(n1585) );
  EN U2008 ( .A(n10246), .B(n10732), .Z(n1586) );
  EN U2009 ( .A(n10243), .B(n10732), .Z(n1587) );
  EN U2010 ( .A(n10240), .B(n10732), .Z(n1588) );
  EN U2011 ( .A(n10237), .B(n10732), .Z(n1589) );
  EN U2012 ( .A(n10234), .B(n10732), .Z(n1590) );
  EN U2013 ( .A(n10231), .B(n10732), .Z(n1591) );
  EN U2014 ( .A(n10228), .B(n10732), .Z(n1592) );
  EN U2015 ( .A(n10225), .B(n10732), .Z(n1593) );
  EN U2016 ( .A(n10222), .B(n10731), .Z(n1594) );
  EN U2017 ( .A(n10219), .B(n10731), .Z(n1595) );
  EN U2018 ( .A(n10216), .B(n10731), .Z(n1596) );
  EN U2019 ( .A(n10213), .B(n10731), .Z(n1597) );
  EN U2020 ( .A(n10210), .B(n10731), .Z(n1598) );
  EN U2021 ( .A(n10207), .B(n10731), .Z(n1599) );
  EN U2022 ( .A(n10204), .B(n10731), .Z(n1600) );
  EN U2023 ( .A(n10201), .B(n10731), .Z(n1601) );
  EN U2024 ( .A(n10198), .B(n10731), .Z(n1602) );
  EN U2025 ( .A(n10195), .B(n10731), .Z(n1603) );
  EN U2026 ( .A(n10192), .B(n10731), .Z(n1604) );
  EN U2027 ( .A(n10189), .B(n10731), .Z(n1605) );
  EN U2028 ( .A(n10186), .B(n10731), .Z(n1606) );
  EN U2029 ( .A(n10183), .B(n10731), .Z(n1607) );
  EN U2030 ( .A(n10180), .B(n10730), .Z(n1608) );
  EN U2031 ( .A(n10177), .B(n10730), .Z(n1609) );
  EN U2032 ( .A(n10174), .B(n10730), .Z(n1610) );
  EN U2033 ( .A(n10171), .B(n10730), .Z(n1611) );
  EN U2034 ( .A(n10168), .B(n10730), .Z(n1612) );
  EN U2035 ( .A(n10165), .B(n10730), .Z(n1613) );
  EN U2036 ( .A(n10162), .B(n10730), .Z(n1614) );
  EN U2037 ( .A(n10159), .B(n10730), .Z(n1615) );
  EN U2038 ( .A(n10156), .B(n10730), .Z(n1616) );
  EN U2039 ( .A(n10153), .B(n10730), .Z(n1617) );
  EN U2040 ( .A(n10150), .B(n10730), .Z(n1618) );
  EN U2041 ( .A(n10147), .B(n10730), .Z(n1619) );
  EN U2042 ( .A(n10144), .B(n10730), .Z(n1620) );
  EN U2043 ( .A(n10141), .B(n10730), .Z(n1621) );
  EN U2044 ( .A(n10138), .B(n10729), .Z(n1622) );
  EN U2045 ( .A(n10135), .B(n10729), .Z(n1623) );
  EN U2046 ( .A(n10132), .B(n10729), .Z(n1624) );
  EN U2047 ( .A(n10129), .B(n10729), .Z(n1625) );
  EN U2048 ( .A(n10126), .B(n10729), .Z(n1626) );
  EN U2049 ( .A(n10123), .B(n10729), .Z(n1627) );
  EN U2050 ( .A(n10120), .B(n10729), .Z(n1628) );
  EN U2051 ( .A(n10117), .B(n10729), .Z(n1629) );
  EN U2052 ( .A(n10114), .B(n10729), .Z(n1630) );
  EN U2053 ( .A(n10111), .B(n10729), .Z(n1631) );
  EN U2054 ( .A(n10108), .B(n10729), .Z(n1632) );
  EN U2055 ( .A(n10105), .B(n10729), .Z(n1633) );
  EN U2056 ( .A(n10102), .B(n10729), .Z(n1634) );
  EN U2057 ( .A(n10099), .B(n10729), .Z(n1635) );
  EN U2058 ( .A(n10096), .B(n10728), .Z(n1636) );
  EN U2059 ( .A(n10093), .B(n10728), .Z(n1637) );
  EN U2060 ( .A(n10090), .B(n10728), .Z(n1638) );
  EN U2061 ( .A(n10087), .B(n10728), .Z(n1639) );
  EN U2062 ( .A(n10084), .B(n10728), .Z(n1640) );
  EN U2063 ( .A(n10081), .B(n10728), .Z(n1641) );
  EN U2064 ( .A(n10078), .B(n10728), .Z(n1642) );
  EN U2065 ( .A(n10075), .B(n10728), .Z(n1643) );
  EN U2066 ( .A(n10072), .B(n10728), .Z(n1644) );
  EN U2067 ( .A(n10069), .B(n10728), .Z(n1645) );
  EN U2068 ( .A(n10066), .B(n10728), .Z(n1646) );
  EN U2069 ( .A(n10063), .B(n10728), .Z(n1647) );
  EN U2070 ( .A(n10060), .B(n10728), .Z(n1648) );
  AO4 U2071 ( .A(n10408), .B(n1585), .C(n1586), .D(n10572), .Z(n3729) );
  AO4 U2072 ( .A(n10408), .B(n1586), .C(n1587), .D(n10572), .Z(n3730) );
  AO4 U2073 ( .A(n10408), .B(n1587), .C(n1588), .D(n10572), .Z(n3731) );
  AO4 U2074 ( .A(n10408), .B(n1588), .C(n1589), .D(n10572), .Z(n3732) );
  AO4 U2075 ( .A(n10408), .B(n1589), .C(n1590), .D(n10572), .Z(n3733) );
  AO4 U2076 ( .A(n10408), .B(n1590), .C(n1591), .D(n10572), .Z(n3734) );
  AO4 U2077 ( .A(n10408), .B(n1591), .C(n1592), .D(n10572), .Z(n3735) );
  AO4 U2078 ( .A(n10408), .B(n1592), .C(n1593), .D(n10572), .Z(n3736) );
  AO4 U2079 ( .A(n10408), .B(n1593), .C(n1594), .D(n10572), .Z(n3737) );
  AO4 U2080 ( .A(n10408), .B(n1594), .C(n1595), .D(n10572), .Z(n3738) );
  AO4 U2081 ( .A(n10407), .B(n1595), .C(n1596), .D(n10572), .Z(n3739) );
  AO4 U2082 ( .A(n10407), .B(n1596), .C(n1597), .D(n10571), .Z(n3740) );
  AO4 U2083 ( .A(n10407), .B(n1597), .C(n1598), .D(n10571), .Z(n3741) );
  AO4 U2084 ( .A(n10407), .B(n1598), .C(n1599), .D(n10571), .Z(n3742) );
  AO4 U2085 ( .A(n10407), .B(n1599), .C(n1600), .D(n10571), .Z(n3743) );
  AO4 U2086 ( .A(n10407), .B(n1600), .C(n1601), .D(n10571), .Z(n3744) );
  AO4 U2087 ( .A(n10407), .B(n1601), .C(n1602), .D(n10571), .Z(n3745) );
  AO4 U2088 ( .A(n10407), .B(n1602), .C(n1603), .D(n10571), .Z(n3746) );
  AO4 U2089 ( .A(n10407), .B(n1603), .C(n1604), .D(n10571), .Z(n3747) );
  AO4 U2090 ( .A(n10407), .B(n1604), .C(n1605), .D(n10571), .Z(n3748) );
  AO4 U2091 ( .A(n10407), .B(n1605), .C(n1606), .D(n10571), .Z(n3749) );
  AO4 U2092 ( .A(n10407), .B(n1606), .C(n1607), .D(n10571), .Z(n3750) );
  AO4 U2093 ( .A(n10407), .B(n1607), .C(n1608), .D(n10571), .Z(n3751) );
  AO4 U2094 ( .A(n10407), .B(n1608), .C(n1609), .D(n10571), .Z(n3752) );
  AO4 U2095 ( .A(n10406), .B(n1609), .C(n1610), .D(n10571), .Z(n3753) );
  AO4 U2096 ( .A(n10406), .B(n1610), .C(n1611), .D(n10570), .Z(n3754) );
  AO4 U2097 ( .A(n10406), .B(n1611), .C(n1612), .D(n10570), .Z(n3755) );
  AO4 U2098 ( .A(n10406), .B(n1612), .C(n1613), .D(n10570), .Z(n3756) );
  AO4 U2099 ( .A(n10406), .B(n1613), .C(n1614), .D(n10570), .Z(n3757) );
  AO4 U2100 ( .A(n10406), .B(n1614), .C(n1615), .D(n10570), .Z(n3758) );
  AO4 U2101 ( .A(n10406), .B(n1615), .C(n1616), .D(n10570), .Z(n3759) );
  AO4 U2102 ( .A(n10406), .B(n1616), .C(n1617), .D(n10570), .Z(n3760) );
  AO4 U2103 ( .A(n10406), .B(n1617), .C(n1618), .D(n10570), .Z(n3761) );
  AO4 U2104 ( .A(n10406), .B(n1618), .C(n1619), .D(n10570), .Z(n3762) );
  AO4 U2105 ( .A(n10406), .B(n1619), .C(n1620), .D(n10570), .Z(n3763) );
  AO4 U2106 ( .A(n10406), .B(n1620), .C(n1621), .D(n10570), .Z(n3764) );
  AO4 U2107 ( .A(n10406), .B(n1621), .C(n1622), .D(n10570), .Z(n3765) );
  AO4 U2108 ( .A(n10406), .B(n1622), .C(n1623), .D(n10570), .Z(n3766) );
  AO4 U2109 ( .A(n10405), .B(n1623), .C(n1624), .D(n10570), .Z(n3767) );
  AO4 U2110 ( .A(n10405), .B(n1624), .C(n1625), .D(n10569), .Z(n3768) );
  AO4 U2111 ( .A(n10405), .B(n1625), .C(n1626), .D(n10569), .Z(n3769) );
  AO4 U2112 ( .A(n10405), .B(n1626), .C(n1627), .D(n10569), .Z(n3770) );
  AO4 U2113 ( .A(n10405), .B(n1627), .C(n1628), .D(n10569), .Z(n3771) );
  AO4 U2114 ( .A(n10405), .B(n1628), .C(n1629), .D(n10569), .Z(n3772) );
  AO4 U2115 ( .A(n10405), .B(n1629), .C(n1630), .D(n10569), .Z(n3773) );
  AO4 U2116 ( .A(n10405), .B(n1630), .C(n1631), .D(n10569), .Z(n3774) );
  AO4 U2117 ( .A(n10405), .B(n1631), .C(n1632), .D(n10569), .Z(n3775) );
  AO4 U2118 ( .A(n10405), .B(n1632), .C(n1633), .D(n10569), .Z(n3776) );
  AO4 U2119 ( .A(n10405), .B(n1633), .C(n1634), .D(n10569), .Z(n3777) );
  AO4 U2120 ( .A(n10405), .B(n1634), .C(n1635), .D(n10569), .Z(n3778) );
  AO4 U2121 ( .A(n10405), .B(n1635), .C(n1636), .D(n10569), .Z(n3779) );
  AO4 U2122 ( .A(n10405), .B(n1636), .C(n1637), .D(n10569), .Z(n3780) );
  AO4 U2123 ( .A(n10404), .B(n1637), .C(n1638), .D(n10569), .Z(n3781) );
  AO4 U2124 ( .A(n10404), .B(n1638), .C(n1639), .D(n10568), .Z(n3782) );
  AO4 U2125 ( .A(n10404), .B(n1639), .C(n1640), .D(n10568), .Z(n3783) );
  AO4 U2126 ( .A(n10404), .B(n1640), .C(n1641), .D(n10568), .Z(n3784) );
  AO4 U2127 ( .A(n10404), .B(n1641), .C(n1642), .D(n10568), .Z(n3785) );
  AO4 U2128 ( .A(n10404), .B(n1642), .C(n1643), .D(n10568), .Z(n3786) );
  AO4 U2129 ( .A(n10404), .B(n1643), .C(n1644), .D(n10568), .Z(n3787) );
  AO4 U2130 ( .A(n10404), .B(n1644), .C(n1645), .D(n10568), .Z(n3788) );
  AO4 U2131 ( .A(n10404), .B(n1645), .C(n1646), .D(n10568), .Z(n3789) );
  AO4 U2132 ( .A(n10404), .B(n1646), .C(n1647), .D(n10568), .Z(n3790) );
  AO4 U2133 ( .A(n10404), .B(n1647), .C(n1648), .D(n10568), .Z(n3791) );
  AO4 U2134 ( .A(n10404), .B(n1648), .C(n10568), .D(n1391), .Z(n3792) );
  AO4 U2135 ( .A(n10568), .B(n1584), .C(n10404), .D(n1391), .Z(n5839) );
  EN U2136 ( .A(n10253), .B(n10727), .Z(n1650) );
  EN U2137 ( .A(n10246), .B(n10727), .Z(n1651) );
  EN U2138 ( .A(n10243), .B(n10727), .Z(n1652) );
  EN U2139 ( .A(n10240), .B(n10727), .Z(n1653) );
  EN U2140 ( .A(n10237), .B(n10727), .Z(n1654) );
  EN U2141 ( .A(n10234), .B(n10727), .Z(n1655) );
  EN U2142 ( .A(n10231), .B(n10727), .Z(n1656) );
  EN U2143 ( .A(n10228), .B(n10727), .Z(n1657) );
  EN U2144 ( .A(n10225), .B(n10727), .Z(n1658) );
  EN U2145 ( .A(n10222), .B(n10726), .Z(n1659) );
  EN U2146 ( .A(n10219), .B(n10726), .Z(n1660) );
  EN U2147 ( .A(n10216), .B(n10726), .Z(n1661) );
  EN U2148 ( .A(n10213), .B(n10726), .Z(n1662) );
  EN U2149 ( .A(n10210), .B(n10726), .Z(n1663) );
  EN U2150 ( .A(n10207), .B(n10726), .Z(n1664) );
  EN U2151 ( .A(n10204), .B(n10726), .Z(n1665) );
  EN U2152 ( .A(n10201), .B(n10726), .Z(n1666) );
  EN U2153 ( .A(n10198), .B(n10726), .Z(n1667) );
  EN U2154 ( .A(n10195), .B(n10726), .Z(n1668) );
  EN U2155 ( .A(n10192), .B(n10726), .Z(n1669) );
  EN U2156 ( .A(n10189), .B(n10726), .Z(n1670) );
  EN U2157 ( .A(n10186), .B(n10726), .Z(n1671) );
  EN U2158 ( .A(n10183), .B(n10726), .Z(n1672) );
  EN U2159 ( .A(n10180), .B(n10725), .Z(n1673) );
  EN U2160 ( .A(n10177), .B(n10725), .Z(n1674) );
  EN U2161 ( .A(n10174), .B(n10725), .Z(n1675) );
  EN U2162 ( .A(n10171), .B(n10725), .Z(n1676) );
  EN U2163 ( .A(n10168), .B(n10725), .Z(n1677) );
  EN U2164 ( .A(n10165), .B(n10725), .Z(n1678) );
  EN U2165 ( .A(n10162), .B(n10725), .Z(n1679) );
  EN U2166 ( .A(n10159), .B(n10725), .Z(n1680) );
  EN U2167 ( .A(n10156), .B(n10725), .Z(n1681) );
  EN U2168 ( .A(n10153), .B(n10725), .Z(n1682) );
  EN U2169 ( .A(n10150), .B(n10725), .Z(n1683) );
  EN U2170 ( .A(n10147), .B(n10725), .Z(n1684) );
  EN U2171 ( .A(n10144), .B(n10725), .Z(n1685) );
  EN U2172 ( .A(n10141), .B(n10725), .Z(n1686) );
  EN U2173 ( .A(n10138), .B(n10724), .Z(n1687) );
  EN U2174 ( .A(n10135), .B(n10724), .Z(n1688) );
  EN U2175 ( .A(n10132), .B(n10724), .Z(n1689) );
  EN U2176 ( .A(n10129), .B(n10724), .Z(n1690) );
  EN U2177 ( .A(n10126), .B(n10724), .Z(n1691) );
  EN U2178 ( .A(n10123), .B(n10724), .Z(n1692) );
  EN U2179 ( .A(n10120), .B(n10724), .Z(n1693) );
  EN U2180 ( .A(n10117), .B(n10724), .Z(n1694) );
  EN U2181 ( .A(n10114), .B(n10724), .Z(n1695) );
  EN U2182 ( .A(n10111), .B(n10724), .Z(n1696) );
  EN U2183 ( .A(n10108), .B(n10724), .Z(n1697) );
  EN U2184 ( .A(n10105), .B(n10724), .Z(n1698) );
  EN U2185 ( .A(n10102), .B(n10724), .Z(n1699) );
  EN U2186 ( .A(n10099), .B(n10724), .Z(n1700) );
  EN U2187 ( .A(n10096), .B(n10723), .Z(n1701) );
  EN U2188 ( .A(n10093), .B(n10723), .Z(n1702) );
  EN U2189 ( .A(n10090), .B(n10723), .Z(n1703) );
  EN U2190 ( .A(n10087), .B(n10723), .Z(n1704) );
  EN U2191 ( .A(n10084), .B(n10723), .Z(n1705) );
  EN U2192 ( .A(n10081), .B(n10723), .Z(n1706) );
  EN U2193 ( .A(n10078), .B(n10723), .Z(n1707) );
  EN U2194 ( .A(n10075), .B(n10723), .Z(n1708) );
  EN U2195 ( .A(n10072), .B(n10723), .Z(n1709) );
  EN U2196 ( .A(n10069), .B(n10723), .Z(n1710) );
  EN U2197 ( .A(n10066), .B(n10723), .Z(n1711) );
  EN U2198 ( .A(n10063), .B(n10723), .Z(n1712) );
  EN U2199 ( .A(n10060), .B(n10723), .Z(n1713) );
  AO4 U2200 ( .A(n10403), .B(n1650), .C(n1651), .D(n10567), .Z(n3795) );
  AO4 U2201 ( .A(n10403), .B(n1651), .C(n1652), .D(n10567), .Z(n3796) );
  AO4 U2202 ( .A(n10403), .B(n1652), .C(n1653), .D(n10567), .Z(n3797) );
  AO4 U2203 ( .A(n10403), .B(n1653), .C(n1654), .D(n10567), .Z(n3798) );
  AO4 U2204 ( .A(n10403), .B(n1654), .C(n1655), .D(n10567), .Z(n3799) );
  AO4 U2205 ( .A(n10403), .B(n1655), .C(n1656), .D(n10567), .Z(n3800) );
  AO4 U2206 ( .A(n10403), .B(n1656), .C(n1657), .D(n10567), .Z(n3801) );
  AO4 U2207 ( .A(n10403), .B(n1657), .C(n1658), .D(n10567), .Z(n3802) );
  AO4 U2208 ( .A(n10403), .B(n1658), .C(n1659), .D(n10567), .Z(n3803) );
  AO4 U2209 ( .A(n10403), .B(n1659), .C(n1660), .D(n10567), .Z(n3804) );
  AO4 U2210 ( .A(n10402), .B(n1660), .C(n1661), .D(n10567), .Z(n3805) );
  AO4 U2211 ( .A(n10402), .B(n1661), .C(n1662), .D(n10566), .Z(n3806) );
  AO4 U2212 ( .A(n10402), .B(n1662), .C(n1663), .D(n10566), .Z(n3807) );
  AO4 U2213 ( .A(n10402), .B(n1663), .C(n1664), .D(n10566), .Z(n3808) );
  AO4 U2214 ( .A(n10402), .B(n1664), .C(n1665), .D(n10566), .Z(n3809) );
  AO4 U2215 ( .A(n10402), .B(n1665), .C(n1666), .D(n10566), .Z(n3810) );
  AO4 U2216 ( .A(n10402), .B(n1666), .C(n1667), .D(n10566), .Z(n3811) );
  AO4 U2217 ( .A(n10402), .B(n1667), .C(n1668), .D(n10566), .Z(n3812) );
  AO4 U2218 ( .A(n10402), .B(n1668), .C(n1669), .D(n10566), .Z(n3813) );
  AO4 U2219 ( .A(n10402), .B(n1669), .C(n1670), .D(n10566), .Z(n3814) );
  AO4 U2220 ( .A(n10402), .B(n1670), .C(n1671), .D(n10566), .Z(n3815) );
  AO4 U2221 ( .A(n10402), .B(n1671), .C(n1672), .D(n10566), .Z(n3816) );
  AO4 U2222 ( .A(n10402), .B(n1672), .C(n1673), .D(n10566), .Z(n3817) );
  AO4 U2223 ( .A(n10402), .B(n1673), .C(n1674), .D(n10566), .Z(n3818) );
  AO4 U2224 ( .A(n10401), .B(n1674), .C(n1675), .D(n10566), .Z(n3819) );
  AO4 U2225 ( .A(n10401), .B(n1675), .C(n1676), .D(n10565), .Z(n3820) );
  AO4 U2226 ( .A(n10401), .B(n1676), .C(n1677), .D(n10565), .Z(n3821) );
  AO4 U2227 ( .A(n10401), .B(n1677), .C(n1678), .D(n10565), .Z(n3822) );
  AO4 U2228 ( .A(n10401), .B(n1678), .C(n1679), .D(n10565), .Z(n3823) );
  AO4 U2229 ( .A(n10401), .B(n1679), .C(n1680), .D(n10565), .Z(n3824) );
  AO4 U2230 ( .A(n10401), .B(n1680), .C(n1681), .D(n10565), .Z(n3825) );
  AO4 U2231 ( .A(n10401), .B(n1681), .C(n1682), .D(n10565), .Z(n3826) );
  AO4 U2232 ( .A(n10401), .B(n1682), .C(n1683), .D(n10565), .Z(n3827) );
  AO4 U2233 ( .A(n10401), .B(n1683), .C(n1684), .D(n10565), .Z(n3828) );
  AO4 U2234 ( .A(n10401), .B(n1684), .C(n1685), .D(n10565), .Z(n3829) );
  AO4 U2235 ( .A(n10401), .B(n1685), .C(n1686), .D(n10565), .Z(n3830) );
  AO4 U2236 ( .A(n10401), .B(n1686), .C(n1687), .D(n10565), .Z(n3831) );
  AO4 U2237 ( .A(n10401), .B(n1687), .C(n1688), .D(n10565), .Z(n3832) );
  AO4 U2238 ( .A(n10400), .B(n1688), .C(n1689), .D(n10565), .Z(n3833) );
  AO4 U2239 ( .A(n10400), .B(n1689), .C(n1690), .D(n10564), .Z(n3834) );
  AO4 U2240 ( .A(n10400), .B(n1690), .C(n1691), .D(n10564), .Z(n3835) );
  AO4 U2241 ( .A(n10400), .B(n1691), .C(n1692), .D(n10564), .Z(n3836) );
  AO4 U2242 ( .A(n10400), .B(n1692), .C(n1693), .D(n10564), .Z(n3837) );
  AO4 U2243 ( .A(n10400), .B(n1693), .C(n1694), .D(n10564), .Z(n3838) );
  AO4 U2244 ( .A(n10400), .B(n1694), .C(n1695), .D(n10564), .Z(n3839) );
  AO4 U2245 ( .A(n10400), .B(n1695), .C(n1696), .D(n10564), .Z(n3840) );
  AO4 U2246 ( .A(n10400), .B(n1696), .C(n1697), .D(n10564), .Z(n3841) );
  AO4 U2247 ( .A(n10400), .B(n1697), .C(n1698), .D(n10564), .Z(n3842) );
  AO4 U2248 ( .A(n10400), .B(n1698), .C(n1699), .D(n10564), .Z(n3843) );
  AO4 U2249 ( .A(n10400), .B(n1699), .C(n1700), .D(n10564), .Z(n3844) );
  AO4 U2250 ( .A(n10400), .B(n1700), .C(n1701), .D(n10564), .Z(n3845) );
  AO4 U2251 ( .A(n10400), .B(n1701), .C(n1702), .D(n10564), .Z(n3846) );
  AO4 U2252 ( .A(n10399), .B(n1702), .C(n1703), .D(n10564), .Z(n3847) );
  AO4 U2253 ( .A(n10399), .B(n1703), .C(n1704), .D(n10563), .Z(n3848) );
  AO4 U2254 ( .A(n10399), .B(n1704), .C(n1705), .D(n10563), .Z(n3849) );
  AO4 U2255 ( .A(n10399), .B(n1705), .C(n1706), .D(n10563), .Z(n3850) );
  AO4 U2256 ( .A(n10399), .B(n1706), .C(n1707), .D(n10563), .Z(n3851) );
  AO4 U2257 ( .A(n10399), .B(n1707), .C(n1708), .D(n10563), .Z(n3852) );
  AO4 U2258 ( .A(n10399), .B(n1708), .C(n1709), .D(n10563), .Z(n3853) );
  AO4 U2259 ( .A(n10399), .B(n1709), .C(n1710), .D(n10563), .Z(n3854) );
  AO4 U2260 ( .A(n10399), .B(n1710), .C(n1711), .D(n10563), .Z(n3855) );
  AO4 U2261 ( .A(n10399), .B(n1711), .C(n1712), .D(n10563), .Z(n3856) );
  AO4 U2262 ( .A(n10399), .B(n1712), .C(n1713), .D(n10563), .Z(n3857) );
  AO4 U2263 ( .A(n10399), .B(n1713), .C(n10563), .D(n1392), .Z(n3858) );
  AO4 U2264 ( .A(n10563), .B(n1649), .C(n10399), .D(n1392), .Z(n5840) );
  EN U2265 ( .A(n10253), .B(n10722), .Z(n1715) );
  EN U2266 ( .A(n10246), .B(n10722), .Z(n1716) );
  EN U2267 ( .A(n10243), .B(n10722), .Z(n1717) );
  EN U2268 ( .A(n10240), .B(n10722), .Z(n1718) );
  EN U2269 ( .A(n10237), .B(n10722), .Z(n1719) );
  EN U2270 ( .A(n10234), .B(n10722), .Z(n1720) );
  EN U2271 ( .A(n10231), .B(n10722), .Z(n1721) );
  EN U2272 ( .A(n10228), .B(n10722), .Z(n1722) );
  EN U2273 ( .A(n10225), .B(n10722), .Z(n1723) );
  EN U2274 ( .A(n10222), .B(n10721), .Z(n1724) );
  EN U2275 ( .A(n10219), .B(n10721), .Z(n1725) );
  EN U2276 ( .A(n10216), .B(n10721), .Z(n1726) );
  EN U2277 ( .A(n10213), .B(n10721), .Z(n1727) );
  EN U2278 ( .A(n10210), .B(n10721), .Z(n1728) );
  EN U2279 ( .A(n10207), .B(n10721), .Z(n1729) );
  EN U2280 ( .A(n10204), .B(n10721), .Z(n1730) );
  EN U2281 ( .A(n10201), .B(n10721), .Z(n1731) );
  EN U2282 ( .A(n10198), .B(n10721), .Z(n1732) );
  EN U2283 ( .A(n10195), .B(n10721), .Z(n1733) );
  EN U2284 ( .A(n10192), .B(n10721), .Z(n1734) );
  EN U2285 ( .A(n10189), .B(n10721), .Z(n1735) );
  EN U2286 ( .A(n10186), .B(n10721), .Z(n1736) );
  EN U2287 ( .A(n10183), .B(n10721), .Z(n1737) );
  EN U2288 ( .A(n10180), .B(n10720), .Z(n1738) );
  EN U2289 ( .A(n10177), .B(n10720), .Z(n1739) );
  EN U2290 ( .A(n10174), .B(n10720), .Z(n1740) );
  EN U2291 ( .A(n10171), .B(n10720), .Z(n1741) );
  EN U2292 ( .A(n10168), .B(n10720), .Z(n1742) );
  EN U2293 ( .A(n10165), .B(n10720), .Z(n1743) );
  EN U2294 ( .A(n10162), .B(n10720), .Z(n1744) );
  EN U2295 ( .A(n10159), .B(n10720), .Z(n1745) );
  EN U2296 ( .A(n10156), .B(n10720), .Z(n1746) );
  EN U2297 ( .A(n10153), .B(n10720), .Z(n1747) );
  EN U2298 ( .A(n10150), .B(n10720), .Z(n1748) );
  EN U2299 ( .A(n10147), .B(n10720), .Z(n1749) );
  EN U2300 ( .A(n10144), .B(n10720), .Z(n1750) );
  EN U2301 ( .A(n10141), .B(n10720), .Z(n1751) );
  EN U2302 ( .A(n10138), .B(n10719), .Z(n1752) );
  EN U2303 ( .A(n10135), .B(n10719), .Z(n1753) );
  EN U2304 ( .A(n10132), .B(n10719), .Z(n1754) );
  EN U2305 ( .A(n10129), .B(n10719), .Z(n1755) );
  EN U2306 ( .A(n10126), .B(n10719), .Z(n1756) );
  EN U2307 ( .A(n10123), .B(n10719), .Z(n1757) );
  EN U2308 ( .A(n10120), .B(n10719), .Z(n1758) );
  EN U2309 ( .A(n10117), .B(n10719), .Z(n1759) );
  EN U2310 ( .A(n10114), .B(n10719), .Z(n1760) );
  EN U2311 ( .A(n10111), .B(n10719), .Z(n1761) );
  EN U2312 ( .A(n10108), .B(n10719), .Z(n1762) );
  EN U2313 ( .A(n10105), .B(n10719), .Z(n1763) );
  EN U2314 ( .A(n10102), .B(n10719), .Z(n1764) );
  EN U2315 ( .A(n10099), .B(n10719), .Z(n1765) );
  EN U2316 ( .A(n10096), .B(n10718), .Z(n1766) );
  EN U2317 ( .A(n10093), .B(n10718), .Z(n1767) );
  EN U2318 ( .A(n10090), .B(n10718), .Z(n1768) );
  EN U2319 ( .A(n10087), .B(n10718), .Z(n1769) );
  EN U2320 ( .A(n10084), .B(n10718), .Z(n1770) );
  EN U2321 ( .A(n10081), .B(n10718), .Z(n1771) );
  EN U2322 ( .A(n10078), .B(n10718), .Z(n1772) );
  EN U2323 ( .A(n10075), .B(n10718), .Z(n1773) );
  EN U2324 ( .A(n10072), .B(n10718), .Z(n1774) );
  EN U2325 ( .A(n10069), .B(n10718), .Z(n1775) );
  EN U2326 ( .A(n10066), .B(n10718), .Z(n1776) );
  EN U2327 ( .A(n10063), .B(n10718), .Z(n1777) );
  EN U2328 ( .A(n10060), .B(n10718), .Z(n1778) );
  AO4 U2329 ( .A(n10398), .B(n1715), .C(n1716), .D(n10562), .Z(n3861) );
  AO4 U2330 ( .A(n10398), .B(n1716), .C(n1717), .D(n10562), .Z(n3862) );
  AO4 U2331 ( .A(n10398), .B(n1717), .C(n1718), .D(n10562), .Z(n3863) );
  AO4 U2332 ( .A(n10398), .B(n1718), .C(n1719), .D(n10562), .Z(n3864) );
  AO4 U2333 ( .A(n10398), .B(n1719), .C(n1720), .D(n10562), .Z(n3865) );
  AO4 U2334 ( .A(n10398), .B(n1720), .C(n1721), .D(n10562), .Z(n3866) );
  AO4 U2335 ( .A(n10398), .B(n1721), .C(n1722), .D(n10562), .Z(n3867) );
  AO4 U2336 ( .A(n10398), .B(n1722), .C(n1723), .D(n10562), .Z(n3868) );
  AO4 U2337 ( .A(n10398), .B(n1723), .C(n1724), .D(n10562), .Z(n3869) );
  AO4 U2338 ( .A(n10398), .B(n1724), .C(n1725), .D(n10562), .Z(n3870) );
  AO4 U2339 ( .A(n10397), .B(n1725), .C(n1726), .D(n10562), .Z(n3871) );
  AO4 U2340 ( .A(n10397), .B(n1726), .C(n1727), .D(n10561), .Z(n3872) );
  AO4 U2341 ( .A(n10397), .B(n1727), .C(n1728), .D(n10561), .Z(n3873) );
  AO4 U2342 ( .A(n10397), .B(n1728), .C(n1729), .D(n10561), .Z(n3874) );
  AO4 U2343 ( .A(n10397), .B(n1729), .C(n1730), .D(n10561), .Z(n3875) );
  AO4 U2344 ( .A(n10397), .B(n1730), .C(n1731), .D(n10561), .Z(n3876) );
  AO4 U2345 ( .A(n10397), .B(n1731), .C(n1732), .D(n10561), .Z(n3877) );
  AO4 U2346 ( .A(n10397), .B(n1732), .C(n1733), .D(n10561), .Z(n3878) );
  AO4 U2347 ( .A(n10397), .B(n1733), .C(n1734), .D(n10561), .Z(n3879) );
  AO4 U2348 ( .A(n10397), .B(n1734), .C(n1735), .D(n10561), .Z(n3880) );
  AO4 U2349 ( .A(n10397), .B(n1735), .C(n1736), .D(n10561), .Z(n3881) );
  AO4 U2350 ( .A(n10397), .B(n1736), .C(n1737), .D(n10561), .Z(n3882) );
  AO4 U2351 ( .A(n10397), .B(n1737), .C(n1738), .D(n10561), .Z(n3883) );
  AO4 U2352 ( .A(n10397), .B(n1738), .C(n1739), .D(n10561), .Z(n3884) );
  AO4 U2353 ( .A(n10396), .B(n1739), .C(n1740), .D(n10561), .Z(n3885) );
  AO4 U2354 ( .A(n10396), .B(n1740), .C(n1741), .D(n10560), .Z(n3886) );
  AO4 U2355 ( .A(n10396), .B(n1741), .C(n1742), .D(n10560), .Z(n3887) );
  AO4 U2356 ( .A(n10396), .B(n1742), .C(n1743), .D(n10560), .Z(n3888) );
  AO4 U2357 ( .A(n10396), .B(n1743), .C(n1744), .D(n10560), .Z(n3889) );
  AO4 U2358 ( .A(n10396), .B(n1744), .C(n1745), .D(n10560), .Z(n3890) );
  AO4 U2359 ( .A(n10396), .B(n1745), .C(n1746), .D(n10560), .Z(n3891) );
  AO4 U2360 ( .A(n10396), .B(n1746), .C(n1747), .D(n10560), .Z(n3892) );
  AO4 U2361 ( .A(n10396), .B(n1747), .C(n1748), .D(n10560), .Z(n3893) );
  AO4 U2362 ( .A(n10396), .B(n1748), .C(n1749), .D(n10560), .Z(n3894) );
  AO4 U2363 ( .A(n10396), .B(n1749), .C(n1750), .D(n10560), .Z(n3895) );
  AO4 U2364 ( .A(n10396), .B(n1750), .C(n1751), .D(n10560), .Z(n3896) );
  AO4 U2365 ( .A(n10396), .B(n1751), .C(n1752), .D(n10560), .Z(n3897) );
  AO4 U2366 ( .A(n10396), .B(n1752), .C(n1753), .D(n10560), .Z(n3898) );
  AO4 U2367 ( .A(n10395), .B(n1753), .C(n1754), .D(n10560), .Z(n3899) );
  AO4 U2368 ( .A(n10395), .B(n1754), .C(n1755), .D(n10559), .Z(n3900) );
  AO4 U2369 ( .A(n10395), .B(n1755), .C(n1756), .D(n10559), .Z(n3901) );
  AO4 U2370 ( .A(n10395), .B(n1756), .C(n1757), .D(n10559), .Z(n3902) );
  AO4 U2371 ( .A(n10395), .B(n1757), .C(n1758), .D(n10559), .Z(n3903) );
  AO4 U2372 ( .A(n10395), .B(n1758), .C(n1759), .D(n10559), .Z(n3904) );
  AO4 U2373 ( .A(n10395), .B(n1759), .C(n1760), .D(n10559), .Z(n3905) );
  AO4 U2374 ( .A(n10395), .B(n1760), .C(n1761), .D(n10559), .Z(n3906) );
  AO4 U2375 ( .A(n10395), .B(n1761), .C(n1762), .D(n10559), .Z(n3907) );
  AO4 U2376 ( .A(n10395), .B(n1762), .C(n1763), .D(n10559), .Z(n3908) );
  AO4 U2377 ( .A(n10395), .B(n1763), .C(n1764), .D(n10559), .Z(n3909) );
  AO4 U2378 ( .A(n10395), .B(n1764), .C(n1765), .D(n10559), .Z(n3910) );
  AO4 U2379 ( .A(n10395), .B(n1765), .C(n1766), .D(n10559), .Z(n3911) );
  AO4 U2380 ( .A(n10395), .B(n1766), .C(n1767), .D(n10559), .Z(n3912) );
  AO4 U2381 ( .A(n10394), .B(n1767), .C(n1768), .D(n10559), .Z(n3913) );
  AO4 U2382 ( .A(n10394), .B(n1768), .C(n1769), .D(n10558), .Z(n3914) );
  AO4 U2383 ( .A(n10394), .B(n1769), .C(n1770), .D(n10558), .Z(n3915) );
  AO4 U2384 ( .A(n10394), .B(n1770), .C(n1771), .D(n10558), .Z(n3916) );
  AO4 U2385 ( .A(n10394), .B(n1771), .C(n1772), .D(n10558), .Z(n3917) );
  AO4 U2386 ( .A(n10394), .B(n1772), .C(n1773), .D(n10558), .Z(n3918) );
  AO4 U2387 ( .A(n10394), .B(n1773), .C(n1774), .D(n10558), .Z(n3919) );
  AO4 U2388 ( .A(n10394), .B(n1774), .C(n1775), .D(n10558), .Z(n3920) );
  AO4 U2389 ( .A(n10394), .B(n1775), .C(n1776), .D(n10558), .Z(n3921) );
  AO4 U2390 ( .A(n10394), .B(n1776), .C(n1777), .D(n10558), .Z(n3922) );
  AO4 U2391 ( .A(n10394), .B(n1777), .C(n1778), .D(n10558), .Z(n3923) );
  AO4 U2392 ( .A(n10394), .B(n1778), .C(n10558), .D(n1393), .Z(n3924) );
  AO4 U2393 ( .A(n10558), .B(n1714), .C(n10394), .D(n1393), .Z(n5841) );
  EN U2394 ( .A(n10253), .B(n10717), .Z(n1780) );
  EN U2395 ( .A(n10246), .B(n10717), .Z(n1781) );
  EN U2396 ( .A(n10243), .B(n10717), .Z(n1782) );
  EN U2397 ( .A(n10240), .B(n10717), .Z(n1783) );
  EN U2398 ( .A(n10237), .B(n10717), .Z(n1784) );
  EN U2399 ( .A(n10234), .B(n10717), .Z(n1785) );
  EN U2400 ( .A(n10231), .B(n10717), .Z(n1786) );
  EN U2401 ( .A(n10228), .B(n10717), .Z(n1787) );
  EN U2402 ( .A(n10225), .B(n10717), .Z(n1788) );
  EN U2403 ( .A(n10222), .B(n10716), .Z(n1789) );
  EN U2404 ( .A(n10219), .B(n10716), .Z(n1790) );
  EN U2405 ( .A(n10216), .B(n10716), .Z(n1791) );
  EN U2406 ( .A(n10213), .B(n10716), .Z(n1792) );
  EN U2407 ( .A(n10210), .B(n10716), .Z(n1793) );
  EN U2408 ( .A(n10207), .B(n10716), .Z(n1794) );
  EN U2409 ( .A(n10204), .B(n10716), .Z(n1795) );
  EN U2410 ( .A(n10201), .B(n10716), .Z(n1796) );
  EN U2411 ( .A(n10198), .B(n10716), .Z(n1797) );
  EN U2412 ( .A(n10195), .B(n10716), .Z(n1798) );
  EN U2413 ( .A(n10192), .B(n10716), .Z(n1799) );
  EN U2414 ( .A(n10189), .B(n10716), .Z(n1800) );
  EN U2415 ( .A(n10186), .B(n10716), .Z(n1801) );
  EN U2416 ( .A(n10183), .B(n10716), .Z(n1802) );
  EN U2417 ( .A(n10180), .B(n10715), .Z(n1803) );
  EN U2418 ( .A(n10177), .B(n10715), .Z(n1804) );
  EN U2419 ( .A(n10174), .B(n10715), .Z(n1805) );
  EN U2420 ( .A(n10171), .B(n10715), .Z(n1806) );
  EN U2421 ( .A(n10168), .B(n10715), .Z(n1807) );
  EN U2422 ( .A(n10165), .B(n10715), .Z(n1808) );
  EN U2423 ( .A(n10162), .B(n10715), .Z(n1809) );
  EN U2424 ( .A(n10159), .B(n10715), .Z(n1810) );
  EN U2425 ( .A(n10156), .B(n10715), .Z(n1811) );
  EN U2426 ( .A(n10153), .B(n10715), .Z(n1812) );
  EN U2427 ( .A(n10150), .B(n10715), .Z(n1813) );
  EN U2428 ( .A(n10147), .B(n10715), .Z(n1814) );
  EN U2429 ( .A(n10144), .B(n10715), .Z(n1815) );
  EN U2430 ( .A(n10141), .B(n10715), .Z(n1816) );
  EN U2431 ( .A(n10138), .B(n10714), .Z(n1817) );
  EN U2432 ( .A(n10135), .B(n10714), .Z(n1818) );
  EN U2433 ( .A(n10132), .B(n10714), .Z(n1819) );
  EN U2434 ( .A(n10129), .B(n10714), .Z(n1820) );
  EN U2435 ( .A(n10126), .B(n10714), .Z(n1821) );
  EN U2436 ( .A(n10123), .B(n10714), .Z(n1822) );
  EN U2437 ( .A(n10120), .B(n10714), .Z(n1823) );
  EN U2438 ( .A(n10117), .B(n10714), .Z(n1824) );
  EN U2439 ( .A(n10114), .B(n10714), .Z(n1825) );
  EN U2440 ( .A(n10111), .B(n10714), .Z(n1826) );
  EN U2441 ( .A(n10108), .B(n10714), .Z(n1827) );
  EN U2442 ( .A(n10105), .B(n10714), .Z(n1828) );
  EN U2443 ( .A(n10102), .B(n10714), .Z(n1829) );
  EN U2444 ( .A(n10099), .B(n10714), .Z(n1830) );
  EN U2445 ( .A(n10096), .B(n10713), .Z(n1831) );
  EN U2446 ( .A(n10093), .B(n10713), .Z(n1832) );
  EN U2447 ( .A(n10090), .B(n10713), .Z(n1833) );
  EN U2448 ( .A(n10087), .B(n10713), .Z(n1834) );
  EN U2449 ( .A(n10084), .B(n10713), .Z(n1835) );
  EN U2450 ( .A(n10081), .B(n10713), .Z(n1836) );
  EN U2451 ( .A(n10078), .B(n10713), .Z(n1837) );
  EN U2452 ( .A(n10075), .B(n10713), .Z(n1838) );
  EN U2453 ( .A(n10072), .B(n10713), .Z(n1839) );
  EN U2454 ( .A(n10069), .B(n10713), .Z(n1840) );
  EN U2455 ( .A(n10066), .B(n10713), .Z(n1841) );
  EN U2456 ( .A(n10063), .B(n10713), .Z(n1842) );
  EN U2457 ( .A(n10060), .B(n10713), .Z(n1843) );
  AO4 U2458 ( .A(n10393), .B(n1780), .C(n1781), .D(n10557), .Z(n3927) );
  AO4 U2459 ( .A(n10393), .B(n1781), .C(n1782), .D(n10557), .Z(n3928) );
  AO4 U2460 ( .A(n10393), .B(n1782), .C(n1783), .D(n10557), .Z(n3929) );
  AO4 U2461 ( .A(n10393), .B(n1783), .C(n1784), .D(n10557), .Z(n3930) );
  AO4 U2462 ( .A(n10393), .B(n1784), .C(n1785), .D(n10557), .Z(n3931) );
  AO4 U2463 ( .A(n10393), .B(n1785), .C(n1786), .D(n10557), .Z(n3932) );
  AO4 U2464 ( .A(n10393), .B(n1786), .C(n1787), .D(n10557), .Z(n3933) );
  AO4 U2465 ( .A(n10393), .B(n1787), .C(n1788), .D(n10557), .Z(n3934) );
  AO4 U2466 ( .A(n10393), .B(n1788), .C(n1789), .D(n10557), .Z(n3935) );
  AO4 U2467 ( .A(n10393), .B(n1789), .C(n1790), .D(n10557), .Z(n3936) );
  AO4 U2468 ( .A(n10392), .B(n1790), .C(n1791), .D(n10557), .Z(n3937) );
  AO4 U2469 ( .A(n10392), .B(n1791), .C(n1792), .D(n10556), .Z(n3938) );
  AO4 U2470 ( .A(n10392), .B(n1792), .C(n1793), .D(n10556), .Z(n3939) );
  AO4 U2471 ( .A(n10392), .B(n1793), .C(n1794), .D(n10556), .Z(n3940) );
  AO4 U2472 ( .A(n10392), .B(n1794), .C(n1795), .D(n10556), .Z(n3941) );
  AO4 U2473 ( .A(n10392), .B(n1795), .C(n1796), .D(n10556), .Z(n3942) );
  AO4 U2474 ( .A(n10392), .B(n1796), .C(n1797), .D(n10556), .Z(n3943) );
  AO4 U2475 ( .A(n10392), .B(n1797), .C(n1798), .D(n10556), .Z(n3944) );
  AO4 U2476 ( .A(n10392), .B(n1798), .C(n1799), .D(n10556), .Z(n3945) );
  AO4 U2477 ( .A(n10392), .B(n1799), .C(n1800), .D(n10556), .Z(n3946) );
  AO4 U2478 ( .A(n10392), .B(n1800), .C(n1801), .D(n10556), .Z(n3947) );
  AO4 U2479 ( .A(n10392), .B(n1801), .C(n1802), .D(n10556), .Z(n3948) );
  AO4 U2480 ( .A(n10392), .B(n1802), .C(n1803), .D(n10556), .Z(n3949) );
  AO4 U2481 ( .A(n10392), .B(n1803), .C(n1804), .D(n10556), .Z(n3950) );
  AO4 U2482 ( .A(n10391), .B(n1804), .C(n1805), .D(n10556), .Z(n3951) );
  AO4 U2483 ( .A(n10391), .B(n1805), .C(n1806), .D(n10555), .Z(n3952) );
  AO4 U2484 ( .A(n10391), .B(n1806), .C(n1807), .D(n10555), .Z(n3953) );
  AO4 U2485 ( .A(n10391), .B(n1807), .C(n1808), .D(n10555), .Z(n3954) );
  AO4 U2486 ( .A(n10391), .B(n1808), .C(n1809), .D(n10555), .Z(n3955) );
  AO4 U2487 ( .A(n10391), .B(n1809), .C(n1810), .D(n10555), .Z(n3956) );
  AO4 U2488 ( .A(n10391), .B(n1810), .C(n1811), .D(n10555), .Z(n3957) );
  AO4 U2489 ( .A(n10391), .B(n1811), .C(n1812), .D(n10555), .Z(n3958) );
  AO4 U2490 ( .A(n10391), .B(n1812), .C(n1813), .D(n10555), .Z(n3959) );
  AO4 U2491 ( .A(n10391), .B(n1813), .C(n1814), .D(n10555), .Z(n3960) );
  AO4 U2492 ( .A(n10391), .B(n1814), .C(n1815), .D(n10555), .Z(n3961) );
  AO4 U2493 ( .A(n10391), .B(n1815), .C(n1816), .D(n10555), .Z(n3962) );
  AO4 U2494 ( .A(n10391), .B(n1816), .C(n1817), .D(n10555), .Z(n3963) );
  AO4 U2495 ( .A(n10391), .B(n1817), .C(n1818), .D(n10555), .Z(n3964) );
  AO4 U2496 ( .A(n10390), .B(n1818), .C(n1819), .D(n10555), .Z(n3965) );
  AO4 U2497 ( .A(n10390), .B(n1819), .C(n1820), .D(n10554), .Z(n3966) );
  AO4 U2498 ( .A(n10390), .B(n1820), .C(n1821), .D(n10554), .Z(n3967) );
  AO4 U2499 ( .A(n10390), .B(n1821), .C(n1822), .D(n10554), .Z(n3968) );
  AO4 U2500 ( .A(n10390), .B(n1822), .C(n1823), .D(n10554), .Z(n3969) );
  AO4 U2501 ( .A(n10390), .B(n1823), .C(n1824), .D(n10554), .Z(n3970) );
  AO4 U2502 ( .A(n10390), .B(n1824), .C(n1825), .D(n10554), .Z(n3971) );
  AO4 U2503 ( .A(n10390), .B(n1825), .C(n1826), .D(n10554), .Z(n3972) );
  AO4 U2504 ( .A(n10390), .B(n1826), .C(n1827), .D(n10554), .Z(n3973) );
  AO4 U2505 ( .A(n10390), .B(n1827), .C(n1828), .D(n10554), .Z(n3974) );
  AO4 U2506 ( .A(n10390), .B(n1828), .C(n1829), .D(n10554), .Z(n3975) );
  AO4 U2507 ( .A(n10390), .B(n1829), .C(n1830), .D(n10554), .Z(n3976) );
  AO4 U2508 ( .A(n10390), .B(n1830), .C(n1831), .D(n10554), .Z(n3977) );
  AO4 U2509 ( .A(n10390), .B(n1831), .C(n1832), .D(n10554), .Z(n3978) );
  AO4 U2510 ( .A(n10389), .B(n1832), .C(n1833), .D(n10554), .Z(n3979) );
  AO4 U2511 ( .A(n10389), .B(n1833), .C(n1834), .D(n10553), .Z(n3980) );
  AO4 U2512 ( .A(n10389), .B(n1834), .C(n1835), .D(n10553), .Z(n3981) );
  AO4 U2513 ( .A(n10389), .B(n1835), .C(n1836), .D(n10553), .Z(n3982) );
  AO4 U2514 ( .A(n10389), .B(n1836), .C(n1837), .D(n10553), .Z(n3983) );
  AO4 U2515 ( .A(n10389), .B(n1837), .C(n1838), .D(n10553), .Z(n3984) );
  AO4 U2516 ( .A(n10389), .B(n1838), .C(n1839), .D(n10553), .Z(n3985) );
  AO4 U2517 ( .A(n10389), .B(n1839), .C(n1840), .D(n10553), .Z(n3986) );
  AO4 U2518 ( .A(n10389), .B(n1840), .C(n1841), .D(n10553), .Z(n3987) );
  AO4 U2519 ( .A(n10389), .B(n1841), .C(n1842), .D(n10553), .Z(n3988) );
  AO4 U2520 ( .A(n10389), .B(n1842), .C(n1843), .D(n10553), .Z(n3989) );
  AO4 U2521 ( .A(n10389), .B(n1843), .C(n10553), .D(n1394), .Z(n3990) );
  AO4 U2522 ( .A(n10553), .B(n1779), .C(n10389), .D(n1394), .Z(n5842) );
  EN U2523 ( .A(n10253), .B(n10712), .Z(n1845) );
  EN U2524 ( .A(n10246), .B(n10712), .Z(n1846) );
  EN U2525 ( .A(n10243), .B(n10712), .Z(n1847) );
  EN U2526 ( .A(n10240), .B(n10712), .Z(n1848) );
  EN U2527 ( .A(n10237), .B(n10712), .Z(n1849) );
  EN U2528 ( .A(n10234), .B(n10712), .Z(n1850) );
  EN U2529 ( .A(n10231), .B(n10712), .Z(n1851) );
  EN U2530 ( .A(n10228), .B(n10712), .Z(n1852) );
  EN U2531 ( .A(n10225), .B(n10712), .Z(n1853) );
  EN U2532 ( .A(n10222), .B(n10711), .Z(n1854) );
  EN U2533 ( .A(n10219), .B(n10711), .Z(n1855) );
  EN U2534 ( .A(n10216), .B(n10711), .Z(n1856) );
  EN U2535 ( .A(n10213), .B(n10711), .Z(n1857) );
  EN U2536 ( .A(n10210), .B(n10711), .Z(n1858) );
  EN U2537 ( .A(n10207), .B(n10711), .Z(n1859) );
  EN U2538 ( .A(n10204), .B(n10711), .Z(n1860) );
  EN U2539 ( .A(n10201), .B(n10711), .Z(n1861) );
  EN U2540 ( .A(n10198), .B(n10711), .Z(n1862) );
  EN U2541 ( .A(n10195), .B(n10711), .Z(n1863) );
  EN U2542 ( .A(n10192), .B(n10711), .Z(n1864) );
  EN U2543 ( .A(n10189), .B(n10711), .Z(n1865) );
  EN U2544 ( .A(n10186), .B(n10711), .Z(n1866) );
  EN U2545 ( .A(n10183), .B(n10711), .Z(n1867) );
  EN U2546 ( .A(n10180), .B(n10710), .Z(n1868) );
  EN U2547 ( .A(n10177), .B(n10710), .Z(n1869) );
  EN U2548 ( .A(n10174), .B(n10710), .Z(n1870) );
  EN U2549 ( .A(n10171), .B(n10710), .Z(n1871) );
  EN U2550 ( .A(n10168), .B(n10710), .Z(n1872) );
  EN U2551 ( .A(n10165), .B(n10710), .Z(n1873) );
  EN U2552 ( .A(n10162), .B(n10710), .Z(n1874) );
  EN U2553 ( .A(n10159), .B(n10710), .Z(n1875) );
  EN U2554 ( .A(n10156), .B(n10710), .Z(n1876) );
  EN U2555 ( .A(n10153), .B(n10710), .Z(n1877) );
  EN U2556 ( .A(n10150), .B(n10710), .Z(n1878) );
  EN U2557 ( .A(n10147), .B(n10710), .Z(n1879) );
  EN U2558 ( .A(n10144), .B(n10710), .Z(n1880) );
  EN U2559 ( .A(n10141), .B(n10710), .Z(n1881) );
  EN U2560 ( .A(n10138), .B(n10709), .Z(n1882) );
  EN U2561 ( .A(n10135), .B(n10709), .Z(n1883) );
  EN U2562 ( .A(n10132), .B(n10709), .Z(n1884) );
  EN U2563 ( .A(n10129), .B(n10709), .Z(n1885) );
  EN U2564 ( .A(n10126), .B(n10709), .Z(n1886) );
  EN U2565 ( .A(n10123), .B(n10709), .Z(n1887) );
  EN U2566 ( .A(n10120), .B(n10709), .Z(n1888) );
  EN U2567 ( .A(n10117), .B(n10709), .Z(n1889) );
  EN U2568 ( .A(n10114), .B(n10709), .Z(n1890) );
  EN U2569 ( .A(n10111), .B(n10709), .Z(n1891) );
  EN U2570 ( .A(n10108), .B(n10709), .Z(n1892) );
  EN U2571 ( .A(n10105), .B(n10709), .Z(n1893) );
  EN U2572 ( .A(n10102), .B(n10709), .Z(n1894) );
  EN U2573 ( .A(n10099), .B(n10709), .Z(n1895) );
  EN U2574 ( .A(n10096), .B(n10708), .Z(n1896) );
  EN U2575 ( .A(n10093), .B(n10708), .Z(n1897) );
  EN U2576 ( .A(n10090), .B(n10708), .Z(n1898) );
  EN U2577 ( .A(n10087), .B(n10708), .Z(n1899) );
  EN U2578 ( .A(n10084), .B(n10708), .Z(n1900) );
  EN U2579 ( .A(n10081), .B(n10708), .Z(n1901) );
  EN U2580 ( .A(n10078), .B(n10708), .Z(n1902) );
  EN U2581 ( .A(n10075), .B(n10708), .Z(n1903) );
  EN U2582 ( .A(n10072), .B(n10708), .Z(n1904) );
  EN U2583 ( .A(n10069), .B(n10708), .Z(n1905) );
  EN U2584 ( .A(n10066), .B(n10708), .Z(n1906) );
  EN U2585 ( .A(n10063), .B(n10708), .Z(n1907) );
  EN U2586 ( .A(n10060), .B(n10708), .Z(n1908) );
  AO4 U2587 ( .A(n10388), .B(n1845), .C(n1846), .D(n10552), .Z(n3993) );
  AO4 U2588 ( .A(n10388), .B(n1846), .C(n1847), .D(n10552), .Z(n3994) );
  AO4 U2589 ( .A(n10388), .B(n1847), .C(n1848), .D(n10552), .Z(n3995) );
  AO4 U2590 ( .A(n10388), .B(n1848), .C(n1849), .D(n10552), .Z(n3996) );
  AO4 U2591 ( .A(n10388), .B(n1849), .C(n1850), .D(n10552), .Z(n3997) );
  AO4 U2592 ( .A(n10388), .B(n1850), .C(n1851), .D(n10552), .Z(n3998) );
  AO4 U2593 ( .A(n10388), .B(n1851), .C(n1852), .D(n10552), .Z(n3999) );
  AO4 U2594 ( .A(n10388), .B(n1852), .C(n1853), .D(n10552), .Z(n4000) );
  AO4 U2595 ( .A(n10388), .B(n1853), .C(n1854), .D(n10552), .Z(n4001) );
  AO4 U2596 ( .A(n10388), .B(n1854), .C(n1855), .D(n10552), .Z(n4002) );
  AO4 U2597 ( .A(n10387), .B(n1855), .C(n1856), .D(n10552), .Z(n4003) );
  AO4 U2598 ( .A(n10387), .B(n1856), .C(n1857), .D(n10551), .Z(n4004) );
  AO4 U2599 ( .A(n10387), .B(n1857), .C(n1858), .D(n10551), .Z(n4005) );
  AO4 U2600 ( .A(n10387), .B(n1858), .C(n1859), .D(n10551), .Z(n4006) );
  AO4 U2601 ( .A(n10387), .B(n1859), .C(n1860), .D(n10551), .Z(n4007) );
  AO4 U2602 ( .A(n10387), .B(n1860), .C(n1861), .D(n10551), .Z(n4008) );
  AO4 U2603 ( .A(n10387), .B(n1861), .C(n1862), .D(n10551), .Z(n4009) );
  AO4 U2604 ( .A(n10387), .B(n1862), .C(n1863), .D(n10551), .Z(n4010) );
  AO4 U2605 ( .A(n10387), .B(n1863), .C(n1864), .D(n10551), .Z(n4011) );
  AO4 U2606 ( .A(n10387), .B(n1864), .C(n1865), .D(n10551), .Z(n4012) );
  AO4 U2607 ( .A(n10387), .B(n1865), .C(n1866), .D(n10551), .Z(n4013) );
  AO4 U2608 ( .A(n10387), .B(n1866), .C(n1867), .D(n10551), .Z(n4014) );
  AO4 U2609 ( .A(n10387), .B(n1867), .C(n1868), .D(n10551), .Z(n4015) );
  AO4 U2610 ( .A(n10387), .B(n1868), .C(n1869), .D(n10551), .Z(n4016) );
  AO4 U2611 ( .A(n10386), .B(n1869), .C(n1870), .D(n10551), .Z(n4017) );
  AO4 U2612 ( .A(n10386), .B(n1870), .C(n1871), .D(n10550), .Z(n4018) );
  AO4 U2613 ( .A(n10386), .B(n1871), .C(n1872), .D(n10550), .Z(n4019) );
  AO4 U2614 ( .A(n10386), .B(n1872), .C(n1873), .D(n10550), .Z(n4020) );
  AO4 U2615 ( .A(n10386), .B(n1873), .C(n1874), .D(n10550), .Z(n4021) );
  AO4 U2616 ( .A(n10386), .B(n1874), .C(n1875), .D(n10550), .Z(n4022) );
  AO4 U2617 ( .A(n10386), .B(n1875), .C(n1876), .D(n10550), .Z(n4023) );
  AO4 U2618 ( .A(n10386), .B(n1876), .C(n1877), .D(n10550), .Z(n4024) );
  AO4 U2619 ( .A(n10386), .B(n1877), .C(n1878), .D(n10550), .Z(n4025) );
  AO4 U2620 ( .A(n10386), .B(n1878), .C(n1879), .D(n10550), .Z(n4026) );
  AO4 U2621 ( .A(n10386), .B(n1879), .C(n1880), .D(n10550), .Z(n4027) );
  AO4 U2622 ( .A(n10386), .B(n1880), .C(n1881), .D(n10550), .Z(n4028) );
  AO4 U2623 ( .A(n10386), .B(n1881), .C(n1882), .D(n10550), .Z(n4029) );
  AO4 U2624 ( .A(n10386), .B(n1882), .C(n1883), .D(n10550), .Z(n4030) );
  AO4 U2625 ( .A(n10385), .B(n1883), .C(n1884), .D(n10550), .Z(n4031) );
  AO4 U2626 ( .A(n10385), .B(n1884), .C(n1885), .D(n10549), .Z(n4032) );
  AO4 U2627 ( .A(n10385), .B(n1885), .C(n1886), .D(n10549), .Z(n4033) );
  AO4 U2628 ( .A(n10385), .B(n1886), .C(n1887), .D(n10549), .Z(n4034) );
  AO4 U2629 ( .A(n10385), .B(n1887), .C(n1888), .D(n10549), .Z(n4035) );
  AO4 U2630 ( .A(n10385), .B(n1888), .C(n1889), .D(n10549), .Z(n4036) );
  AO4 U2631 ( .A(n10385), .B(n1889), .C(n1890), .D(n10549), .Z(n4037) );
  AO4 U2632 ( .A(n10385), .B(n1890), .C(n1891), .D(n10549), .Z(n4038) );
  AO4 U2633 ( .A(n10385), .B(n1891), .C(n1892), .D(n10549), .Z(n4039) );
  AO4 U2634 ( .A(n10385), .B(n1892), .C(n1893), .D(n10549), .Z(n4040) );
  AO4 U2635 ( .A(n10385), .B(n1893), .C(n1894), .D(n10549), .Z(n4041) );
  AO4 U2636 ( .A(n10385), .B(n1894), .C(n1895), .D(n10549), .Z(n4042) );
  AO4 U2637 ( .A(n10385), .B(n1895), .C(n1896), .D(n10549), .Z(n4043) );
  AO4 U2638 ( .A(n10385), .B(n1896), .C(n1897), .D(n10549), .Z(n4044) );
  AO4 U2639 ( .A(n10384), .B(n1897), .C(n1898), .D(n10549), .Z(n4045) );
  AO4 U2640 ( .A(n10384), .B(n1898), .C(n1899), .D(n10548), .Z(n4046) );
  AO4 U2641 ( .A(n10384), .B(n1899), .C(n1900), .D(n10548), .Z(n4047) );
  AO4 U2642 ( .A(n10384), .B(n1900), .C(n1901), .D(n10548), .Z(n4048) );
  AO4 U2643 ( .A(n10384), .B(n1901), .C(n1902), .D(n10548), .Z(n4049) );
  AO4 U2644 ( .A(n10384), .B(n1902), .C(n1903), .D(n10548), .Z(n4050) );
  AO4 U2645 ( .A(n10384), .B(n1903), .C(n1904), .D(n10548), .Z(n4051) );
  AO4 U2646 ( .A(n10384), .B(n1904), .C(n1905), .D(n10548), .Z(n4052) );
  AO4 U2647 ( .A(n10384), .B(n1905), .C(n1906), .D(n10548), .Z(n4053) );
  AO4 U2648 ( .A(n10384), .B(n1906), .C(n1907), .D(n10548), .Z(n4054) );
  AO4 U2649 ( .A(n10384), .B(n1907), .C(n1908), .D(n10548), .Z(n4055) );
  AO4 U2650 ( .A(n10384), .B(n1908), .C(n10548), .D(n1395), .Z(n4056) );
  AO4 U2651 ( .A(n10548), .B(n1844), .C(n10384), .D(n1395), .Z(n5843) );
  EN U2652 ( .A(n10253), .B(n10707), .Z(n1910) );
  EN U2653 ( .A(n10246), .B(n10707), .Z(n1911) );
  EN U2654 ( .A(n10243), .B(n10707), .Z(n1912) );
  EN U2655 ( .A(n10240), .B(n10707), .Z(n1913) );
  EN U2656 ( .A(n10237), .B(n10707), .Z(n1914) );
  EN U2657 ( .A(n10234), .B(n10707), .Z(n1915) );
  EN U2658 ( .A(n10231), .B(n10707), .Z(n1916) );
  EN U2659 ( .A(n10228), .B(n10707), .Z(n1917) );
  EN U2660 ( .A(n10225), .B(n10707), .Z(n1918) );
  EN U2661 ( .A(n10222), .B(n10706), .Z(n1919) );
  EN U2662 ( .A(n10219), .B(n10706), .Z(n1920) );
  EN U2663 ( .A(n10216), .B(n10706), .Z(n1921) );
  EN U2664 ( .A(n10213), .B(n10706), .Z(n1922) );
  EN U2665 ( .A(n10210), .B(n10706), .Z(n1923) );
  EN U2666 ( .A(n10207), .B(n10706), .Z(n1924) );
  EN U2667 ( .A(n10204), .B(n10706), .Z(n1925) );
  EN U2668 ( .A(n10201), .B(n10706), .Z(n1926) );
  EN U2669 ( .A(n10198), .B(n10706), .Z(n1927) );
  EN U2670 ( .A(n10195), .B(n10706), .Z(n1928) );
  EN U2671 ( .A(n10192), .B(n10706), .Z(n1929) );
  EN U2672 ( .A(n10189), .B(n10706), .Z(n1930) );
  EN U2673 ( .A(n10186), .B(n10706), .Z(n1931) );
  EN U2674 ( .A(n10183), .B(n10706), .Z(n1932) );
  EN U2675 ( .A(n10180), .B(n10705), .Z(n1933) );
  EN U2676 ( .A(n10177), .B(n10705), .Z(n1934) );
  EN U2677 ( .A(n10174), .B(n10705), .Z(n1935) );
  EN U2678 ( .A(n10171), .B(n10705), .Z(n1936) );
  EN U2679 ( .A(n10168), .B(n10705), .Z(n1937) );
  EN U2680 ( .A(n10165), .B(n10705), .Z(n1938) );
  EN U2681 ( .A(n10162), .B(n10705), .Z(n1939) );
  EN U2682 ( .A(n10159), .B(n10705), .Z(n1940) );
  EN U2683 ( .A(n10156), .B(n10705), .Z(n1941) );
  EN U2684 ( .A(n10153), .B(n10705), .Z(n1942) );
  EN U2685 ( .A(n10150), .B(n10705), .Z(n1943) );
  EN U2686 ( .A(n10147), .B(n10705), .Z(n1944) );
  EN U2687 ( .A(n10144), .B(n10705), .Z(n1945) );
  EN U2688 ( .A(n10141), .B(n10705), .Z(n1946) );
  EN U2689 ( .A(n10138), .B(n10704), .Z(n1947) );
  EN U2690 ( .A(n10135), .B(n10704), .Z(n1948) );
  EN U2691 ( .A(n10132), .B(n10704), .Z(n1949) );
  EN U2692 ( .A(n10129), .B(n10704), .Z(n1950) );
  EN U2693 ( .A(n10126), .B(n10704), .Z(n1951) );
  EN U2694 ( .A(n10123), .B(n10704), .Z(n1952) );
  EN U2695 ( .A(n10120), .B(n10704), .Z(n1953) );
  EN U2696 ( .A(n10117), .B(n10704), .Z(n1954) );
  EN U2697 ( .A(n10114), .B(n10704), .Z(n1955) );
  EN U2698 ( .A(n10111), .B(n10704), .Z(n1956) );
  EN U2699 ( .A(n10108), .B(n10704), .Z(n1957) );
  EN U2700 ( .A(n10105), .B(n10704), .Z(n1958) );
  EN U2701 ( .A(n10102), .B(n10704), .Z(n1959) );
  EN U2702 ( .A(n10099), .B(n10704), .Z(n1960) );
  EN U2703 ( .A(n10096), .B(n10703), .Z(n1961) );
  EN U2704 ( .A(n10093), .B(n10703), .Z(n1962) );
  EN U2705 ( .A(n10090), .B(n10703), .Z(n1963) );
  EN U2706 ( .A(n10087), .B(n10703), .Z(n1964) );
  EN U2707 ( .A(n10084), .B(n10703), .Z(n1965) );
  EN U2708 ( .A(n10081), .B(n10703), .Z(n1966) );
  EN U2709 ( .A(n10078), .B(n10703), .Z(n1967) );
  EN U2710 ( .A(n10075), .B(n10703), .Z(n1968) );
  EN U2711 ( .A(n10072), .B(n10703), .Z(n1969) );
  EN U2712 ( .A(n10069), .B(n10703), .Z(n1970) );
  EN U2713 ( .A(n10066), .B(n10703), .Z(n1971) );
  EN U2714 ( .A(n10063), .B(n10703), .Z(n1972) );
  EN U2715 ( .A(n10060), .B(n10703), .Z(n1973) );
  AO4 U2716 ( .A(n10383), .B(n1910), .C(n1911), .D(n10547), .Z(n4059) );
  AO4 U2717 ( .A(n10383), .B(n1911), .C(n1912), .D(n10547), .Z(n4060) );
  AO4 U2718 ( .A(n10383), .B(n1912), .C(n1913), .D(n10547), .Z(n4061) );
  AO4 U2719 ( .A(n10383), .B(n1913), .C(n1914), .D(n10547), .Z(n4062) );
  AO4 U2720 ( .A(n10383), .B(n1914), .C(n1915), .D(n10547), .Z(n4063) );
  AO4 U2721 ( .A(n10383), .B(n1915), .C(n1916), .D(n10547), .Z(n4064) );
  AO4 U2722 ( .A(n10383), .B(n1916), .C(n1917), .D(n10547), .Z(n4065) );
  AO4 U2723 ( .A(n10383), .B(n1917), .C(n1918), .D(n10547), .Z(n4066) );
  AO4 U2724 ( .A(n10383), .B(n1918), .C(n1919), .D(n10547), .Z(n4067) );
  AO4 U2725 ( .A(n10383), .B(n1919), .C(n1920), .D(n10547), .Z(n4068) );
  AO4 U2726 ( .A(n10382), .B(n1920), .C(n1921), .D(n10547), .Z(n4069) );
  AO4 U2727 ( .A(n10382), .B(n1921), .C(n1922), .D(n10546), .Z(n4070) );
  AO4 U2728 ( .A(n10382), .B(n1922), .C(n1923), .D(n10546), .Z(n4071) );
  AO4 U2729 ( .A(n10382), .B(n1923), .C(n1924), .D(n10546), .Z(n4072) );
  AO4 U2730 ( .A(n10382), .B(n1924), .C(n1925), .D(n10546), .Z(n4073) );
  AO4 U2731 ( .A(n10382), .B(n1925), .C(n1926), .D(n10546), .Z(n4074) );
  AO4 U2732 ( .A(n10382), .B(n1926), .C(n1927), .D(n10546), .Z(n4075) );
  AO4 U2733 ( .A(n10382), .B(n1927), .C(n1928), .D(n10546), .Z(n4076) );
  AO4 U2734 ( .A(n10382), .B(n1928), .C(n1929), .D(n10546), .Z(n4077) );
  AO4 U2735 ( .A(n10382), .B(n1929), .C(n1930), .D(n10546), .Z(n4078) );
  AO4 U2736 ( .A(n10382), .B(n1930), .C(n1931), .D(n10546), .Z(n4079) );
  AO4 U2737 ( .A(n10382), .B(n1931), .C(n1932), .D(n10546), .Z(n4080) );
  AO4 U2738 ( .A(n10382), .B(n1932), .C(n1933), .D(n10546), .Z(n4081) );
  AO4 U2739 ( .A(n10382), .B(n1933), .C(n1934), .D(n10546), .Z(n4082) );
  AO4 U2740 ( .A(n10381), .B(n1934), .C(n1935), .D(n10546), .Z(n4083) );
  AO4 U2741 ( .A(n10381), .B(n1935), .C(n1936), .D(n10545), .Z(n4084) );
  AO4 U2742 ( .A(n10381), .B(n1936), .C(n1937), .D(n10545), .Z(n4085) );
  AO4 U2743 ( .A(n10381), .B(n1937), .C(n1938), .D(n10545), .Z(n4086) );
  AO4 U2744 ( .A(n10381), .B(n1938), .C(n1939), .D(n10545), .Z(n4087) );
  AO4 U2745 ( .A(n10381), .B(n1939), .C(n1940), .D(n10545), .Z(n4088) );
  AO4 U2746 ( .A(n10381), .B(n1940), .C(n1941), .D(n10545), .Z(n4089) );
  AO4 U2747 ( .A(n10381), .B(n1941), .C(n1942), .D(n10545), .Z(n4090) );
  AO4 U2748 ( .A(n10381), .B(n1942), .C(n1943), .D(n10545), .Z(n4091) );
  AO4 U2749 ( .A(n10381), .B(n1943), .C(n1944), .D(n10545), .Z(n4092) );
  AO4 U2750 ( .A(n10381), .B(n1944), .C(n1945), .D(n10545), .Z(n4093) );
  AO4 U2751 ( .A(n10381), .B(n1945), .C(n1946), .D(n10545), .Z(n4094) );
  AO4 U2752 ( .A(n10381), .B(n1946), .C(n1947), .D(n10545), .Z(n4095) );
  AO4 U2753 ( .A(n10381), .B(n1947), .C(n1948), .D(n10545), .Z(n4096) );
  AO4 U2754 ( .A(n10380), .B(n1948), .C(n1949), .D(n10545), .Z(n4097) );
  AO4 U2755 ( .A(n10380), .B(n1949), .C(n1950), .D(n10544), .Z(n4098) );
  AO4 U2756 ( .A(n10380), .B(n1950), .C(n1951), .D(n10544), .Z(n4099) );
  AO4 U2757 ( .A(n10380), .B(n1951), .C(n1952), .D(n10544), .Z(n4100) );
  AO4 U2758 ( .A(n10380), .B(n1952), .C(n1953), .D(n10544), .Z(n4101) );
  AO4 U2759 ( .A(n10380), .B(n1953), .C(n1954), .D(n10544), .Z(n4102) );
  AO4 U2760 ( .A(n10380), .B(n1954), .C(n1955), .D(n10544), .Z(n4103) );
  AO4 U2761 ( .A(n10380), .B(n1955), .C(n1956), .D(n10544), .Z(n4104) );
  AO4 U2762 ( .A(n10380), .B(n1956), .C(n1957), .D(n10544), .Z(n4105) );
  AO4 U2763 ( .A(n10380), .B(n1957), .C(n1958), .D(n10544), .Z(n4106) );
  AO4 U2764 ( .A(n10380), .B(n1958), .C(n1959), .D(n10544), .Z(n4107) );
  AO4 U2765 ( .A(n10380), .B(n1959), .C(n1960), .D(n10544), .Z(n4108) );
  AO4 U2766 ( .A(n10380), .B(n1960), .C(n1961), .D(n10544), .Z(n4109) );
  AO4 U2767 ( .A(n10380), .B(n1961), .C(n1962), .D(n10544), .Z(n4110) );
  AO4 U2768 ( .A(n10379), .B(n1962), .C(n1963), .D(n10544), .Z(n4111) );
  AO4 U2769 ( .A(n10379), .B(n1963), .C(n1964), .D(n10543), .Z(n4112) );
  AO4 U2770 ( .A(n10379), .B(n1964), .C(n1965), .D(n10543), .Z(n4113) );
  AO4 U2771 ( .A(n10379), .B(n1965), .C(n1966), .D(n10543), .Z(n4114) );
  AO4 U2772 ( .A(n10379), .B(n1966), .C(n1967), .D(n10543), .Z(n4115) );
  AO4 U2773 ( .A(n10379), .B(n1967), .C(n1968), .D(n10543), .Z(n4116) );
  AO4 U2774 ( .A(n10379), .B(n1968), .C(n1969), .D(n10543), .Z(n4117) );
  AO4 U2775 ( .A(n10379), .B(n1969), .C(n1970), .D(n10543), .Z(n4118) );
  AO4 U2776 ( .A(n10379), .B(n1970), .C(n1971), .D(n10543), .Z(n4119) );
  AO4 U2777 ( .A(n10379), .B(n1971), .C(n1972), .D(n10543), .Z(n4120) );
  AO4 U2778 ( .A(n10379), .B(n1972), .C(n1973), .D(n10543), .Z(n4121) );
  AO4 U2779 ( .A(n10379), .B(n1973), .C(n10543), .D(n1396), .Z(n4122) );
  AO4 U2780 ( .A(n10543), .B(n1909), .C(n10379), .D(n1396), .Z(n5844) );
  EN U2781 ( .A(n10253), .B(n10702), .Z(n1975) );
  EN U2782 ( .A(n10246), .B(n10702), .Z(n1976) );
  EN U2783 ( .A(n10243), .B(n10702), .Z(n1977) );
  EN U2784 ( .A(n10240), .B(n10702), .Z(n1978) );
  EN U2785 ( .A(n10237), .B(n10702), .Z(n1979) );
  EN U2786 ( .A(n10234), .B(n10702), .Z(n1980) );
  EN U2787 ( .A(n10231), .B(n10702), .Z(n1981) );
  EN U2788 ( .A(n10228), .B(n10702), .Z(n1982) );
  EN U2789 ( .A(n10225), .B(n10702), .Z(n1983) );
  EN U2790 ( .A(n10222), .B(n10701), .Z(n1984) );
  EN U2791 ( .A(n10219), .B(n10701), .Z(n1985) );
  EN U2792 ( .A(n10216), .B(n10701), .Z(n1986) );
  EN U2793 ( .A(n10213), .B(n10701), .Z(n1987) );
  EN U2794 ( .A(n10210), .B(n10701), .Z(n1988) );
  EN U2795 ( .A(n10207), .B(n10701), .Z(n1989) );
  EN U2796 ( .A(n10204), .B(n10701), .Z(n1990) );
  EN U2797 ( .A(n10201), .B(n10701), .Z(n1991) );
  EN U2798 ( .A(n10198), .B(n10701), .Z(n1992) );
  EN U2799 ( .A(n10195), .B(n10701), .Z(n1993) );
  EN U2800 ( .A(n10192), .B(n10701), .Z(n1994) );
  EN U2801 ( .A(n10189), .B(n10701), .Z(n1995) );
  EN U2802 ( .A(n10186), .B(n10701), .Z(n1996) );
  EN U2803 ( .A(n10183), .B(n10701), .Z(n1997) );
  EN U2804 ( .A(n10180), .B(n10700), .Z(n1998) );
  EN U2805 ( .A(n10177), .B(n10700), .Z(n1999) );
  EN U2806 ( .A(n10174), .B(n10700), .Z(n2000) );
  EN U2807 ( .A(n10171), .B(n10700), .Z(n2001) );
  EN U2808 ( .A(n10168), .B(n10700), .Z(n2002) );
  EN U2809 ( .A(n10165), .B(n10700), .Z(n2003) );
  EN U2810 ( .A(n10162), .B(n10700), .Z(n2004) );
  EN U2811 ( .A(n10159), .B(n10700), .Z(n2005) );
  EN U2812 ( .A(n10156), .B(n10700), .Z(n2006) );
  EN U2813 ( .A(n10153), .B(n10700), .Z(n2007) );
  EN U2814 ( .A(n10150), .B(n10700), .Z(n2008) );
  EN U2815 ( .A(n10147), .B(n10700), .Z(n2009) );
  EN U2816 ( .A(n10144), .B(n10700), .Z(n2010) );
  EN U2817 ( .A(n10141), .B(n10700), .Z(n2011) );
  EN U2818 ( .A(n10138), .B(n10699), .Z(n2012) );
  EN U2819 ( .A(n10135), .B(n10699), .Z(n2013) );
  EN U2820 ( .A(n10132), .B(n10699), .Z(n2014) );
  EN U2821 ( .A(n10129), .B(n10699), .Z(n2015) );
  EN U2822 ( .A(n10126), .B(n10699), .Z(n2016) );
  EN U2823 ( .A(n10123), .B(n10699), .Z(n2017) );
  EN U2824 ( .A(n10120), .B(n10699), .Z(n2018) );
  EN U2825 ( .A(n10117), .B(n10699), .Z(n2019) );
  EN U2826 ( .A(n10114), .B(n10699), .Z(n2020) );
  EN U2827 ( .A(n10111), .B(n10699), .Z(n2021) );
  EN U2828 ( .A(n10108), .B(n10699), .Z(n2022) );
  EN U2829 ( .A(n10105), .B(n10699), .Z(n2023) );
  EN U2830 ( .A(n10102), .B(n10699), .Z(n2024) );
  EN U2831 ( .A(n10099), .B(n10699), .Z(n2025) );
  EN U2832 ( .A(n10096), .B(n10698), .Z(n2026) );
  EN U2833 ( .A(n10093), .B(n10698), .Z(n2027) );
  EN U2834 ( .A(n10090), .B(n10698), .Z(n2028) );
  EN U2835 ( .A(n10087), .B(n10698), .Z(n2029) );
  EN U2836 ( .A(n10084), .B(n10698), .Z(n2030) );
  EN U2837 ( .A(n10081), .B(n10698), .Z(n2031) );
  EN U2838 ( .A(n10078), .B(n10698), .Z(n2032) );
  EN U2839 ( .A(n10075), .B(n10698), .Z(n2033) );
  EN U2840 ( .A(n10072), .B(n10698), .Z(n2034) );
  EN U2841 ( .A(n10069), .B(n10698), .Z(n2035) );
  EN U2842 ( .A(n10066), .B(n10698), .Z(n2036) );
  EN U2843 ( .A(n10063), .B(n10698), .Z(n2037) );
  EN U2844 ( .A(n10060), .B(n10698), .Z(n2038) );
  AO4 U2845 ( .A(n10378), .B(n1975), .C(n1976), .D(n10542), .Z(n4125) );
  AO4 U2846 ( .A(n10378), .B(n1976), .C(n1977), .D(n10542), .Z(n4126) );
  AO4 U2847 ( .A(n10378), .B(n1977), .C(n1978), .D(n10542), .Z(n4127) );
  AO4 U2848 ( .A(n10378), .B(n1978), .C(n1979), .D(n10542), .Z(n4128) );
  AO4 U2849 ( .A(n10378), .B(n1979), .C(n1980), .D(n10542), .Z(n4129) );
  AO4 U2850 ( .A(n10378), .B(n1980), .C(n1981), .D(n10542), .Z(n4130) );
  AO4 U2851 ( .A(n10378), .B(n1981), .C(n1982), .D(n10542), .Z(n4131) );
  AO4 U2852 ( .A(n10378), .B(n1982), .C(n1983), .D(n10542), .Z(n4132) );
  AO4 U2853 ( .A(n10378), .B(n1983), .C(n1984), .D(n10542), .Z(n4133) );
  AO4 U2854 ( .A(n10378), .B(n1984), .C(n1985), .D(n10542), .Z(n4134) );
  AO4 U2855 ( .A(n10377), .B(n1985), .C(n1986), .D(n10542), .Z(n4135) );
  AO4 U2856 ( .A(n10377), .B(n1986), .C(n1987), .D(n10541), .Z(n4136) );
  AO4 U2857 ( .A(n10377), .B(n1987), .C(n1988), .D(n10541), .Z(n4137) );
  AO4 U2858 ( .A(n10377), .B(n1988), .C(n1989), .D(n10541), .Z(n4138) );
  AO4 U2859 ( .A(n10377), .B(n1989), .C(n1990), .D(n10541), .Z(n4139) );
  AO4 U2860 ( .A(n10377), .B(n1990), .C(n1991), .D(n10541), .Z(n4140) );
  AO4 U2861 ( .A(n10377), .B(n1991), .C(n1992), .D(n10541), .Z(n4141) );
  AO4 U2862 ( .A(n10377), .B(n1992), .C(n1993), .D(n10541), .Z(n4142) );
  AO4 U2863 ( .A(n10377), .B(n1993), .C(n1994), .D(n10541), .Z(n4143) );
  AO4 U2864 ( .A(n10377), .B(n1994), .C(n1995), .D(n10541), .Z(n4144) );
  AO4 U2865 ( .A(n10377), .B(n1995), .C(n1996), .D(n10541), .Z(n4145) );
  AO4 U2866 ( .A(n10377), .B(n1996), .C(n1997), .D(n10541), .Z(n4146) );
  AO4 U2867 ( .A(n10377), .B(n1997), .C(n1998), .D(n10541), .Z(n4147) );
  AO4 U2868 ( .A(n10377), .B(n1998), .C(n1999), .D(n10541), .Z(n4148) );
  AO4 U2869 ( .A(n10376), .B(n1999), .C(n2000), .D(n10541), .Z(n4149) );
  AO4 U2870 ( .A(n10376), .B(n2000), .C(n2001), .D(n10540), .Z(n4150) );
  AO4 U2871 ( .A(n10376), .B(n2001), .C(n2002), .D(n10540), .Z(n4151) );
  AO4 U2872 ( .A(n10376), .B(n2002), .C(n2003), .D(n10540), .Z(n4152) );
  AO4 U2873 ( .A(n10376), .B(n2003), .C(n2004), .D(n10540), .Z(n4153) );
  AO4 U2874 ( .A(n10376), .B(n2004), .C(n2005), .D(n10540), .Z(n4154) );
  AO4 U2875 ( .A(n10376), .B(n2005), .C(n2006), .D(n10540), .Z(n4155) );
  AO4 U2876 ( .A(n10376), .B(n2006), .C(n2007), .D(n10540), .Z(n4156) );
  AO4 U2877 ( .A(n10376), .B(n2007), .C(n2008), .D(n10540), .Z(n4157) );
  AO4 U2878 ( .A(n10376), .B(n2008), .C(n2009), .D(n10540), .Z(n4158) );
  AO4 U2879 ( .A(n10376), .B(n2009), .C(n2010), .D(n10540), .Z(n4159) );
  AO4 U2880 ( .A(n10376), .B(n2010), .C(n2011), .D(n10540), .Z(n4160) );
  AO4 U2881 ( .A(n10376), .B(n2011), .C(n2012), .D(n10540), .Z(n4161) );
  AO4 U2882 ( .A(n10376), .B(n2012), .C(n2013), .D(n10540), .Z(n4162) );
  AO4 U2883 ( .A(n10375), .B(n2013), .C(n2014), .D(n10540), .Z(n4163) );
  AO4 U2884 ( .A(n10375), .B(n2014), .C(n2015), .D(n10539), .Z(n4164) );
  AO4 U2885 ( .A(n10375), .B(n2015), .C(n2016), .D(n10539), .Z(n4165) );
  AO4 U2886 ( .A(n10375), .B(n2016), .C(n2017), .D(n10539), .Z(n4166) );
  AO4 U2887 ( .A(n10375), .B(n2017), .C(n2018), .D(n10539), .Z(n4167) );
  AO4 U2888 ( .A(n10375), .B(n2018), .C(n2019), .D(n10539), .Z(n4168) );
  AO4 U2889 ( .A(n10375), .B(n2019), .C(n2020), .D(n10539), .Z(n4169) );
  AO4 U2890 ( .A(n10375), .B(n2020), .C(n2021), .D(n10539), .Z(n4170) );
  AO4 U2891 ( .A(n10375), .B(n2021), .C(n2022), .D(n10539), .Z(n4171) );
  AO4 U2892 ( .A(n10375), .B(n2022), .C(n2023), .D(n10539), .Z(n4172) );
  AO4 U2893 ( .A(n10375), .B(n2023), .C(n2024), .D(n10539), .Z(n4173) );
  AO4 U2894 ( .A(n10375), .B(n2024), .C(n2025), .D(n10539), .Z(n4174) );
  AO4 U2895 ( .A(n10375), .B(n2025), .C(n2026), .D(n10539), .Z(n4175) );
  AO4 U2896 ( .A(n10375), .B(n2026), .C(n2027), .D(n10539), .Z(n4176) );
  AO4 U2897 ( .A(n10374), .B(n2027), .C(n2028), .D(n10539), .Z(n4177) );
  AO4 U2898 ( .A(n10374), .B(n2028), .C(n2029), .D(n10538), .Z(n4178) );
  AO4 U2899 ( .A(n10374), .B(n2029), .C(n2030), .D(n10538), .Z(n4179) );
  AO4 U2900 ( .A(n10374), .B(n2030), .C(n2031), .D(n10538), .Z(n4180) );
  AO4 U2901 ( .A(n10374), .B(n2031), .C(n2032), .D(n10538), .Z(n4181) );
  AO4 U2902 ( .A(n10374), .B(n2032), .C(n2033), .D(n10538), .Z(n4182) );
  AO4 U2903 ( .A(n10374), .B(n2033), .C(n2034), .D(n10538), .Z(n4183) );
  AO4 U2904 ( .A(n10374), .B(n2034), .C(n2035), .D(n10538), .Z(n4184) );
  AO4 U2905 ( .A(n10374), .B(n2035), .C(n2036), .D(n10538), .Z(n4185) );
  AO4 U2906 ( .A(n10374), .B(n2036), .C(n2037), .D(n10538), .Z(n4186) );
  AO4 U2907 ( .A(n10374), .B(n2037), .C(n2038), .D(n10538), .Z(n4187) );
  AO4 U2908 ( .A(n10374), .B(n2038), .C(n10538), .D(n1397), .Z(n4188) );
  AO4 U2909 ( .A(n10538), .B(n1974), .C(n10374), .D(n1397), .Z(n5845) );
  EN U2910 ( .A(n10253), .B(n10697), .Z(n2040) );
  EN U2911 ( .A(n10246), .B(n10697), .Z(n2041) );
  EN U2912 ( .A(n10243), .B(n10697), .Z(n2042) );
  EN U2913 ( .A(n10240), .B(n10697), .Z(n2043) );
  EN U2914 ( .A(n10237), .B(n10697), .Z(n2044) );
  EN U2915 ( .A(n10234), .B(n10697), .Z(n2045) );
  EN U2916 ( .A(n10231), .B(n10697), .Z(n2046) );
  EN U2917 ( .A(n10228), .B(n10697), .Z(n2047) );
  EN U2918 ( .A(n10225), .B(n10697), .Z(n2048) );
  EN U2919 ( .A(n10222), .B(n10696), .Z(n2049) );
  EN U2920 ( .A(n10219), .B(n10696), .Z(n2050) );
  EN U2921 ( .A(n10216), .B(n10696), .Z(n2051) );
  EN U2922 ( .A(n10213), .B(n10696), .Z(n2052) );
  EN U2923 ( .A(n10210), .B(n10696), .Z(n2053) );
  EN U2924 ( .A(n10207), .B(n10696), .Z(n2054) );
  EN U2925 ( .A(n10204), .B(n10696), .Z(n2055) );
  EN U2926 ( .A(n10201), .B(n10696), .Z(n2056) );
  EN U2927 ( .A(n10198), .B(n10696), .Z(n2057) );
  EN U2928 ( .A(n10195), .B(n10696), .Z(n2058) );
  EN U2929 ( .A(n10192), .B(n10696), .Z(n2059) );
  EN U2930 ( .A(n10189), .B(n10696), .Z(n2060) );
  EN U2931 ( .A(n10186), .B(n10696), .Z(n2061) );
  EN U2932 ( .A(n10183), .B(n10696), .Z(n2062) );
  EN U2933 ( .A(n10180), .B(n10695), .Z(n2063) );
  EN U2934 ( .A(n10177), .B(n10695), .Z(n2064) );
  EN U2935 ( .A(n10174), .B(n10695), .Z(n2065) );
  EN U2936 ( .A(n10171), .B(n10695), .Z(n2066) );
  EN U2937 ( .A(n10168), .B(n10695), .Z(n2067) );
  EN U2938 ( .A(n10165), .B(n10695), .Z(n2068) );
  EN U2939 ( .A(n10162), .B(n10695), .Z(n2069) );
  EN U2940 ( .A(n10159), .B(n10695), .Z(n2070) );
  EN U2941 ( .A(n10156), .B(n10695), .Z(n2071) );
  EN U2942 ( .A(n10153), .B(n10695), .Z(n2072) );
  EN U2943 ( .A(n10150), .B(n10695), .Z(n2073) );
  EN U2944 ( .A(n10147), .B(n10695), .Z(n2074) );
  EN U2945 ( .A(n10144), .B(n10695), .Z(n2075) );
  EN U2946 ( .A(n10141), .B(n10695), .Z(n2076) );
  EN U2947 ( .A(n10138), .B(n10694), .Z(n2077) );
  EN U2948 ( .A(n10135), .B(n10694), .Z(n2078) );
  EN U2949 ( .A(n10132), .B(n10694), .Z(n2079) );
  EN U2950 ( .A(n10129), .B(n10694), .Z(n2080) );
  EN U2951 ( .A(n10126), .B(n10694), .Z(n2081) );
  EN U2952 ( .A(n10123), .B(n10694), .Z(n2082) );
  EN U2953 ( .A(n10120), .B(n10694), .Z(n2083) );
  EN U2954 ( .A(n10117), .B(n10694), .Z(n2084) );
  EN U2955 ( .A(n10114), .B(n10694), .Z(n2085) );
  EN U2956 ( .A(n10111), .B(n10694), .Z(n2086) );
  EN U2957 ( .A(n10108), .B(n10694), .Z(n2087) );
  EN U2958 ( .A(n10105), .B(n10694), .Z(n2088) );
  EN U2959 ( .A(n10102), .B(n10694), .Z(n2089) );
  EN U2960 ( .A(n10099), .B(n10694), .Z(n2090) );
  EN U2961 ( .A(n10096), .B(n10693), .Z(n2091) );
  EN U2962 ( .A(n10093), .B(n10693), .Z(n2092) );
  EN U2963 ( .A(n10090), .B(n10693), .Z(n2093) );
  EN U2964 ( .A(n10087), .B(n10693), .Z(n2094) );
  EN U2965 ( .A(n10084), .B(n10693), .Z(n2095) );
  EN U2966 ( .A(n10081), .B(n10693), .Z(n2096) );
  EN U2967 ( .A(n10078), .B(n10693), .Z(n2097) );
  EN U2968 ( .A(n10075), .B(n10693), .Z(n2098) );
  EN U2969 ( .A(n10072), .B(n10693), .Z(n2099) );
  EN U2970 ( .A(n10069), .B(n10693), .Z(n2100) );
  EN U2971 ( .A(n10066), .B(n10693), .Z(n2101) );
  EN U2972 ( .A(n10063), .B(n10693), .Z(n2102) );
  EN U2973 ( .A(n10060), .B(n10693), .Z(n2103) );
  AO4 U2974 ( .A(n10373), .B(n2040), .C(n2041), .D(n10537), .Z(n4191) );
  AO4 U2975 ( .A(n10373), .B(n2041), .C(n2042), .D(n10537), .Z(n4192) );
  AO4 U2976 ( .A(n10373), .B(n2042), .C(n2043), .D(n10537), .Z(n4193) );
  AO4 U2977 ( .A(n10373), .B(n2043), .C(n2044), .D(n10537), .Z(n4194) );
  AO4 U2978 ( .A(n10373), .B(n2044), .C(n2045), .D(n10537), .Z(n4195) );
  AO4 U2979 ( .A(n10373), .B(n2045), .C(n2046), .D(n10537), .Z(n4196) );
  AO4 U2980 ( .A(n10373), .B(n2046), .C(n2047), .D(n10537), .Z(n4197) );
  AO4 U2981 ( .A(n10373), .B(n2047), .C(n2048), .D(n10537), .Z(n4198) );
  AO4 U2982 ( .A(n10373), .B(n2048), .C(n2049), .D(n10537), .Z(n4199) );
  AO4 U2983 ( .A(n10373), .B(n2049), .C(n2050), .D(n10537), .Z(n4200) );
  AO4 U2984 ( .A(n10372), .B(n2050), .C(n2051), .D(n10537), .Z(n4201) );
  AO4 U2985 ( .A(n10372), .B(n2051), .C(n2052), .D(n10536), .Z(n4202) );
  AO4 U2986 ( .A(n10372), .B(n2052), .C(n2053), .D(n10536), .Z(n4203) );
  AO4 U2987 ( .A(n10372), .B(n2053), .C(n2054), .D(n10536), .Z(n4204) );
  AO4 U2988 ( .A(n10372), .B(n2054), .C(n2055), .D(n10536), .Z(n4205) );
  AO4 U2989 ( .A(n10372), .B(n2055), .C(n2056), .D(n10536), .Z(n4206) );
  AO4 U2990 ( .A(n10372), .B(n2056), .C(n2057), .D(n10536), .Z(n4207) );
  AO4 U2991 ( .A(n10372), .B(n2057), .C(n2058), .D(n10536), .Z(n4208) );
  AO4 U2992 ( .A(n10372), .B(n2058), .C(n2059), .D(n10536), .Z(n4209) );
  AO4 U2993 ( .A(n10372), .B(n2059), .C(n2060), .D(n10536), .Z(n4210) );
  AO4 U2994 ( .A(n10372), .B(n2060), .C(n2061), .D(n10536), .Z(n4211) );
  AO4 U2995 ( .A(n10372), .B(n2061), .C(n2062), .D(n10536), .Z(n4212) );
  AO4 U2996 ( .A(n10372), .B(n2062), .C(n2063), .D(n10536), .Z(n4213) );
  AO4 U2997 ( .A(n10372), .B(n2063), .C(n2064), .D(n10536), .Z(n4214) );
  AO4 U2998 ( .A(n10371), .B(n2064), .C(n2065), .D(n10536), .Z(n4215) );
  AO4 U2999 ( .A(n10371), .B(n2065), .C(n2066), .D(n10535), .Z(n4216) );
  AO4 U3000 ( .A(n10371), .B(n2066), .C(n2067), .D(n10535), .Z(n4217) );
  AO4 U3001 ( .A(n10371), .B(n2067), .C(n2068), .D(n10535), .Z(n4218) );
  AO4 U3002 ( .A(n10371), .B(n2068), .C(n2069), .D(n10535), .Z(n4219) );
  AO4 U3003 ( .A(n10371), .B(n2069), .C(n2070), .D(n10535), .Z(n4220) );
  AO4 U3004 ( .A(n10371), .B(n2070), .C(n2071), .D(n10535), .Z(n4221) );
  AO4 U3005 ( .A(n10371), .B(n2071), .C(n2072), .D(n10535), .Z(n4222) );
  AO4 U3006 ( .A(n10371), .B(n2072), .C(n2073), .D(n10535), .Z(n4223) );
  AO4 U3007 ( .A(n10371), .B(n2073), .C(n2074), .D(n10535), .Z(n4224) );
  AO4 U3008 ( .A(n10371), .B(n2074), .C(n2075), .D(n10535), .Z(n4225) );
  AO4 U3009 ( .A(n10371), .B(n2075), .C(n2076), .D(n10535), .Z(n4226) );
  AO4 U3010 ( .A(n10371), .B(n2076), .C(n2077), .D(n10535), .Z(n4227) );
  AO4 U3011 ( .A(n10371), .B(n2077), .C(n2078), .D(n10535), .Z(n4228) );
  AO4 U3012 ( .A(n10370), .B(n2078), .C(n2079), .D(n10535), .Z(n4229) );
  AO4 U3013 ( .A(n10370), .B(n2079), .C(n2080), .D(n10534), .Z(n4230) );
  AO4 U3014 ( .A(n10370), .B(n2080), .C(n2081), .D(n10534), .Z(n4231) );
  AO4 U3015 ( .A(n10370), .B(n2081), .C(n2082), .D(n10534), .Z(n4232) );
  AO4 U3016 ( .A(n10370), .B(n2082), .C(n2083), .D(n10534), .Z(n4233) );
  AO4 U3017 ( .A(n10370), .B(n2083), .C(n2084), .D(n10534), .Z(n4234) );
  AO4 U3018 ( .A(n10370), .B(n2084), .C(n2085), .D(n10534), .Z(n4235) );
  AO4 U3019 ( .A(n10370), .B(n2085), .C(n2086), .D(n10534), .Z(n4236) );
  AO4 U3020 ( .A(n10370), .B(n2086), .C(n2087), .D(n10534), .Z(n4237) );
  AO4 U3021 ( .A(n10370), .B(n2087), .C(n2088), .D(n10534), .Z(n4238) );
  AO4 U3022 ( .A(n10370), .B(n2088), .C(n2089), .D(n10534), .Z(n4239) );
  AO4 U3023 ( .A(n10370), .B(n2089), .C(n2090), .D(n10534), .Z(n4240) );
  AO4 U3024 ( .A(n10370), .B(n2090), .C(n2091), .D(n10534), .Z(n4241) );
  AO4 U3025 ( .A(n10370), .B(n2091), .C(n2092), .D(n10534), .Z(n4242) );
  AO4 U3026 ( .A(n10369), .B(n2092), .C(n2093), .D(n10534), .Z(n4243) );
  AO4 U3027 ( .A(n10369), .B(n2093), .C(n2094), .D(n10533), .Z(n4244) );
  AO4 U3028 ( .A(n10369), .B(n2094), .C(n2095), .D(n10533), .Z(n4245) );
  AO4 U3029 ( .A(n10369), .B(n2095), .C(n2096), .D(n10533), .Z(n4246) );
  AO4 U3030 ( .A(n10369), .B(n2096), .C(n2097), .D(n10533), .Z(n4247) );
  AO4 U3031 ( .A(n10369), .B(n2097), .C(n2098), .D(n10533), .Z(n4248) );
  AO4 U3032 ( .A(n10369), .B(n2098), .C(n2099), .D(n10533), .Z(n4249) );
  AO4 U3033 ( .A(n10369), .B(n2099), .C(n2100), .D(n10533), .Z(n4250) );
  AO4 U3034 ( .A(n10369), .B(n2100), .C(n2101), .D(n10533), .Z(n4251) );
  AO4 U3035 ( .A(n10369), .B(n2101), .C(n2102), .D(n10533), .Z(n4252) );
  AO4 U3036 ( .A(n10369), .B(n2102), .C(n2103), .D(n10533), .Z(n4253) );
  AO4 U3037 ( .A(n10369), .B(n2103), .C(n10533), .D(n1398), .Z(n4254) );
  AO4 U3038 ( .A(n10533), .B(n2039), .C(n10369), .D(n1398), .Z(n5846) );
  EN U3039 ( .A(n10253), .B(n10692), .Z(n2105) );
  EN U3040 ( .A(n10246), .B(n10692), .Z(n2106) );
  EN U3041 ( .A(n10243), .B(n10692), .Z(n2107) );
  EN U3042 ( .A(n10240), .B(n10692), .Z(n2108) );
  EN U3043 ( .A(n10237), .B(n10692), .Z(n2109) );
  EN U3044 ( .A(n10234), .B(n10692), .Z(n2110) );
  EN U3045 ( .A(n10231), .B(n10692), .Z(n2111) );
  EN U3046 ( .A(n10228), .B(n10692), .Z(n2112) );
  EN U3047 ( .A(n10225), .B(n10692), .Z(n2113) );
  EN U3048 ( .A(n10222), .B(n10691), .Z(n2114) );
  EN U3049 ( .A(n10219), .B(n10691), .Z(n2115) );
  EN U3050 ( .A(n10216), .B(n10691), .Z(n2116) );
  EN U3051 ( .A(n10213), .B(n10691), .Z(n2117) );
  EN U3052 ( .A(n10210), .B(n10691), .Z(n2118) );
  EN U3053 ( .A(n10207), .B(n10691), .Z(n2119) );
  EN U3054 ( .A(n10204), .B(n10691), .Z(n2120) );
  EN U3055 ( .A(n10201), .B(n10691), .Z(n2121) );
  EN U3056 ( .A(n10198), .B(n10691), .Z(n2122) );
  EN U3057 ( .A(n10195), .B(n10691), .Z(n2123) );
  EN U3058 ( .A(n10192), .B(n10691), .Z(n2124) );
  EN U3059 ( .A(n10189), .B(n10691), .Z(n2125) );
  EN U3060 ( .A(n10186), .B(n10691), .Z(n2126) );
  EN U3061 ( .A(n10183), .B(n10691), .Z(n2127) );
  EN U3062 ( .A(n10180), .B(n10690), .Z(n2128) );
  EN U3063 ( .A(n10177), .B(n10690), .Z(n2129) );
  EN U3064 ( .A(n10174), .B(n10690), .Z(n2130) );
  EN U3065 ( .A(n10171), .B(n10690), .Z(n2131) );
  EN U3066 ( .A(n10168), .B(n10690), .Z(n2132) );
  EN U3067 ( .A(n10165), .B(n10690), .Z(n2133) );
  EN U3068 ( .A(n10162), .B(n10690), .Z(n2134) );
  EN U3069 ( .A(n10159), .B(n10690), .Z(n2135) );
  EN U3070 ( .A(n10156), .B(n10690), .Z(n2136) );
  EN U3071 ( .A(n10153), .B(n10690), .Z(n2137) );
  EN U3072 ( .A(n10150), .B(n10690), .Z(n2138) );
  EN U3073 ( .A(n10147), .B(n10690), .Z(n2139) );
  EN U3074 ( .A(n10144), .B(n10690), .Z(n2140) );
  EN U3075 ( .A(n10141), .B(n10690), .Z(n2141) );
  EN U3076 ( .A(n10138), .B(n10689), .Z(n2142) );
  EN U3077 ( .A(n10135), .B(n10689), .Z(n2143) );
  EN U3078 ( .A(n10132), .B(n10689), .Z(n2144) );
  EN U3079 ( .A(n10129), .B(n10689), .Z(n2145) );
  EN U3080 ( .A(n10126), .B(n10689), .Z(n2146) );
  EN U3081 ( .A(n10123), .B(n10689), .Z(n2147) );
  EN U3082 ( .A(n10120), .B(n10689), .Z(n2148) );
  EN U3083 ( .A(n10117), .B(n10689), .Z(n2149) );
  EN U3084 ( .A(n10114), .B(n10689), .Z(n2150) );
  EN U3085 ( .A(n10111), .B(n10689), .Z(n2151) );
  EN U3086 ( .A(n10108), .B(n10689), .Z(n2152) );
  EN U3087 ( .A(n10105), .B(n10689), .Z(n2153) );
  EN U3088 ( .A(n10102), .B(n10689), .Z(n2154) );
  EN U3089 ( .A(n10099), .B(n10689), .Z(n2155) );
  EN U3090 ( .A(n10096), .B(n10688), .Z(n2156) );
  EN U3091 ( .A(n10093), .B(n10688), .Z(n2157) );
  EN U3092 ( .A(n10090), .B(n10688), .Z(n2158) );
  EN U3093 ( .A(n10087), .B(n10688), .Z(n2159) );
  EN U3094 ( .A(n10084), .B(n10688), .Z(n2160) );
  EN U3095 ( .A(n10081), .B(n10688), .Z(n2161) );
  EN U3096 ( .A(n10078), .B(n10688), .Z(n2162) );
  EN U3097 ( .A(n10075), .B(n10688), .Z(n2163) );
  EN U3098 ( .A(n10072), .B(n10688), .Z(n2164) );
  EN U3099 ( .A(n10069), .B(n10688), .Z(n2165) );
  EN U3100 ( .A(n10066), .B(n10688), .Z(n2166) );
  EN U3101 ( .A(n10063), .B(n10688), .Z(n2167) );
  EN U3102 ( .A(n10060), .B(n10688), .Z(n2168) );
  AO4 U3103 ( .A(n10368), .B(n2105), .C(n2106), .D(n10532), .Z(n4257) );
  AO4 U3104 ( .A(n10368), .B(n2106), .C(n2107), .D(n10532), .Z(n4258) );
  AO4 U3105 ( .A(n10368), .B(n2107), .C(n2108), .D(n10532), .Z(n4259) );
  AO4 U3106 ( .A(n10368), .B(n2108), .C(n2109), .D(n10532), .Z(n4260) );
  AO4 U3107 ( .A(n10368), .B(n2109), .C(n2110), .D(n10532), .Z(n4261) );
  AO4 U3108 ( .A(n10368), .B(n2110), .C(n2111), .D(n10532), .Z(n4262) );
  AO4 U3109 ( .A(n10368), .B(n2111), .C(n2112), .D(n10532), .Z(n4263) );
  AO4 U3110 ( .A(n10368), .B(n2112), .C(n2113), .D(n10532), .Z(n4264) );
  AO4 U3111 ( .A(n10368), .B(n2113), .C(n2114), .D(n10532), .Z(n4265) );
  AO4 U3112 ( .A(n10368), .B(n2114), .C(n2115), .D(n10532), .Z(n4266) );
  AO4 U3113 ( .A(n10367), .B(n2115), .C(n2116), .D(n10532), .Z(n4267) );
  AO4 U3114 ( .A(n10367), .B(n2116), .C(n2117), .D(n10531), .Z(n4268) );
  AO4 U3115 ( .A(n10367), .B(n2117), .C(n2118), .D(n10531), .Z(n4269) );
  AO4 U3116 ( .A(n10367), .B(n2118), .C(n2119), .D(n10531), .Z(n4270) );
  AO4 U3117 ( .A(n10367), .B(n2119), .C(n2120), .D(n10531), .Z(n4271) );
  AO4 U3118 ( .A(n10367), .B(n2120), .C(n2121), .D(n10531), .Z(n4272) );
  AO4 U3119 ( .A(n10367), .B(n2121), .C(n2122), .D(n10531), .Z(n4273) );
  AO4 U3120 ( .A(n10367), .B(n2122), .C(n2123), .D(n10531), .Z(n4274) );
  AO4 U3121 ( .A(n10367), .B(n2123), .C(n2124), .D(n10531), .Z(n4275) );
  AO4 U3122 ( .A(n10367), .B(n2124), .C(n2125), .D(n10531), .Z(n4276) );
  AO4 U3123 ( .A(n10367), .B(n2125), .C(n2126), .D(n10531), .Z(n4277) );
  AO4 U3124 ( .A(n10367), .B(n2126), .C(n2127), .D(n10531), .Z(n4278) );
  AO4 U3125 ( .A(n10367), .B(n2127), .C(n2128), .D(n10531), .Z(n4279) );
  AO4 U3126 ( .A(n10367), .B(n2128), .C(n2129), .D(n10531), .Z(n4280) );
  AO4 U3127 ( .A(n10366), .B(n2129), .C(n2130), .D(n10531), .Z(n4281) );
  AO4 U3128 ( .A(n10366), .B(n2130), .C(n2131), .D(n10530), .Z(n4282) );
  AO4 U3129 ( .A(n10366), .B(n2131), .C(n2132), .D(n10530), .Z(n4283) );
  AO4 U3130 ( .A(n10366), .B(n2132), .C(n2133), .D(n10530), .Z(n4284) );
  AO4 U3131 ( .A(n10366), .B(n2133), .C(n2134), .D(n10530), .Z(n4285) );
  AO4 U3132 ( .A(n10366), .B(n2134), .C(n2135), .D(n10530), .Z(n4286) );
  AO4 U3133 ( .A(n10366), .B(n2135), .C(n2136), .D(n10530), .Z(n4287) );
  AO4 U3134 ( .A(n10366), .B(n2136), .C(n2137), .D(n10530), .Z(n4288) );
  AO4 U3135 ( .A(n10366), .B(n2137), .C(n2138), .D(n10530), .Z(n4289) );
  AO4 U3136 ( .A(n10366), .B(n2138), .C(n2139), .D(n10530), .Z(n4290) );
  AO4 U3137 ( .A(n10366), .B(n2139), .C(n2140), .D(n10530), .Z(n4291) );
  AO4 U3138 ( .A(n10366), .B(n2140), .C(n2141), .D(n10530), .Z(n4292) );
  AO4 U3139 ( .A(n10366), .B(n2141), .C(n2142), .D(n10530), .Z(n4293) );
  AO4 U3140 ( .A(n10366), .B(n2142), .C(n2143), .D(n10530), .Z(n4294) );
  AO4 U3141 ( .A(n10365), .B(n2143), .C(n2144), .D(n10530), .Z(n4295) );
  AO4 U3142 ( .A(n10365), .B(n2144), .C(n2145), .D(n10529), .Z(n4296) );
  AO4 U3143 ( .A(n10365), .B(n2145), .C(n2146), .D(n10529), .Z(n4297) );
  AO4 U3144 ( .A(n10365), .B(n2146), .C(n2147), .D(n10529), .Z(n4298) );
  AO4 U3145 ( .A(n10365), .B(n2147), .C(n2148), .D(n10529), .Z(n4299) );
  AO4 U3146 ( .A(n10365), .B(n2148), .C(n2149), .D(n10529), .Z(n4300) );
  AO4 U3147 ( .A(n10365), .B(n2149), .C(n2150), .D(n10529), .Z(n4301) );
  AO4 U3148 ( .A(n10365), .B(n2150), .C(n2151), .D(n10529), .Z(n4302) );
  AO4 U3149 ( .A(n10365), .B(n2151), .C(n2152), .D(n10529), .Z(n4303) );
  AO4 U3150 ( .A(n10365), .B(n2152), .C(n2153), .D(n10529), .Z(n4304) );
  AO4 U3151 ( .A(n10365), .B(n2153), .C(n2154), .D(n10529), .Z(n4305) );
  AO4 U3152 ( .A(n10365), .B(n2154), .C(n2155), .D(n10529), .Z(n4306) );
  AO4 U3153 ( .A(n10365), .B(n2155), .C(n2156), .D(n10529), .Z(n4307) );
  AO4 U3154 ( .A(n10365), .B(n2156), .C(n2157), .D(n10529), .Z(n4308) );
  AO4 U3155 ( .A(n10364), .B(n2157), .C(n2158), .D(n10529), .Z(n4309) );
  AO4 U3156 ( .A(n10364), .B(n2158), .C(n2159), .D(n10528), .Z(n4310) );
  AO4 U3157 ( .A(n10364), .B(n2159), .C(n2160), .D(n10528), .Z(n4311) );
  AO4 U3158 ( .A(n10364), .B(n2160), .C(n2161), .D(n10528), .Z(n4312) );
  AO4 U3159 ( .A(n10364), .B(n2161), .C(n2162), .D(n10528), .Z(n4313) );
  AO4 U3160 ( .A(n10364), .B(n2162), .C(n2163), .D(n10528), .Z(n4314) );
  AO4 U3161 ( .A(n10364), .B(n2163), .C(n2164), .D(n10528), .Z(n4315) );
  AO4 U3162 ( .A(n10364), .B(n2164), .C(n2165), .D(n10528), .Z(n4316) );
  AO4 U3163 ( .A(n10364), .B(n2165), .C(n2166), .D(n10528), .Z(n4317) );
  AO4 U3164 ( .A(n10364), .B(n2166), .C(n2167), .D(n10528), .Z(n4318) );
  AO4 U3165 ( .A(n10364), .B(n2167), .C(n2168), .D(n10528), .Z(n4319) );
  AO4 U3166 ( .A(n10364), .B(n2168), .C(n10528), .D(n1399), .Z(n4320) );
  AO4 U3167 ( .A(n10528), .B(n2104), .C(n10364), .D(n1399), .Z(n5847) );
  EN U3168 ( .A(n10253), .B(n10687), .Z(n2170) );
  EN U3169 ( .A(n10246), .B(n10687), .Z(n2171) );
  EN U3170 ( .A(n10243), .B(n10687), .Z(n2172) );
  EN U3171 ( .A(n10240), .B(n10687), .Z(n2173) );
  EN U3172 ( .A(n10237), .B(n10687), .Z(n2174) );
  EN U3173 ( .A(n10234), .B(n10687), .Z(n2175) );
  EN U3174 ( .A(n10231), .B(n10687), .Z(n2176) );
  EN U3175 ( .A(n10228), .B(n10687), .Z(n2177) );
  EN U3176 ( .A(n10225), .B(n10687), .Z(n2178) );
  EN U3177 ( .A(n10222), .B(n10686), .Z(n2179) );
  EN U3178 ( .A(n10219), .B(n10686), .Z(n2180) );
  EN U3179 ( .A(n10216), .B(n10686), .Z(n2181) );
  EN U3180 ( .A(n10213), .B(n10686), .Z(n2182) );
  EN U3181 ( .A(n10210), .B(n10686), .Z(n2183) );
  EN U3182 ( .A(n10207), .B(n10686), .Z(n2184) );
  EN U3183 ( .A(n10204), .B(n10686), .Z(n2185) );
  EN U3184 ( .A(n10201), .B(n10686), .Z(n2186) );
  EN U3185 ( .A(n10198), .B(n10686), .Z(n2187) );
  EN U3186 ( .A(n10195), .B(n10686), .Z(n2188) );
  EN U3187 ( .A(n10192), .B(n10686), .Z(n2189) );
  EN U3188 ( .A(n10189), .B(n10686), .Z(n2190) );
  EN U3189 ( .A(n10186), .B(n10686), .Z(n2191) );
  EN U3190 ( .A(n10183), .B(n10686), .Z(n2192) );
  EN U3191 ( .A(n10180), .B(n10685), .Z(n2193) );
  EN U3192 ( .A(n10177), .B(n10685), .Z(n2194) );
  EN U3193 ( .A(n10174), .B(n10685), .Z(n2195) );
  EN U3194 ( .A(n10171), .B(n10685), .Z(n2196) );
  EN U3195 ( .A(n10168), .B(n10685), .Z(n2197) );
  EN U3196 ( .A(n10165), .B(n10685), .Z(n2198) );
  EN U3197 ( .A(n10162), .B(n10685), .Z(n2199) );
  EN U3198 ( .A(n10159), .B(n10685), .Z(n2200) );
  EN U3199 ( .A(n10156), .B(n10685), .Z(n2201) );
  EN U3200 ( .A(n10153), .B(n10685), .Z(n2202) );
  EN U3201 ( .A(n10150), .B(n10685), .Z(n2203) );
  EN U3202 ( .A(n10147), .B(n10685), .Z(n2204) );
  EN U3203 ( .A(n10144), .B(n10685), .Z(n2205) );
  EN U3204 ( .A(n10141), .B(n10685), .Z(n2206) );
  EN U3205 ( .A(n10138), .B(n10684), .Z(n2207) );
  EN U3206 ( .A(n10135), .B(n10684), .Z(n2208) );
  EN U3207 ( .A(n10132), .B(n10684), .Z(n2209) );
  EN U3208 ( .A(n10129), .B(n10684), .Z(n2210) );
  EN U3209 ( .A(n10126), .B(n10684), .Z(n2211) );
  EN U3210 ( .A(n10123), .B(n10684), .Z(n2212) );
  EN U3211 ( .A(n10120), .B(n10684), .Z(n2213) );
  EN U3212 ( .A(n10117), .B(n10684), .Z(n2214) );
  EN U3213 ( .A(n10114), .B(n10684), .Z(n2215) );
  EN U3214 ( .A(n10111), .B(n10684), .Z(n2216) );
  EN U3215 ( .A(n10108), .B(n10684), .Z(n2217) );
  EN U3216 ( .A(n10105), .B(n10684), .Z(n2218) );
  EN U3217 ( .A(n10102), .B(n10684), .Z(n2219) );
  EN U3218 ( .A(n10099), .B(n10684), .Z(n2220) );
  EN U3219 ( .A(n10096), .B(n10683), .Z(n2221) );
  EN U3220 ( .A(n10093), .B(n10683), .Z(n2222) );
  EN U3221 ( .A(n10090), .B(n10683), .Z(n2223) );
  EN U3222 ( .A(n10087), .B(n10683), .Z(n2224) );
  EN U3223 ( .A(n10084), .B(n10683), .Z(n2225) );
  EN U3224 ( .A(n10081), .B(n10683), .Z(n2226) );
  EN U3225 ( .A(n10078), .B(n10683), .Z(n2227) );
  EN U3226 ( .A(n10075), .B(n10683), .Z(n2228) );
  EN U3227 ( .A(n10072), .B(n10683), .Z(n2229) );
  EN U3228 ( .A(n10069), .B(n10683), .Z(n2230) );
  EN U3229 ( .A(n10066), .B(n10683), .Z(n2231) );
  EN U3230 ( .A(n10063), .B(n10683), .Z(n2232) );
  EN U3231 ( .A(n10060), .B(n10683), .Z(n2233) );
  AO4 U3232 ( .A(n10363), .B(n2170), .C(n2171), .D(n10527), .Z(n4323) );
  AO4 U3233 ( .A(n10363), .B(n2171), .C(n2172), .D(n10527), .Z(n4324) );
  AO4 U3234 ( .A(n10363), .B(n2172), .C(n2173), .D(n10527), .Z(n4325) );
  AO4 U3235 ( .A(n10363), .B(n2173), .C(n2174), .D(n10527), .Z(n4326) );
  AO4 U3236 ( .A(n10363), .B(n2174), .C(n2175), .D(n10527), .Z(n4327) );
  AO4 U3237 ( .A(n10363), .B(n2175), .C(n2176), .D(n10527), .Z(n4328) );
  AO4 U3238 ( .A(n10363), .B(n2176), .C(n2177), .D(n10527), .Z(n4329) );
  AO4 U3239 ( .A(n10363), .B(n2177), .C(n2178), .D(n10527), .Z(n4330) );
  AO4 U3240 ( .A(n10363), .B(n2178), .C(n2179), .D(n10527), .Z(n4331) );
  AO4 U3241 ( .A(n10363), .B(n2179), .C(n2180), .D(n10527), .Z(n4332) );
  AO4 U3242 ( .A(n10362), .B(n2180), .C(n2181), .D(n10527), .Z(n4333) );
  AO4 U3243 ( .A(n10362), .B(n2181), .C(n2182), .D(n10526), .Z(n4334) );
  AO4 U3244 ( .A(n10362), .B(n2182), .C(n2183), .D(n10526), .Z(n4335) );
  AO4 U3245 ( .A(n10362), .B(n2183), .C(n2184), .D(n10526), .Z(n4336) );
  AO4 U3246 ( .A(n10362), .B(n2184), .C(n2185), .D(n10526), .Z(n4337) );
  AO4 U3247 ( .A(n10362), .B(n2185), .C(n2186), .D(n10526), .Z(n4338) );
  AO4 U3248 ( .A(n10362), .B(n2186), .C(n2187), .D(n10526), .Z(n4339) );
  AO4 U3249 ( .A(n10362), .B(n2187), .C(n2188), .D(n10526), .Z(n4340) );
  AO4 U3250 ( .A(n10362), .B(n2188), .C(n2189), .D(n10526), .Z(n4341) );
  AO4 U3251 ( .A(n10362), .B(n2189), .C(n2190), .D(n10526), .Z(n4342) );
  AO4 U3252 ( .A(n10362), .B(n2190), .C(n2191), .D(n10526), .Z(n4343) );
  AO4 U3253 ( .A(n10362), .B(n2191), .C(n2192), .D(n10526), .Z(n4344) );
  AO4 U3254 ( .A(n10362), .B(n2192), .C(n2193), .D(n10526), .Z(n4345) );
  AO4 U3255 ( .A(n10362), .B(n2193), .C(n2194), .D(n10526), .Z(n4346) );
  AO4 U3256 ( .A(n10361), .B(n2194), .C(n2195), .D(n10526), .Z(n4347) );
  AO4 U3257 ( .A(n10361), .B(n2195), .C(n2196), .D(n10525), .Z(n4348) );
  AO4 U3258 ( .A(n10361), .B(n2196), .C(n2197), .D(n10525), .Z(n4349) );
  AO4 U3259 ( .A(n10361), .B(n2197), .C(n2198), .D(n10525), .Z(n4350) );
  AO4 U3260 ( .A(n10361), .B(n2198), .C(n2199), .D(n10525), .Z(n4351) );
  AO4 U3261 ( .A(n10361), .B(n2199), .C(n2200), .D(n10525), .Z(n4352) );
  AO4 U3262 ( .A(n10361), .B(n2200), .C(n2201), .D(n10525), .Z(n4353) );
  AO4 U3263 ( .A(n10361), .B(n2201), .C(n2202), .D(n10525), .Z(n4354) );
  AO4 U3264 ( .A(n10361), .B(n2202), .C(n2203), .D(n10525), .Z(n4355) );
  AO4 U3265 ( .A(n10361), .B(n2203), .C(n2204), .D(n10525), .Z(n4356) );
  AO4 U3266 ( .A(n10361), .B(n2204), .C(n2205), .D(n10525), .Z(n4357) );
  AO4 U3267 ( .A(n10361), .B(n2205), .C(n2206), .D(n10525), .Z(n4358) );
  AO4 U3268 ( .A(n10361), .B(n2206), .C(n2207), .D(n10525), .Z(n4359) );
  AO4 U3269 ( .A(n10361), .B(n2207), .C(n2208), .D(n10525), .Z(n4360) );
  AO4 U3270 ( .A(n10360), .B(n2208), .C(n2209), .D(n10525), .Z(n4361) );
  AO4 U3271 ( .A(n10360), .B(n2209), .C(n2210), .D(n10524), .Z(n4362) );
  AO4 U3272 ( .A(n10360), .B(n2210), .C(n2211), .D(n10524), .Z(n4363) );
  AO4 U3273 ( .A(n10360), .B(n2211), .C(n2212), .D(n10524), .Z(n4364) );
  AO4 U3274 ( .A(n10360), .B(n2212), .C(n2213), .D(n10524), .Z(n4365) );
  AO4 U3275 ( .A(n10360), .B(n2213), .C(n2214), .D(n10524), .Z(n4366) );
  AO4 U3276 ( .A(n10360), .B(n2214), .C(n2215), .D(n10524), .Z(n4367) );
  AO4 U3277 ( .A(n10360), .B(n2215), .C(n2216), .D(n10524), .Z(n4368) );
  AO4 U3278 ( .A(n10360), .B(n2216), .C(n2217), .D(n10524), .Z(n4369) );
  AO4 U3279 ( .A(n10360), .B(n2217), .C(n2218), .D(n10524), .Z(n4370) );
  AO4 U3280 ( .A(n10360), .B(n2218), .C(n2219), .D(n10524), .Z(n4371) );
  AO4 U3281 ( .A(n10360), .B(n2219), .C(n2220), .D(n10524), .Z(n4372) );
  AO4 U3282 ( .A(n10360), .B(n2220), .C(n2221), .D(n10524), .Z(n4373) );
  AO4 U3283 ( .A(n10360), .B(n2221), .C(n2222), .D(n10524), .Z(n4374) );
  AO4 U3284 ( .A(n10359), .B(n2222), .C(n2223), .D(n10524), .Z(n4375) );
  AO4 U3285 ( .A(n10359), .B(n2223), .C(n2224), .D(n10523), .Z(n4376) );
  AO4 U3286 ( .A(n10359), .B(n2224), .C(n2225), .D(n10523), .Z(n4377) );
  AO4 U3287 ( .A(n10359), .B(n2225), .C(n2226), .D(n10523), .Z(n4378) );
  AO4 U3288 ( .A(n10359), .B(n2226), .C(n2227), .D(n10523), .Z(n4379) );
  AO4 U3289 ( .A(n10359), .B(n2227), .C(n2228), .D(n10523), .Z(n4380) );
  AO4 U3290 ( .A(n10359), .B(n2228), .C(n2229), .D(n10523), .Z(n4381) );
  AO4 U3291 ( .A(n10359), .B(n2229), .C(n2230), .D(n10523), .Z(n4382) );
  AO4 U3292 ( .A(n10359), .B(n2230), .C(n2231), .D(n10523), .Z(n4383) );
  AO4 U3293 ( .A(n10359), .B(n2231), .C(n2232), .D(n10523), .Z(n4384) );
  AO4 U3294 ( .A(n10359), .B(n2232), .C(n2233), .D(n10523), .Z(n4385) );
  AO4 U3295 ( .A(n10359), .B(n2233), .C(n10523), .D(n1400), .Z(n4386) );
  AO4 U3296 ( .A(n10523), .B(n2169), .C(n10359), .D(n1400), .Z(n5848) );
  EN U3297 ( .A(n10253), .B(n10682), .Z(n2235) );
  EN U3298 ( .A(n10245), .B(n10682), .Z(n2236) );
  EN U3299 ( .A(n10242), .B(n10682), .Z(n2237) );
  EN U3300 ( .A(n10239), .B(n10682), .Z(n2238) );
  EN U3301 ( .A(n10236), .B(n10682), .Z(n2239) );
  EN U3302 ( .A(n10233), .B(n10682), .Z(n2240) );
  EN U3303 ( .A(n10230), .B(n10682), .Z(n2241) );
  EN U3304 ( .A(n10227), .B(n10682), .Z(n2242) );
  EN U3305 ( .A(n10224), .B(n10682), .Z(n2243) );
  EN U3306 ( .A(n10221), .B(n10681), .Z(n2244) );
  EN U3307 ( .A(n10218), .B(n10681), .Z(n2245) );
  EN U3308 ( .A(n10215), .B(n10681), .Z(n2246) );
  EN U3309 ( .A(n10212), .B(n10681), .Z(n2247) );
  EN U3310 ( .A(n10209), .B(n10681), .Z(n2248) );
  EN U3311 ( .A(n10206), .B(n10681), .Z(n2249) );
  EN U3312 ( .A(n10203), .B(n10681), .Z(n2250) );
  EN U3313 ( .A(n10200), .B(n10681), .Z(n2251) );
  EN U3314 ( .A(n10197), .B(n10681), .Z(n2252) );
  EN U3315 ( .A(n10194), .B(n10681), .Z(n2253) );
  EN U3316 ( .A(n10191), .B(n10681), .Z(n2254) );
  EN U3317 ( .A(n10188), .B(n10681), .Z(n2255) );
  EN U3318 ( .A(n10185), .B(n10681), .Z(n2256) );
  EN U3319 ( .A(n10182), .B(n10681), .Z(n2257) );
  EN U3320 ( .A(n10179), .B(n10680), .Z(n2258) );
  EN U3321 ( .A(n10176), .B(n10680), .Z(n2259) );
  EN U3322 ( .A(n10173), .B(n10680), .Z(n2260) );
  EN U3323 ( .A(n10170), .B(n10680), .Z(n2261) );
  EN U3324 ( .A(n10167), .B(n10680), .Z(n2262) );
  EN U3325 ( .A(n10164), .B(n10680), .Z(n2263) );
  EN U3326 ( .A(n10161), .B(n10680), .Z(n2264) );
  EN U3327 ( .A(n10158), .B(n10680), .Z(n2265) );
  EN U3328 ( .A(n10155), .B(n10680), .Z(n2266) );
  EN U3329 ( .A(n10152), .B(n10680), .Z(n2267) );
  EN U3330 ( .A(n10149), .B(n10680), .Z(n2268) );
  EN U3331 ( .A(n10146), .B(n10680), .Z(n2269) );
  EN U3332 ( .A(n10143), .B(n10680), .Z(n2270) );
  EN U3333 ( .A(n10140), .B(n10680), .Z(n2271) );
  EN U3334 ( .A(n10137), .B(n10679), .Z(n2272) );
  EN U3335 ( .A(n10134), .B(n10679), .Z(n2273) );
  EN U3336 ( .A(n10131), .B(n10679), .Z(n2274) );
  EN U3337 ( .A(n10128), .B(n10679), .Z(n2275) );
  EN U3338 ( .A(n10125), .B(n10679), .Z(n2276) );
  EN U3339 ( .A(n10122), .B(n10679), .Z(n2277) );
  EN U3340 ( .A(n10119), .B(n10679), .Z(n2278) );
  EN U3341 ( .A(n10116), .B(n10679), .Z(n2279) );
  EN U3342 ( .A(n10113), .B(n10679), .Z(n2280) );
  EN U3343 ( .A(n10110), .B(n10679), .Z(n2281) );
  EN U3344 ( .A(n10107), .B(n10679), .Z(n2282) );
  EN U3345 ( .A(n10104), .B(n10679), .Z(n2283) );
  EN U3346 ( .A(n10101), .B(n10679), .Z(n2284) );
  EN U3347 ( .A(n10098), .B(n10679), .Z(n2285) );
  EN U3348 ( .A(n10095), .B(n10678), .Z(n2286) );
  EN U3349 ( .A(n10092), .B(n10678), .Z(n2287) );
  EN U3350 ( .A(n10089), .B(n10678), .Z(n2288) );
  EN U3351 ( .A(n10086), .B(n10678), .Z(n2289) );
  EN U3352 ( .A(n10083), .B(n10678), .Z(n2290) );
  EN U3353 ( .A(n10080), .B(n10678), .Z(n2291) );
  EN U3354 ( .A(n10077), .B(n10678), .Z(n2292) );
  EN U3355 ( .A(n10074), .B(n10678), .Z(n2293) );
  EN U3356 ( .A(n10071), .B(n10678), .Z(n2294) );
  EN U3357 ( .A(n10068), .B(n10678), .Z(n2295) );
  EN U3358 ( .A(n10065), .B(n10678), .Z(n2296) );
  EN U3359 ( .A(n10062), .B(n10678), .Z(n2297) );
  EN U3360 ( .A(n10059), .B(n10678), .Z(n2298) );
  AO4 U3361 ( .A(n10358), .B(n2235), .C(n2236), .D(n10522), .Z(n4389) );
  AO4 U3362 ( .A(n10358), .B(n2236), .C(n2237), .D(n10522), .Z(n4390) );
  AO4 U3363 ( .A(n10358), .B(n2237), .C(n2238), .D(n10522), .Z(n4391) );
  AO4 U3364 ( .A(n10358), .B(n2238), .C(n2239), .D(n10522), .Z(n4392) );
  AO4 U3365 ( .A(n10358), .B(n2239), .C(n2240), .D(n10522), .Z(n4393) );
  AO4 U3366 ( .A(n10358), .B(n2240), .C(n2241), .D(n10522), .Z(n4394) );
  AO4 U3367 ( .A(n10358), .B(n2241), .C(n2242), .D(n10522), .Z(n4395) );
  AO4 U3368 ( .A(n10358), .B(n2242), .C(n2243), .D(n10522), .Z(n4396) );
  AO4 U3369 ( .A(n10358), .B(n2243), .C(n2244), .D(n10522), .Z(n4397) );
  AO4 U3370 ( .A(n10358), .B(n2244), .C(n2245), .D(n10522), .Z(n4398) );
  AO4 U3371 ( .A(n10357), .B(n2245), .C(n2246), .D(n10522), .Z(n4399) );
  AO4 U3372 ( .A(n10357), .B(n2246), .C(n2247), .D(n10521), .Z(n4400) );
  AO4 U3373 ( .A(n10357), .B(n2247), .C(n2248), .D(n10521), .Z(n4401) );
  AO4 U3374 ( .A(n10357), .B(n2248), .C(n2249), .D(n10521), .Z(n4402) );
  AO4 U3375 ( .A(n10357), .B(n2249), .C(n2250), .D(n10521), .Z(n4403) );
  AO4 U3376 ( .A(n10357), .B(n2250), .C(n2251), .D(n10521), .Z(n4404) );
  AO4 U3377 ( .A(n10357), .B(n2251), .C(n2252), .D(n10521), .Z(n4405) );
  AO4 U3378 ( .A(n10357), .B(n2252), .C(n2253), .D(n10521), .Z(n4406) );
  AO4 U3379 ( .A(n10357), .B(n2253), .C(n2254), .D(n10521), .Z(n4407) );
  AO4 U3380 ( .A(n10357), .B(n2254), .C(n2255), .D(n10521), .Z(n4408) );
  AO4 U3381 ( .A(n10357), .B(n2255), .C(n2256), .D(n10521), .Z(n4409) );
  AO4 U3382 ( .A(n10357), .B(n2256), .C(n2257), .D(n10521), .Z(n4410) );
  AO4 U3383 ( .A(n10357), .B(n2257), .C(n2258), .D(n10521), .Z(n4411) );
  AO4 U3384 ( .A(n10357), .B(n2258), .C(n2259), .D(n10521), .Z(n4412) );
  AO4 U3385 ( .A(n10356), .B(n2259), .C(n2260), .D(n10521), .Z(n4413) );
  AO4 U3386 ( .A(n10356), .B(n2260), .C(n2261), .D(n10520), .Z(n4414) );
  AO4 U3387 ( .A(n10356), .B(n2261), .C(n2262), .D(n10520), .Z(n4415) );
  AO4 U3388 ( .A(n10356), .B(n2262), .C(n2263), .D(n10520), .Z(n4416) );
  AO4 U3389 ( .A(n10356), .B(n2263), .C(n2264), .D(n10520), .Z(n4417) );
  AO4 U3390 ( .A(n10356), .B(n2264), .C(n2265), .D(n10520), .Z(n4418) );
  AO4 U3391 ( .A(n10356), .B(n2265), .C(n2266), .D(n10520), .Z(n4419) );
  AO4 U3392 ( .A(n10356), .B(n2266), .C(n2267), .D(n10520), .Z(n4420) );
  AO4 U3393 ( .A(n10356), .B(n2267), .C(n2268), .D(n10520), .Z(n4421) );
  AO4 U3394 ( .A(n10356), .B(n2268), .C(n2269), .D(n10520), .Z(n4422) );
  AO4 U3395 ( .A(n10356), .B(n2269), .C(n2270), .D(n10520), .Z(n4423) );
  AO4 U3396 ( .A(n10356), .B(n2270), .C(n2271), .D(n10520), .Z(n4424) );
  AO4 U3397 ( .A(n10356), .B(n2271), .C(n2272), .D(n10520), .Z(n4425) );
  AO4 U3398 ( .A(n10356), .B(n2272), .C(n2273), .D(n10520), .Z(n4426) );
  AO4 U3399 ( .A(n10355), .B(n2273), .C(n2274), .D(n10520), .Z(n4427) );
  AO4 U3400 ( .A(n10355), .B(n2274), .C(n2275), .D(n10519), .Z(n4428) );
  AO4 U3401 ( .A(n10355), .B(n2275), .C(n2276), .D(n10519), .Z(n4429) );
  AO4 U3402 ( .A(n10355), .B(n2276), .C(n2277), .D(n10519), .Z(n4430) );
  AO4 U3403 ( .A(n10355), .B(n2277), .C(n2278), .D(n10519), .Z(n4431) );
  AO4 U3404 ( .A(n10355), .B(n2278), .C(n2279), .D(n10519), .Z(n4432) );
  AO4 U3405 ( .A(n10355), .B(n2279), .C(n2280), .D(n10519), .Z(n4433) );
  AO4 U3406 ( .A(n10355), .B(n2280), .C(n2281), .D(n10519), .Z(n4434) );
  AO4 U3407 ( .A(n10355), .B(n2281), .C(n2282), .D(n10519), .Z(n4435) );
  AO4 U3408 ( .A(n10355), .B(n2282), .C(n2283), .D(n10519), .Z(n4436) );
  AO4 U3409 ( .A(n10355), .B(n2283), .C(n2284), .D(n10519), .Z(n4437) );
  AO4 U3410 ( .A(n10355), .B(n2284), .C(n2285), .D(n10519), .Z(n4438) );
  AO4 U3411 ( .A(n10355), .B(n2285), .C(n2286), .D(n10519), .Z(n4439) );
  AO4 U3412 ( .A(n10355), .B(n2286), .C(n2287), .D(n10519), .Z(n4440) );
  AO4 U3413 ( .A(n10354), .B(n2287), .C(n2288), .D(n10519), .Z(n4441) );
  AO4 U3414 ( .A(n10354), .B(n2288), .C(n2289), .D(n10518), .Z(n4442) );
  AO4 U3415 ( .A(n10354), .B(n2289), .C(n2290), .D(n10518), .Z(n4443) );
  AO4 U3416 ( .A(n10354), .B(n2290), .C(n2291), .D(n10518), .Z(n4444) );
  AO4 U3417 ( .A(n10354), .B(n2291), .C(n2292), .D(n10518), .Z(n4445) );
  AO4 U3418 ( .A(n10354), .B(n2292), .C(n2293), .D(n10518), .Z(n4446) );
  AO4 U3419 ( .A(n10354), .B(n2293), .C(n2294), .D(n10518), .Z(n4447) );
  AO4 U3420 ( .A(n10354), .B(n2294), .C(n2295), .D(n10518), .Z(n4448) );
  AO4 U3421 ( .A(n10354), .B(n2295), .C(n2296), .D(n10518), .Z(n4449) );
  AO4 U3422 ( .A(n10354), .B(n2296), .C(n2297), .D(n10518), .Z(n4450) );
  AO4 U3423 ( .A(n10354), .B(n2297), .C(n2298), .D(n10518), .Z(n4451) );
  AO4 U3424 ( .A(n10354), .B(n2298), .C(n10518), .D(n1401), .Z(n4452) );
  AO4 U3425 ( .A(n10518), .B(n2234), .C(n10354), .D(n1401), .Z(n5849) );
  EN U3426 ( .A(n10253), .B(n10677), .Z(n2300) );
  EN U3427 ( .A(n10245), .B(n10677), .Z(n2301) );
  EN U3428 ( .A(n10242), .B(n10677), .Z(n2302) );
  EN U3429 ( .A(n10239), .B(n10677), .Z(n2303) );
  EN U3430 ( .A(n10236), .B(n10677), .Z(n2304) );
  EN U3431 ( .A(n10233), .B(n10677), .Z(n2305) );
  EN U3432 ( .A(n10230), .B(n10677), .Z(n2306) );
  EN U3433 ( .A(n10227), .B(n10677), .Z(n2307) );
  EN U3434 ( .A(n10224), .B(n10677), .Z(n2308) );
  EN U3435 ( .A(n10221), .B(n10676), .Z(n2309) );
  EN U3436 ( .A(n10218), .B(n10676), .Z(n2310) );
  EN U3437 ( .A(n10215), .B(n10676), .Z(n2311) );
  EN U3438 ( .A(n10212), .B(n10676), .Z(n2312) );
  EN U3439 ( .A(n10209), .B(n10676), .Z(n2313) );
  EN U3440 ( .A(n10206), .B(n10676), .Z(n2314) );
  EN U3441 ( .A(n10203), .B(n10676), .Z(n2315) );
  EN U3442 ( .A(n10200), .B(n10676), .Z(n2316) );
  EN U3443 ( .A(n10197), .B(n10676), .Z(n2317) );
  EN U3444 ( .A(n10194), .B(n10676), .Z(n2318) );
  EN U3445 ( .A(n10191), .B(n10676), .Z(n2319) );
  EN U3446 ( .A(n10188), .B(n10676), .Z(n2320) );
  EN U3447 ( .A(n10185), .B(n10676), .Z(n2321) );
  EN U3448 ( .A(n10182), .B(n10676), .Z(n2322) );
  EN U3449 ( .A(n10179), .B(n10675), .Z(n2323) );
  EN U3450 ( .A(n10176), .B(n10675), .Z(n2324) );
  EN U3451 ( .A(n10173), .B(n10675), .Z(n2325) );
  EN U3452 ( .A(n10170), .B(n10675), .Z(n2326) );
  EN U3453 ( .A(n10167), .B(n10675), .Z(n2327) );
  EN U3454 ( .A(n10164), .B(n10675), .Z(n2328) );
  EN U3455 ( .A(n10161), .B(n10675), .Z(n2329) );
  EN U3456 ( .A(n10158), .B(n10675), .Z(n2330) );
  EN U3457 ( .A(n10155), .B(n10675), .Z(n2331) );
  EN U3458 ( .A(n10152), .B(n10675), .Z(n2332) );
  EN U3459 ( .A(n10149), .B(n10675), .Z(n2333) );
  EN U3460 ( .A(n10146), .B(n10675), .Z(n2334) );
  EN U3461 ( .A(n10143), .B(n10675), .Z(n2335) );
  EN U3462 ( .A(n10140), .B(n10675), .Z(n2336) );
  EN U3463 ( .A(n10137), .B(n10674), .Z(n2337) );
  EN U3464 ( .A(n10134), .B(n10674), .Z(n2338) );
  EN U3465 ( .A(n10131), .B(n10674), .Z(n2339) );
  EN U3466 ( .A(n10128), .B(n10674), .Z(n2340) );
  EN U3467 ( .A(n10125), .B(n10674), .Z(n2341) );
  EN U3468 ( .A(n10122), .B(n10674), .Z(n2342) );
  EN U3469 ( .A(n10119), .B(n10674), .Z(n2343) );
  EN U3470 ( .A(n10116), .B(n10674), .Z(n2344) );
  EN U3471 ( .A(n10113), .B(n10674), .Z(n2345) );
  EN U3472 ( .A(n10110), .B(n10674), .Z(n2346) );
  EN U3473 ( .A(n10107), .B(n10674), .Z(n2347) );
  EN U3474 ( .A(n10104), .B(n10674), .Z(n2348) );
  EN U3475 ( .A(n10101), .B(n10674), .Z(n2349) );
  EN U3476 ( .A(n10098), .B(n10674), .Z(n2350) );
  EN U3477 ( .A(n10095), .B(n10673), .Z(n2351) );
  EN U3478 ( .A(n10092), .B(n10673), .Z(n2352) );
  EN U3479 ( .A(n10089), .B(n10673), .Z(n2353) );
  EN U3480 ( .A(n10086), .B(n10673), .Z(n2354) );
  EN U3481 ( .A(n10083), .B(n10673), .Z(n2355) );
  EN U3482 ( .A(n10080), .B(n10673), .Z(n2356) );
  EN U3483 ( .A(n10077), .B(n10673), .Z(n2357) );
  EN U3484 ( .A(n10074), .B(n10673), .Z(n2358) );
  EN U3485 ( .A(n10071), .B(n10673), .Z(n2359) );
  EN U3486 ( .A(n10068), .B(n10673), .Z(n2360) );
  EN U3487 ( .A(n10065), .B(n10673), .Z(n2361) );
  EN U3488 ( .A(n10062), .B(n10673), .Z(n2362) );
  EN U3489 ( .A(n10059), .B(n10673), .Z(n2363) );
  AO4 U3490 ( .A(n10353), .B(n2300), .C(n2301), .D(n10517), .Z(n4455) );
  AO4 U3491 ( .A(n10353), .B(n2301), .C(n2302), .D(n10517), .Z(n4456) );
  AO4 U3492 ( .A(n10353), .B(n2302), .C(n2303), .D(n10517), .Z(n4457) );
  AO4 U3493 ( .A(n10353), .B(n2303), .C(n2304), .D(n10517), .Z(n4458) );
  AO4 U3494 ( .A(n10353), .B(n2304), .C(n2305), .D(n10517), .Z(n4459) );
  AO4 U3495 ( .A(n10353), .B(n2305), .C(n2306), .D(n10517), .Z(n4460) );
  AO4 U3496 ( .A(n10353), .B(n2306), .C(n2307), .D(n10517), .Z(n4461) );
  AO4 U3497 ( .A(n10353), .B(n2307), .C(n2308), .D(n10517), .Z(n4462) );
  AO4 U3498 ( .A(n10353), .B(n2308), .C(n2309), .D(n10517), .Z(n4463) );
  AO4 U3499 ( .A(n10353), .B(n2309), .C(n2310), .D(n10517), .Z(n4464) );
  AO4 U3500 ( .A(n10352), .B(n2310), .C(n2311), .D(n10517), .Z(n4465) );
  AO4 U3501 ( .A(n10352), .B(n2311), .C(n2312), .D(n10516), .Z(n4466) );
  AO4 U3502 ( .A(n10352), .B(n2312), .C(n2313), .D(n10516), .Z(n4467) );
  AO4 U3503 ( .A(n10352), .B(n2313), .C(n2314), .D(n10516), .Z(n4468) );
  AO4 U3504 ( .A(n10352), .B(n2314), .C(n2315), .D(n10516), .Z(n4469) );
  AO4 U3505 ( .A(n10352), .B(n2315), .C(n2316), .D(n10516), .Z(n4470) );
  AO4 U3506 ( .A(n10352), .B(n2316), .C(n2317), .D(n10516), .Z(n4471) );
  AO4 U3507 ( .A(n10352), .B(n2317), .C(n2318), .D(n10516), .Z(n4472) );
  AO4 U3508 ( .A(n10352), .B(n2318), .C(n2319), .D(n10516), .Z(n4473) );
  AO4 U3509 ( .A(n10352), .B(n2319), .C(n2320), .D(n10516), .Z(n4474) );
  AO4 U3510 ( .A(n10352), .B(n2320), .C(n2321), .D(n10516), .Z(n4475) );
  AO4 U3511 ( .A(n10352), .B(n2321), .C(n2322), .D(n10516), .Z(n4476) );
  AO4 U3512 ( .A(n10352), .B(n2322), .C(n2323), .D(n10516), .Z(n4477) );
  AO4 U3513 ( .A(n10352), .B(n2323), .C(n2324), .D(n10516), .Z(n4478) );
  AO4 U3514 ( .A(n10351), .B(n2324), .C(n2325), .D(n10516), .Z(n4479) );
  AO4 U3515 ( .A(n10351), .B(n2325), .C(n2326), .D(n10515), .Z(n4480) );
  AO4 U3516 ( .A(n10351), .B(n2326), .C(n2327), .D(n10515), .Z(n4481) );
  AO4 U3517 ( .A(n10351), .B(n2327), .C(n2328), .D(n10515), .Z(n4482) );
  AO4 U3518 ( .A(n10351), .B(n2328), .C(n2329), .D(n10515), .Z(n4483) );
  AO4 U3519 ( .A(n10351), .B(n2329), .C(n2330), .D(n10515), .Z(n4484) );
  AO4 U3520 ( .A(n10351), .B(n2330), .C(n2331), .D(n10515), .Z(n4485) );
  AO4 U3521 ( .A(n10351), .B(n2331), .C(n2332), .D(n10515), .Z(n4486) );
  AO4 U3522 ( .A(n10351), .B(n2332), .C(n2333), .D(n10515), .Z(n4487) );
  AO4 U3523 ( .A(n10351), .B(n2333), .C(n2334), .D(n10515), .Z(n4488) );
  AO4 U3524 ( .A(n10351), .B(n2334), .C(n2335), .D(n10515), .Z(n4489) );
  AO4 U3525 ( .A(n10351), .B(n2335), .C(n2336), .D(n10515), .Z(n4490) );
  AO4 U3526 ( .A(n10351), .B(n2336), .C(n2337), .D(n10515), .Z(n4491) );
  AO4 U3527 ( .A(n10351), .B(n2337), .C(n2338), .D(n10515), .Z(n4492) );
  AO4 U3528 ( .A(n10350), .B(n2338), .C(n2339), .D(n10515), .Z(n4493) );
  AO4 U3529 ( .A(n10350), .B(n2339), .C(n2340), .D(n10514), .Z(n4494) );
  AO4 U3530 ( .A(n10350), .B(n2340), .C(n2341), .D(n10514), .Z(n4495) );
  AO4 U3531 ( .A(n10350), .B(n2341), .C(n2342), .D(n10514), .Z(n4496) );
  AO4 U3532 ( .A(n10350), .B(n2342), .C(n2343), .D(n10514), .Z(n4497) );
  AO4 U3533 ( .A(n10350), .B(n2343), .C(n2344), .D(n10514), .Z(n4498) );
  AO4 U3534 ( .A(n10350), .B(n2344), .C(n2345), .D(n10514), .Z(n4499) );
  AO4 U3535 ( .A(n10350), .B(n2345), .C(n2346), .D(n10514), .Z(n4500) );
  AO4 U3536 ( .A(n10350), .B(n2346), .C(n2347), .D(n10514), .Z(n4501) );
  AO4 U3537 ( .A(n10350), .B(n2347), .C(n2348), .D(n10514), .Z(n4502) );
  AO4 U3538 ( .A(n10350), .B(n2348), .C(n2349), .D(n10514), .Z(n4503) );
  AO4 U3539 ( .A(n10350), .B(n2349), .C(n2350), .D(n10514), .Z(n4504) );
  AO4 U3540 ( .A(n10350), .B(n2350), .C(n2351), .D(n10514), .Z(n4505) );
  AO4 U3541 ( .A(n10350), .B(n2351), .C(n2352), .D(n10514), .Z(n4506) );
  AO4 U3542 ( .A(n10349), .B(n2352), .C(n2353), .D(n10514), .Z(n4507) );
  AO4 U3543 ( .A(n10349), .B(n2353), .C(n2354), .D(n10513), .Z(n4508) );
  AO4 U3544 ( .A(n10349), .B(n2354), .C(n2355), .D(n10513), .Z(n4509) );
  AO4 U3545 ( .A(n10349), .B(n2355), .C(n2356), .D(n10513), .Z(n4510) );
  AO4 U3546 ( .A(n10349), .B(n2356), .C(n2357), .D(n10513), .Z(n4511) );
  AO4 U3547 ( .A(n10349), .B(n2357), .C(n2358), .D(n10513), .Z(n4512) );
  AO4 U3548 ( .A(n10349), .B(n2358), .C(n2359), .D(n10513), .Z(n4513) );
  AO4 U3549 ( .A(n10349), .B(n2359), .C(n2360), .D(n10513), .Z(n4514) );
  AO4 U3550 ( .A(n10349), .B(n2360), .C(n2361), .D(n10513), .Z(n4515) );
  AO4 U3551 ( .A(n10349), .B(n2361), .C(n2362), .D(n10513), .Z(n4516) );
  AO4 U3552 ( .A(n10349), .B(n2362), .C(n2363), .D(n10513), .Z(n4517) );
  AO4 U3553 ( .A(n10349), .B(n2363), .C(n10513), .D(n1402), .Z(n4518) );
  AO4 U3554 ( .A(n10513), .B(n2299), .C(n10349), .D(n1402), .Z(n5850) );
  EN U3555 ( .A(n10253), .B(n10672), .Z(n2365) );
  EN U3556 ( .A(n10245), .B(n10672), .Z(n2366) );
  EN U3557 ( .A(n10242), .B(n10672), .Z(n2367) );
  EN U3558 ( .A(n10239), .B(n10672), .Z(n2368) );
  EN U3559 ( .A(n10236), .B(n10672), .Z(n2369) );
  EN U3560 ( .A(n10233), .B(n10672), .Z(n2370) );
  EN U3561 ( .A(n10230), .B(n10672), .Z(n2371) );
  EN U3562 ( .A(n10227), .B(n10672), .Z(n2372) );
  EN U3563 ( .A(n10224), .B(n10672), .Z(n2373) );
  EN U3564 ( .A(n10221), .B(n10671), .Z(n2374) );
  EN U3565 ( .A(n10218), .B(n10671), .Z(n2375) );
  EN U3566 ( .A(n10215), .B(n10671), .Z(n2376) );
  EN U3567 ( .A(n10212), .B(n10671), .Z(n2377) );
  EN U3568 ( .A(n10209), .B(n10671), .Z(n2378) );
  EN U3569 ( .A(n10206), .B(n10671), .Z(n2379) );
  EN U3570 ( .A(n10203), .B(n10671), .Z(n2380) );
  EN U3571 ( .A(n10200), .B(n10671), .Z(n2381) );
  EN U3572 ( .A(n10197), .B(n10671), .Z(n2382) );
  EN U3573 ( .A(n10194), .B(n10671), .Z(n2383) );
  EN U3574 ( .A(n10191), .B(n10671), .Z(n2384) );
  EN U3575 ( .A(n10188), .B(n10671), .Z(n2385) );
  EN U3576 ( .A(n10185), .B(n10671), .Z(n2386) );
  EN U3577 ( .A(n10182), .B(n10671), .Z(n2387) );
  EN U3578 ( .A(n10179), .B(n10670), .Z(n2388) );
  EN U3579 ( .A(n10176), .B(n10670), .Z(n2389) );
  EN U3580 ( .A(n10173), .B(n10670), .Z(n2390) );
  EN U3581 ( .A(n10170), .B(n10670), .Z(n2391) );
  EN U3582 ( .A(n10167), .B(n10670), .Z(n2392) );
  EN U3583 ( .A(n10164), .B(n10670), .Z(n2393) );
  EN U3584 ( .A(n10161), .B(n10670), .Z(n2394) );
  EN U3585 ( .A(n10158), .B(n10670), .Z(n2395) );
  EN U3586 ( .A(n10155), .B(n10670), .Z(n2396) );
  EN U3587 ( .A(n10152), .B(n10670), .Z(n2397) );
  EN U3588 ( .A(n10149), .B(n10670), .Z(n2398) );
  EN U3589 ( .A(n10146), .B(n10670), .Z(n2399) );
  EN U3590 ( .A(n10143), .B(n10670), .Z(n2400) );
  EN U3591 ( .A(n10140), .B(n10670), .Z(n2401) );
  EN U3592 ( .A(n10137), .B(n10669), .Z(n2402) );
  EN U3593 ( .A(n10134), .B(n10669), .Z(n2403) );
  EN U3594 ( .A(n10131), .B(n10669), .Z(n2404) );
  EN U3595 ( .A(n10128), .B(n10669), .Z(n2405) );
  EN U3596 ( .A(n10125), .B(n10669), .Z(n2406) );
  EN U3597 ( .A(n10122), .B(n10669), .Z(n2407) );
  EN U3598 ( .A(n10119), .B(n10669), .Z(n2408) );
  EN U3599 ( .A(n10116), .B(n10669), .Z(n2409) );
  EN U3600 ( .A(n10113), .B(n10669), .Z(n2410) );
  EN U3601 ( .A(n10110), .B(n10669), .Z(n2411) );
  EN U3602 ( .A(n10107), .B(n10669), .Z(n2412) );
  EN U3603 ( .A(n10104), .B(n10669), .Z(n2413) );
  EN U3604 ( .A(n10101), .B(n10669), .Z(n2414) );
  EN U3605 ( .A(n10098), .B(n10669), .Z(n2415) );
  EN U3606 ( .A(n10095), .B(n10668), .Z(n2416) );
  EN U3607 ( .A(n10092), .B(n10668), .Z(n2417) );
  EN U3608 ( .A(n10089), .B(n10668), .Z(n2418) );
  EN U3609 ( .A(n10086), .B(n10668), .Z(n2419) );
  EN U3610 ( .A(n10083), .B(n10668), .Z(n2420) );
  EN U3611 ( .A(n10080), .B(n10668), .Z(n2421) );
  EN U3612 ( .A(n10077), .B(n10668), .Z(n2422) );
  EN U3613 ( .A(n10074), .B(n10668), .Z(n2423) );
  EN U3614 ( .A(n10071), .B(n10668), .Z(n2424) );
  EN U3615 ( .A(n10068), .B(n10668), .Z(n2425) );
  EN U3616 ( .A(n10065), .B(n10668), .Z(n2426) );
  EN U3617 ( .A(n10062), .B(n10668), .Z(n2427) );
  EN U3618 ( .A(n10059), .B(n10668), .Z(n2428) );
  AO4 U3619 ( .A(n10348), .B(n2365), .C(n2366), .D(n10512), .Z(n4521) );
  AO4 U3620 ( .A(n10348), .B(n2366), .C(n2367), .D(n10512), .Z(n4522) );
  AO4 U3621 ( .A(n10348), .B(n2367), .C(n2368), .D(n10512), .Z(n4523) );
  AO4 U3622 ( .A(n10348), .B(n2368), .C(n2369), .D(n10512), .Z(n4524) );
  AO4 U3623 ( .A(n10348), .B(n2369), .C(n2370), .D(n10512), .Z(n4525) );
  AO4 U3624 ( .A(n10348), .B(n2370), .C(n2371), .D(n10512), .Z(n4526) );
  AO4 U3625 ( .A(n10348), .B(n2371), .C(n2372), .D(n10512), .Z(n4527) );
  AO4 U3626 ( .A(n10348), .B(n2372), .C(n2373), .D(n10512), .Z(n4528) );
  AO4 U3627 ( .A(n10348), .B(n2373), .C(n2374), .D(n10512), .Z(n4529) );
  AO4 U3628 ( .A(n10348), .B(n2374), .C(n2375), .D(n10512), .Z(n4530) );
  AO4 U3629 ( .A(n10347), .B(n2375), .C(n2376), .D(n10512), .Z(n4531) );
  AO4 U3630 ( .A(n10347), .B(n2376), .C(n2377), .D(n10511), .Z(n4532) );
  AO4 U3631 ( .A(n10347), .B(n2377), .C(n2378), .D(n10511), .Z(n4533) );
  AO4 U3632 ( .A(n10347), .B(n2378), .C(n2379), .D(n10511), .Z(n4534) );
  AO4 U3633 ( .A(n10347), .B(n2379), .C(n2380), .D(n10511), .Z(n4535) );
  AO4 U3634 ( .A(n10347), .B(n2380), .C(n2381), .D(n10511), .Z(n4536) );
  AO4 U3635 ( .A(n10347), .B(n2381), .C(n2382), .D(n10511), .Z(n4537) );
  AO4 U3636 ( .A(n10347), .B(n2382), .C(n2383), .D(n10511), .Z(n4538) );
  AO4 U3637 ( .A(n10347), .B(n2383), .C(n2384), .D(n10511), .Z(n4539) );
  AO4 U3638 ( .A(n10347), .B(n2384), .C(n2385), .D(n10511), .Z(n4540) );
  AO4 U3639 ( .A(n10347), .B(n2385), .C(n2386), .D(n10511), .Z(n4541) );
  AO4 U3640 ( .A(n10347), .B(n2386), .C(n2387), .D(n10511), .Z(n4542) );
  AO4 U3641 ( .A(n10347), .B(n2387), .C(n2388), .D(n10511), .Z(n4543) );
  AO4 U3642 ( .A(n10347), .B(n2388), .C(n2389), .D(n10511), .Z(n4544) );
  AO4 U3643 ( .A(n10346), .B(n2389), .C(n2390), .D(n10511), .Z(n4545) );
  AO4 U3644 ( .A(n10346), .B(n2390), .C(n2391), .D(n10510), .Z(n4546) );
  AO4 U3645 ( .A(n10346), .B(n2391), .C(n2392), .D(n10510), .Z(n4547) );
  AO4 U3646 ( .A(n10346), .B(n2392), .C(n2393), .D(n10510), .Z(n4548) );
  AO4 U3647 ( .A(n10346), .B(n2393), .C(n2394), .D(n10510), .Z(n4549) );
  AO4 U3648 ( .A(n10346), .B(n2394), .C(n2395), .D(n10510), .Z(n4550) );
  AO4 U3649 ( .A(n10346), .B(n2395), .C(n2396), .D(n10510), .Z(n4551) );
  AO4 U3650 ( .A(n10346), .B(n2396), .C(n2397), .D(n10510), .Z(n4552) );
  AO4 U3651 ( .A(n10346), .B(n2397), .C(n2398), .D(n10510), .Z(n4553) );
  AO4 U3652 ( .A(n10346), .B(n2398), .C(n2399), .D(n10510), .Z(n4554) );
  AO4 U3653 ( .A(n10346), .B(n2399), .C(n2400), .D(n10510), .Z(n4555) );
  AO4 U3654 ( .A(n10346), .B(n2400), .C(n2401), .D(n10510), .Z(n4556) );
  AO4 U3655 ( .A(n10346), .B(n2401), .C(n2402), .D(n10510), .Z(n4557) );
  AO4 U3656 ( .A(n10346), .B(n2402), .C(n2403), .D(n10510), .Z(n4558) );
  AO4 U3657 ( .A(n10345), .B(n2403), .C(n2404), .D(n10510), .Z(n4559) );
  AO4 U3658 ( .A(n10345), .B(n2404), .C(n2405), .D(n10509), .Z(n4560) );
  AO4 U3659 ( .A(n10345), .B(n2405), .C(n2406), .D(n10509), .Z(n4561) );
  AO4 U3660 ( .A(n10345), .B(n2406), .C(n2407), .D(n10509), .Z(n4562) );
  AO4 U3661 ( .A(n10345), .B(n2407), .C(n2408), .D(n10509), .Z(n4563) );
  AO4 U3662 ( .A(n10345), .B(n2408), .C(n2409), .D(n10509), .Z(n4564) );
  AO4 U3663 ( .A(n10345), .B(n2409), .C(n2410), .D(n10509), .Z(n4565) );
  AO4 U3664 ( .A(n10345), .B(n2410), .C(n2411), .D(n10509), .Z(n4566) );
  AO4 U3665 ( .A(n10345), .B(n2411), .C(n2412), .D(n10509), .Z(n4567) );
  AO4 U3666 ( .A(n10345), .B(n2412), .C(n2413), .D(n10509), .Z(n4568) );
  AO4 U3667 ( .A(n10345), .B(n2413), .C(n2414), .D(n10509), .Z(n4569) );
  AO4 U3668 ( .A(n10345), .B(n2414), .C(n2415), .D(n10509), .Z(n4570) );
  AO4 U3669 ( .A(n10345), .B(n2415), .C(n2416), .D(n10509), .Z(n4571) );
  AO4 U3670 ( .A(n10345), .B(n2416), .C(n2417), .D(n10509), .Z(n4572) );
  AO4 U3671 ( .A(n10344), .B(n2417), .C(n2418), .D(n10509), .Z(n4573) );
  AO4 U3672 ( .A(n10344), .B(n2418), .C(n2419), .D(n10508), .Z(n4574) );
  AO4 U3673 ( .A(n10344), .B(n2419), .C(n2420), .D(n10508), .Z(n4575) );
  AO4 U3674 ( .A(n10344), .B(n2420), .C(n2421), .D(n10508), .Z(n4576) );
  AO4 U3675 ( .A(n10344), .B(n2421), .C(n2422), .D(n10508), .Z(n4577) );
  AO4 U3676 ( .A(n10344), .B(n2422), .C(n2423), .D(n10508), .Z(n4578) );
  AO4 U3677 ( .A(n10344), .B(n2423), .C(n2424), .D(n10508), .Z(n4579) );
  AO4 U3678 ( .A(n10344), .B(n2424), .C(n2425), .D(n10508), .Z(n4580) );
  AO4 U3679 ( .A(n10344), .B(n2425), .C(n2426), .D(n10508), .Z(n4581) );
  AO4 U3680 ( .A(n10344), .B(n2426), .C(n2427), .D(n10508), .Z(n4582) );
  AO4 U3681 ( .A(n10344), .B(n2427), .C(n2428), .D(n10508), .Z(n4583) );
  AO4 U3682 ( .A(n10344), .B(n2428), .C(n10508), .D(n1403), .Z(n4584) );
  AO4 U3683 ( .A(n10508), .B(n2364), .C(n10344), .D(n1403), .Z(n5851) );
  EN U3684 ( .A(n10252), .B(n10667), .Z(n2430) );
  EN U3685 ( .A(n10245), .B(n10667), .Z(n2431) );
  EN U3686 ( .A(n10242), .B(n10667), .Z(n2432) );
  EN U3687 ( .A(n10239), .B(n10667), .Z(n2433) );
  EN U3688 ( .A(n10236), .B(n10667), .Z(n2434) );
  EN U3689 ( .A(n10233), .B(n10667), .Z(n2435) );
  EN U3690 ( .A(n10230), .B(n10667), .Z(n2436) );
  EN U3691 ( .A(n10227), .B(n10667), .Z(n2437) );
  EN U3692 ( .A(n10224), .B(n10667), .Z(n2438) );
  EN U3693 ( .A(n10221), .B(n10666), .Z(n2439) );
  EN U3694 ( .A(n10218), .B(n10666), .Z(n2440) );
  EN U3695 ( .A(n10215), .B(n10666), .Z(n2441) );
  EN U3696 ( .A(n10212), .B(n10666), .Z(n2442) );
  EN U3697 ( .A(n10209), .B(n10666), .Z(n2443) );
  EN U3698 ( .A(n10206), .B(n10666), .Z(n2444) );
  EN U3699 ( .A(n10203), .B(n10666), .Z(n2445) );
  EN U3700 ( .A(n10200), .B(n10666), .Z(n2446) );
  EN U3701 ( .A(n10197), .B(n10666), .Z(n2447) );
  EN U3702 ( .A(n10194), .B(n10666), .Z(n2448) );
  EN U3703 ( .A(n10191), .B(n10666), .Z(n2449) );
  EN U3704 ( .A(n10188), .B(n10666), .Z(n2450) );
  EN U3705 ( .A(n10185), .B(n10666), .Z(n2451) );
  EN U3706 ( .A(n10182), .B(n10666), .Z(n2452) );
  EN U3707 ( .A(n10179), .B(n10665), .Z(n2453) );
  EN U3708 ( .A(n10176), .B(n10665), .Z(n2454) );
  EN U3709 ( .A(n10173), .B(n10665), .Z(n2455) );
  EN U3710 ( .A(n10170), .B(n10665), .Z(n2456) );
  EN U3711 ( .A(n10167), .B(n10665), .Z(n2457) );
  EN U3712 ( .A(n10164), .B(n10665), .Z(n2458) );
  EN U3713 ( .A(n10161), .B(n10665), .Z(n2459) );
  EN U3714 ( .A(n10158), .B(n10665), .Z(n2460) );
  EN U3715 ( .A(n10155), .B(n10665), .Z(n2461) );
  EN U3716 ( .A(n10152), .B(n10665), .Z(n2462) );
  EN U3717 ( .A(n10149), .B(n10665), .Z(n2463) );
  EN U3718 ( .A(n10146), .B(n10665), .Z(n2464) );
  EN U3719 ( .A(n10143), .B(n10665), .Z(n2465) );
  EN U3720 ( .A(n10140), .B(n10665), .Z(n2466) );
  EN U3721 ( .A(n10137), .B(n10664), .Z(n2467) );
  EN U3722 ( .A(n10134), .B(n10664), .Z(n2468) );
  EN U3723 ( .A(n10131), .B(n10664), .Z(n2469) );
  EN U3724 ( .A(n10128), .B(n10664), .Z(n2470) );
  EN U3725 ( .A(n10125), .B(n10664), .Z(n2471) );
  EN U3726 ( .A(n10122), .B(n10664), .Z(n2472) );
  EN U3727 ( .A(n10119), .B(n10664), .Z(n2473) );
  EN U3728 ( .A(n10116), .B(n10664), .Z(n2474) );
  EN U3729 ( .A(n10113), .B(n10664), .Z(n2475) );
  EN U3730 ( .A(n10110), .B(n10664), .Z(n2476) );
  EN U3731 ( .A(n10107), .B(n10664), .Z(n2477) );
  EN U3732 ( .A(n10104), .B(n10664), .Z(n2478) );
  EN U3733 ( .A(n10101), .B(n10664), .Z(n2479) );
  EN U3734 ( .A(n10098), .B(n10664), .Z(n2480) );
  EN U3735 ( .A(n10095), .B(n10663), .Z(n2481) );
  EN U3736 ( .A(n10092), .B(n10663), .Z(n2482) );
  EN U3737 ( .A(n10089), .B(n10663), .Z(n2483) );
  EN U3738 ( .A(n10086), .B(n10663), .Z(n2484) );
  EN U3739 ( .A(n10083), .B(n10663), .Z(n2485) );
  EN U3740 ( .A(n10080), .B(n10663), .Z(n2486) );
  EN U3741 ( .A(n10077), .B(n10663), .Z(n2487) );
  EN U3742 ( .A(n10074), .B(n10663), .Z(n2488) );
  EN U3743 ( .A(n10071), .B(n10663), .Z(n2489) );
  EN U3744 ( .A(n10068), .B(n10663), .Z(n2490) );
  EN U3745 ( .A(n10065), .B(n10663), .Z(n2491) );
  EN U3746 ( .A(n10062), .B(n10663), .Z(n2492) );
  EN U3747 ( .A(n10059), .B(n10663), .Z(n2493) );
  AO4 U3748 ( .A(n10343), .B(n2430), .C(n2431), .D(n10507), .Z(n4587) );
  AO4 U3749 ( .A(n10343), .B(n2431), .C(n2432), .D(n10507), .Z(n4588) );
  AO4 U3750 ( .A(n10343), .B(n2432), .C(n2433), .D(n10507), .Z(n4589) );
  AO4 U3751 ( .A(n10343), .B(n2433), .C(n2434), .D(n10507), .Z(n4590) );
  AO4 U3752 ( .A(n10343), .B(n2434), .C(n2435), .D(n10507), .Z(n4591) );
  AO4 U3753 ( .A(n10343), .B(n2435), .C(n2436), .D(n10507), .Z(n4592) );
  AO4 U3754 ( .A(n10343), .B(n2436), .C(n2437), .D(n10507), .Z(n4593) );
  AO4 U3755 ( .A(n10343), .B(n2437), .C(n2438), .D(n10507), .Z(n4594) );
  AO4 U3756 ( .A(n10343), .B(n2438), .C(n2439), .D(n10507), .Z(n4595) );
  AO4 U3757 ( .A(n10343), .B(n2439), .C(n2440), .D(n10507), .Z(n4596) );
  AO4 U3758 ( .A(n10342), .B(n2440), .C(n2441), .D(n10507), .Z(n4597) );
  AO4 U3759 ( .A(n10342), .B(n2441), .C(n2442), .D(n10506), .Z(n4598) );
  AO4 U3760 ( .A(n10342), .B(n2442), .C(n2443), .D(n10506), .Z(n4599) );
  AO4 U3761 ( .A(n10342), .B(n2443), .C(n2444), .D(n10506), .Z(n4600) );
  AO4 U3762 ( .A(n10342), .B(n2444), .C(n2445), .D(n10506), .Z(n4601) );
  AO4 U3763 ( .A(n10342), .B(n2445), .C(n2446), .D(n10506), .Z(n4602) );
  AO4 U3764 ( .A(n10342), .B(n2446), .C(n2447), .D(n10506), .Z(n4603) );
  AO4 U3765 ( .A(n10342), .B(n2447), .C(n2448), .D(n10506), .Z(n4604) );
  AO4 U3766 ( .A(n10342), .B(n2448), .C(n2449), .D(n10506), .Z(n4605) );
  AO4 U3767 ( .A(n10342), .B(n2449), .C(n2450), .D(n10506), .Z(n4606) );
  AO4 U3768 ( .A(n10342), .B(n2450), .C(n2451), .D(n10506), .Z(n4607) );
  AO4 U3769 ( .A(n10342), .B(n2451), .C(n2452), .D(n10506), .Z(n4608) );
  AO4 U3770 ( .A(n10342), .B(n2452), .C(n2453), .D(n10506), .Z(n4609) );
  AO4 U3771 ( .A(n10342), .B(n2453), .C(n2454), .D(n10506), .Z(n4610) );
  AO4 U3772 ( .A(n10341), .B(n2454), .C(n2455), .D(n10506), .Z(n4611) );
  AO4 U3773 ( .A(n10341), .B(n2455), .C(n2456), .D(n10505), .Z(n4612) );
  AO4 U3774 ( .A(n10341), .B(n2456), .C(n2457), .D(n10505), .Z(n4613) );
  AO4 U3775 ( .A(n10341), .B(n2457), .C(n2458), .D(n10505), .Z(n4614) );
  AO4 U3776 ( .A(n10341), .B(n2458), .C(n2459), .D(n10505), .Z(n4615) );
  AO4 U3777 ( .A(n10341), .B(n2459), .C(n2460), .D(n10505), .Z(n4616) );
  AO4 U3778 ( .A(n10341), .B(n2460), .C(n2461), .D(n10505), .Z(n4617) );
  AO4 U3779 ( .A(n10341), .B(n2461), .C(n2462), .D(n10505), .Z(n4618) );
  AO4 U3780 ( .A(n10341), .B(n2462), .C(n2463), .D(n10505), .Z(n4619) );
  AO4 U3781 ( .A(n10341), .B(n2463), .C(n2464), .D(n10505), .Z(n4620) );
  AO4 U3782 ( .A(n10341), .B(n2464), .C(n2465), .D(n10505), .Z(n4621) );
  AO4 U3783 ( .A(n10341), .B(n2465), .C(n2466), .D(n10505), .Z(n4622) );
  AO4 U3784 ( .A(n10341), .B(n2466), .C(n2467), .D(n10505), .Z(n4623) );
  AO4 U3785 ( .A(n10341), .B(n2467), .C(n2468), .D(n10505), .Z(n4624) );
  AO4 U3786 ( .A(n10340), .B(n2468), .C(n2469), .D(n10505), .Z(n4625) );
  AO4 U3787 ( .A(n10340), .B(n2469), .C(n2470), .D(n10504), .Z(n4626) );
  AO4 U3788 ( .A(n10340), .B(n2470), .C(n2471), .D(n10504), .Z(n4627) );
  AO4 U3789 ( .A(n10340), .B(n2471), .C(n2472), .D(n10504), .Z(n4628) );
  AO4 U3790 ( .A(n10340), .B(n2472), .C(n2473), .D(n10504), .Z(n4629) );
  AO4 U3791 ( .A(n10340), .B(n2473), .C(n2474), .D(n10504), .Z(n4630) );
  AO4 U3792 ( .A(n10340), .B(n2474), .C(n2475), .D(n10504), .Z(n4631) );
  AO4 U3793 ( .A(n10340), .B(n2475), .C(n2476), .D(n10504), .Z(n4632) );
  AO4 U3794 ( .A(n10340), .B(n2476), .C(n2477), .D(n10504), .Z(n4633) );
  AO4 U3795 ( .A(n10340), .B(n2477), .C(n2478), .D(n10504), .Z(n4634) );
  AO4 U3796 ( .A(n10340), .B(n2478), .C(n2479), .D(n10504), .Z(n4635) );
  AO4 U3797 ( .A(n10340), .B(n2479), .C(n2480), .D(n10504), .Z(n4636) );
  AO4 U3798 ( .A(n10340), .B(n2480), .C(n2481), .D(n10504), .Z(n4637) );
  AO4 U3799 ( .A(n10340), .B(n2481), .C(n2482), .D(n10504), .Z(n4638) );
  AO4 U3800 ( .A(n10339), .B(n2482), .C(n2483), .D(n10504), .Z(n4639) );
  AO4 U3801 ( .A(n10339), .B(n2483), .C(n2484), .D(n10503), .Z(n4640) );
  AO4 U3802 ( .A(n10339), .B(n2484), .C(n2485), .D(n10503), .Z(n4641) );
  AO4 U3803 ( .A(n10339), .B(n2485), .C(n2486), .D(n10503), .Z(n4642) );
  AO4 U3804 ( .A(n10339), .B(n2486), .C(n2487), .D(n10503), .Z(n4643) );
  AO4 U3805 ( .A(n10339), .B(n2487), .C(n2488), .D(n10503), .Z(n4644) );
  AO4 U3806 ( .A(n10339), .B(n2488), .C(n2489), .D(n10503), .Z(n4645) );
  AO4 U3807 ( .A(n10339), .B(n2489), .C(n2490), .D(n10503), .Z(n4646) );
  AO4 U3808 ( .A(n10339), .B(n2490), .C(n2491), .D(n10503), .Z(n4647) );
  AO4 U3809 ( .A(n10339), .B(n2491), .C(n2492), .D(n10503), .Z(n4648) );
  AO4 U3810 ( .A(n10339), .B(n2492), .C(n2493), .D(n10503), .Z(n4649) );
  AO4 U3811 ( .A(n10339), .B(n2493), .C(n10503), .D(n1404), .Z(n4650) );
  AO4 U3812 ( .A(n10503), .B(n2429), .C(n10339), .D(n1404), .Z(n5852) );
  EN U3813 ( .A(n10252), .B(n10662), .Z(n2495) );
  EN U3814 ( .A(n10245), .B(n10662), .Z(n2496) );
  EN U3815 ( .A(n10242), .B(n10662), .Z(n2497) );
  EN U3816 ( .A(n10239), .B(n10662), .Z(n2498) );
  EN U3817 ( .A(n10236), .B(n10662), .Z(n2499) );
  EN U3818 ( .A(n10233), .B(n10662), .Z(n2500) );
  EN U3819 ( .A(n10230), .B(n10662), .Z(n2501) );
  EN U3820 ( .A(n10227), .B(n10662), .Z(n2502) );
  EN U3821 ( .A(n10224), .B(n10662), .Z(n2503) );
  EN U3822 ( .A(n10221), .B(n10661), .Z(n2504) );
  EN U3823 ( .A(n10218), .B(n10661), .Z(n2505) );
  EN U3824 ( .A(n10215), .B(n10661), .Z(n2506) );
  EN U3825 ( .A(n10212), .B(n10661), .Z(n2507) );
  EN U3826 ( .A(n10209), .B(n10661), .Z(n2508) );
  EN U3827 ( .A(n10206), .B(n10661), .Z(n2509) );
  EN U3828 ( .A(n10203), .B(n10661), .Z(n2510) );
  EN U3829 ( .A(n10200), .B(n10661), .Z(n2511) );
  EN U3830 ( .A(n10197), .B(n10661), .Z(n2512) );
  EN U3831 ( .A(n10194), .B(n10661), .Z(n2513) );
  EN U3832 ( .A(n10191), .B(n10661), .Z(n2514) );
  EN U3833 ( .A(n10188), .B(n10661), .Z(n2515) );
  EN U3834 ( .A(n10185), .B(n10661), .Z(n2516) );
  EN U3835 ( .A(n10182), .B(n10661), .Z(n2517) );
  EN U3836 ( .A(n10179), .B(n10660), .Z(n2518) );
  EN U3837 ( .A(n10176), .B(n10660), .Z(n2519) );
  EN U3838 ( .A(n10173), .B(n10660), .Z(n2520) );
  EN U3839 ( .A(n10170), .B(n10660), .Z(n2521) );
  EN U3840 ( .A(n10167), .B(n10660), .Z(n2522) );
  EN U3841 ( .A(n10164), .B(n10660), .Z(n2523) );
  EN U3842 ( .A(n10161), .B(n10660), .Z(n2524) );
  EN U3843 ( .A(n10158), .B(n10660), .Z(n2525) );
  EN U3844 ( .A(n10155), .B(n10660), .Z(n2526) );
  EN U3845 ( .A(n10152), .B(n10660), .Z(n2527) );
  EN U3846 ( .A(n10149), .B(n10660), .Z(n2528) );
  EN U3847 ( .A(n10146), .B(n10660), .Z(n2529) );
  EN U3848 ( .A(n10143), .B(n10660), .Z(n2530) );
  EN U3849 ( .A(n10140), .B(n10660), .Z(n2531) );
  EN U3850 ( .A(n10137), .B(n10659), .Z(n2532) );
  EN U3851 ( .A(n10134), .B(n10659), .Z(n2533) );
  EN U3852 ( .A(n10131), .B(n10659), .Z(n2534) );
  EN U3853 ( .A(n10128), .B(n10659), .Z(n2535) );
  EN U3854 ( .A(n10125), .B(n10659), .Z(n2536) );
  EN U3855 ( .A(n10122), .B(n10659), .Z(n2537) );
  EN U3856 ( .A(n10119), .B(n10659), .Z(n2538) );
  EN U3857 ( .A(n10116), .B(n10659), .Z(n2539) );
  EN U3858 ( .A(n10113), .B(n10659), .Z(n2540) );
  EN U3859 ( .A(n10110), .B(n10659), .Z(n2541) );
  EN U3860 ( .A(n10107), .B(n10659), .Z(n2542) );
  EN U3861 ( .A(n10104), .B(n10659), .Z(n2543) );
  EN U3862 ( .A(n10101), .B(n10659), .Z(n2544) );
  EN U3863 ( .A(n10098), .B(n10659), .Z(n2545) );
  EN U3864 ( .A(n10095), .B(n10658), .Z(n2546) );
  EN U3865 ( .A(n10092), .B(n10658), .Z(n2547) );
  EN U3866 ( .A(n10089), .B(n10658), .Z(n2548) );
  EN U3867 ( .A(n10086), .B(n10658), .Z(n2549) );
  EN U3868 ( .A(n10083), .B(n10658), .Z(n2550) );
  EN U3869 ( .A(n10080), .B(n10658), .Z(n2551) );
  EN U3870 ( .A(n10077), .B(n10658), .Z(n2552) );
  EN U3871 ( .A(n10074), .B(n10658), .Z(n2553) );
  EN U3872 ( .A(n10071), .B(n10658), .Z(n2554) );
  EN U3873 ( .A(n10068), .B(n10658), .Z(n2555) );
  EN U3874 ( .A(n10065), .B(n10658), .Z(n2556) );
  EN U3875 ( .A(n10062), .B(n10658), .Z(n2557) );
  EN U3876 ( .A(n10059), .B(n10658), .Z(n2558) );
  AO4 U3877 ( .A(n10338), .B(n2495), .C(n2496), .D(n10502), .Z(n4653) );
  AO4 U3878 ( .A(n10338), .B(n2496), .C(n2497), .D(n10502), .Z(n4654) );
  AO4 U3879 ( .A(n10338), .B(n2497), .C(n2498), .D(n10502), .Z(n4655) );
  AO4 U3880 ( .A(n10338), .B(n2498), .C(n2499), .D(n10502), .Z(n4656) );
  AO4 U3881 ( .A(n10338), .B(n2499), .C(n2500), .D(n10502), .Z(n4657) );
  AO4 U3882 ( .A(n10338), .B(n2500), .C(n2501), .D(n10502), .Z(n4658) );
  AO4 U3883 ( .A(n10338), .B(n2501), .C(n2502), .D(n10502), .Z(n4659) );
  AO4 U3884 ( .A(n10338), .B(n2502), .C(n2503), .D(n10502), .Z(n4660) );
  AO4 U3885 ( .A(n10338), .B(n2503), .C(n2504), .D(n10502), .Z(n4661) );
  AO4 U3886 ( .A(n10338), .B(n2504), .C(n2505), .D(n10502), .Z(n4662) );
  AO4 U3887 ( .A(n10337), .B(n2505), .C(n2506), .D(n10502), .Z(n4663) );
  AO4 U3888 ( .A(n10337), .B(n2506), .C(n2507), .D(n10501), .Z(n4664) );
  AO4 U3889 ( .A(n10337), .B(n2507), .C(n2508), .D(n10501), .Z(n4665) );
  AO4 U3890 ( .A(n10337), .B(n2508), .C(n2509), .D(n10501), .Z(n4666) );
  AO4 U3891 ( .A(n10337), .B(n2509), .C(n2510), .D(n10501), .Z(n4667) );
  AO4 U3892 ( .A(n10337), .B(n2510), .C(n2511), .D(n10501), .Z(n4668) );
  AO4 U3893 ( .A(n10337), .B(n2511), .C(n2512), .D(n10501), .Z(n4669) );
  AO4 U3894 ( .A(n10337), .B(n2512), .C(n2513), .D(n10501), .Z(n4670) );
  AO4 U3895 ( .A(n10337), .B(n2513), .C(n2514), .D(n10501), .Z(n4671) );
  AO4 U3896 ( .A(n10337), .B(n2514), .C(n2515), .D(n10501), .Z(n4672) );
  AO4 U3897 ( .A(n10337), .B(n2515), .C(n2516), .D(n10501), .Z(n4673) );
  AO4 U3898 ( .A(n10337), .B(n2516), .C(n2517), .D(n10501), .Z(n4674) );
  AO4 U3899 ( .A(n10337), .B(n2517), .C(n2518), .D(n10501), .Z(n4675) );
  AO4 U3900 ( .A(n10337), .B(n2518), .C(n2519), .D(n10501), .Z(n4676) );
  AO4 U3901 ( .A(n10336), .B(n2519), .C(n2520), .D(n10501), .Z(n4677) );
  AO4 U3902 ( .A(n10336), .B(n2520), .C(n2521), .D(n10500), .Z(n4678) );
  AO4 U3903 ( .A(n10336), .B(n2521), .C(n2522), .D(n10500), .Z(n4679) );
  AO4 U3904 ( .A(n10336), .B(n2522), .C(n2523), .D(n10500), .Z(n4680) );
  AO4 U3905 ( .A(n10336), .B(n2523), .C(n2524), .D(n10500), .Z(n4681) );
  AO4 U3906 ( .A(n10336), .B(n2524), .C(n2525), .D(n10500), .Z(n4682) );
  AO4 U3907 ( .A(n10336), .B(n2525), .C(n2526), .D(n10500), .Z(n4683) );
  AO4 U3908 ( .A(n10336), .B(n2526), .C(n2527), .D(n10500), .Z(n4684) );
  AO4 U3909 ( .A(n10336), .B(n2527), .C(n2528), .D(n10500), .Z(n4685) );
  AO4 U3910 ( .A(n10336), .B(n2528), .C(n2529), .D(n10500), .Z(n4686) );
  AO4 U3911 ( .A(n10336), .B(n2529), .C(n2530), .D(n10500), .Z(n4687) );
  AO4 U3912 ( .A(n10336), .B(n2530), .C(n2531), .D(n10500), .Z(n4688) );
  AO4 U3913 ( .A(n10336), .B(n2531), .C(n2532), .D(n10500), .Z(n4689) );
  AO4 U3914 ( .A(n10336), .B(n2532), .C(n2533), .D(n10500), .Z(n4690) );
  AO4 U3915 ( .A(n10335), .B(n2533), .C(n2534), .D(n10500), .Z(n4691) );
  AO4 U3916 ( .A(n10335), .B(n2534), .C(n2535), .D(n10499), .Z(n4692) );
  AO4 U3917 ( .A(n10335), .B(n2535), .C(n2536), .D(n10499), .Z(n4693) );
  AO4 U3918 ( .A(n10335), .B(n2536), .C(n2537), .D(n10499), .Z(n4694) );
  AO4 U3919 ( .A(n10335), .B(n2537), .C(n2538), .D(n10499), .Z(n4695) );
  AO4 U3920 ( .A(n10335), .B(n2538), .C(n2539), .D(n10499), .Z(n4696) );
  AO4 U3921 ( .A(n10335), .B(n2539), .C(n2540), .D(n10499), .Z(n4697) );
  AO4 U3922 ( .A(n10335), .B(n2540), .C(n2541), .D(n10499), .Z(n4698) );
  AO4 U3923 ( .A(n10335), .B(n2541), .C(n2542), .D(n10499), .Z(n4699) );
  AO4 U3924 ( .A(n10335), .B(n2542), .C(n2543), .D(n10499), .Z(n4700) );
  AO4 U3925 ( .A(n10335), .B(n2543), .C(n2544), .D(n10499), .Z(n4701) );
  AO4 U3926 ( .A(n10335), .B(n2544), .C(n2545), .D(n10499), .Z(n4702) );
  AO4 U3927 ( .A(n10335), .B(n2545), .C(n2546), .D(n10499), .Z(n4703) );
  AO4 U3928 ( .A(n10335), .B(n2546), .C(n2547), .D(n10499), .Z(n4704) );
  AO4 U3929 ( .A(n10334), .B(n2547), .C(n2548), .D(n10499), .Z(n4705) );
  AO4 U3930 ( .A(n10334), .B(n2548), .C(n2549), .D(n10498), .Z(n4706) );
  AO4 U3931 ( .A(n10334), .B(n2549), .C(n2550), .D(n10498), .Z(n4707) );
  AO4 U3932 ( .A(n10334), .B(n2550), .C(n2551), .D(n10498), .Z(n4708) );
  AO4 U3933 ( .A(n10334), .B(n2551), .C(n2552), .D(n10498), .Z(n4709) );
  AO4 U3934 ( .A(n10334), .B(n2552), .C(n2553), .D(n10498), .Z(n4710) );
  AO4 U3935 ( .A(n10334), .B(n2553), .C(n2554), .D(n10498), .Z(n4711) );
  AO4 U3936 ( .A(n10334), .B(n2554), .C(n2555), .D(n10498), .Z(n4712) );
  AO4 U3937 ( .A(n10334), .B(n2555), .C(n2556), .D(n10498), .Z(n4713) );
  AO4 U3938 ( .A(n10334), .B(n2556), .C(n2557), .D(n10498), .Z(n4714) );
  AO4 U3939 ( .A(n10334), .B(n2557), .C(n2558), .D(n10498), .Z(n4715) );
  AO4 U3940 ( .A(n10334), .B(n2558), .C(n10498), .D(n1405), .Z(n4716) );
  AO4 U3941 ( .A(n10498), .B(n2494), .C(n10334), .D(n1405), .Z(n5853) );
  EN U3942 ( .A(n10252), .B(n10657), .Z(n2560) );
  EN U3943 ( .A(n10245), .B(n10657), .Z(n2561) );
  EN U3944 ( .A(n10242), .B(n10657), .Z(n2562) );
  EN U3945 ( .A(n10239), .B(n10657), .Z(n2563) );
  EN U3946 ( .A(n10236), .B(n10657), .Z(n2564) );
  EN U3947 ( .A(n10233), .B(n10657), .Z(n2565) );
  EN U3948 ( .A(n10230), .B(n10657), .Z(n2566) );
  EN U3949 ( .A(n10227), .B(n10657), .Z(n2567) );
  EN U3950 ( .A(n10224), .B(n10657), .Z(n2568) );
  EN U3951 ( .A(n10221), .B(n10656), .Z(n2569) );
  EN U3952 ( .A(n10218), .B(n10656), .Z(n2570) );
  EN U3953 ( .A(n10215), .B(n10656), .Z(n2571) );
  EN U3954 ( .A(n10212), .B(n10656), .Z(n2572) );
  EN U3955 ( .A(n10209), .B(n10656), .Z(n2573) );
  EN U3956 ( .A(n10206), .B(n10656), .Z(n2574) );
  EN U3957 ( .A(n10203), .B(n10656), .Z(n2575) );
  EN U3958 ( .A(n10200), .B(n10656), .Z(n2576) );
  EN U3959 ( .A(n10197), .B(n10656), .Z(n2577) );
  EN U3960 ( .A(n10194), .B(n10656), .Z(n2578) );
  EN U3961 ( .A(n10191), .B(n10656), .Z(n2579) );
  EN U3962 ( .A(n10188), .B(n10656), .Z(n2580) );
  EN U3963 ( .A(n10185), .B(n10656), .Z(n2581) );
  EN U3964 ( .A(n10182), .B(n10656), .Z(n2582) );
  EN U3965 ( .A(n10179), .B(n10655), .Z(n2583) );
  EN U3966 ( .A(n10176), .B(n10655), .Z(n2584) );
  EN U3967 ( .A(n10173), .B(n10655), .Z(n2585) );
  EN U3968 ( .A(n10170), .B(n10655), .Z(n2586) );
  EN U3969 ( .A(n10167), .B(n10655), .Z(n2587) );
  EN U3970 ( .A(n10164), .B(n10655), .Z(n2588) );
  EN U3971 ( .A(n10161), .B(n10655), .Z(n2589) );
  EN U3972 ( .A(n10158), .B(n10655), .Z(n2590) );
  EN U3973 ( .A(n10155), .B(n10655), .Z(n2591) );
  EN U3974 ( .A(n10152), .B(n10655), .Z(n2592) );
  EN U3975 ( .A(n10149), .B(n10655), .Z(n2593) );
  EN U3976 ( .A(n10146), .B(n10655), .Z(n2594) );
  EN U3977 ( .A(n10143), .B(n10655), .Z(n2595) );
  EN U3978 ( .A(n10140), .B(n10655), .Z(n2596) );
  EN U3979 ( .A(n10137), .B(n10654), .Z(n2597) );
  EN U3980 ( .A(n10134), .B(n10654), .Z(n2598) );
  EN U3981 ( .A(n10131), .B(n10654), .Z(n2599) );
  EN U3982 ( .A(n10128), .B(n10654), .Z(n2600) );
  EN U3983 ( .A(n10125), .B(n10654), .Z(n2601) );
  EN U3984 ( .A(n10122), .B(n10654), .Z(n2602) );
  EN U3985 ( .A(n10119), .B(n10654), .Z(n2603) );
  EN U3986 ( .A(n10116), .B(n10654), .Z(n2604) );
  EN U3987 ( .A(n10113), .B(n10654), .Z(n2605) );
  EN U3988 ( .A(n10110), .B(n10654), .Z(n2606) );
  EN U3989 ( .A(n10107), .B(n10654), .Z(n2607) );
  EN U3990 ( .A(n10104), .B(n10654), .Z(n2608) );
  EN U3991 ( .A(n10101), .B(n10654), .Z(n2609) );
  EN U3992 ( .A(n10098), .B(n10654), .Z(n2610) );
  EN U3993 ( .A(n10095), .B(n10653), .Z(n2611) );
  EN U3994 ( .A(n10092), .B(n10653), .Z(n2612) );
  EN U3995 ( .A(n10089), .B(n10653), .Z(n2613) );
  EN U3996 ( .A(n10086), .B(n10653), .Z(n2614) );
  EN U3997 ( .A(n10083), .B(n10653), .Z(n2615) );
  EN U3998 ( .A(n10080), .B(n10653), .Z(n2616) );
  EN U3999 ( .A(n10077), .B(n10653), .Z(n2617) );
  EN U4000 ( .A(n10074), .B(n10653), .Z(n2618) );
  EN U4001 ( .A(n10071), .B(n10653), .Z(n2619) );
  EN U4002 ( .A(n10068), .B(n10653), .Z(n2620) );
  EN U4003 ( .A(n10065), .B(n10653), .Z(n2621) );
  EN U4004 ( .A(n10062), .B(n10653), .Z(n2622) );
  EN U4005 ( .A(n10059), .B(n10653), .Z(n2623) );
  AO4 U4006 ( .A(n10333), .B(n2560), .C(n2561), .D(n10497), .Z(n4719) );
  AO4 U4007 ( .A(n10333), .B(n2561), .C(n2562), .D(n10497), .Z(n4720) );
  AO4 U4008 ( .A(n10333), .B(n2562), .C(n2563), .D(n10497), .Z(n4721) );
  AO4 U4009 ( .A(n10333), .B(n2563), .C(n2564), .D(n10497), .Z(n4722) );
  AO4 U4010 ( .A(n10333), .B(n2564), .C(n2565), .D(n10497), .Z(n4723) );
  AO4 U4011 ( .A(n10333), .B(n2565), .C(n2566), .D(n10497), .Z(n4724) );
  AO4 U4012 ( .A(n10333), .B(n2566), .C(n2567), .D(n10497), .Z(n4725) );
  AO4 U4013 ( .A(n10333), .B(n2567), .C(n2568), .D(n10497), .Z(n4726) );
  AO4 U4014 ( .A(n10333), .B(n2568), .C(n2569), .D(n10497), .Z(n4727) );
  AO4 U4015 ( .A(n10333), .B(n2569), .C(n2570), .D(n10497), .Z(n4728) );
  AO4 U4016 ( .A(n10332), .B(n2570), .C(n2571), .D(n10497), .Z(n4729) );
  AO4 U4017 ( .A(n10332), .B(n2571), .C(n2572), .D(n10496), .Z(n4730) );
  AO4 U4018 ( .A(n10332), .B(n2572), .C(n2573), .D(n10496), .Z(n4731) );
  AO4 U4019 ( .A(n10332), .B(n2573), .C(n2574), .D(n10496), .Z(n4732) );
  AO4 U4020 ( .A(n10332), .B(n2574), .C(n2575), .D(n10496), .Z(n4733) );
  AO4 U4021 ( .A(n10332), .B(n2575), .C(n2576), .D(n10496), .Z(n4734) );
  AO4 U4022 ( .A(n10332), .B(n2576), .C(n2577), .D(n10496), .Z(n4735) );
  AO4 U4023 ( .A(n10332), .B(n2577), .C(n2578), .D(n10496), .Z(n4736) );
  AO4 U4024 ( .A(n10332), .B(n2578), .C(n2579), .D(n10496), .Z(n4737) );
  AO4 U4025 ( .A(n10332), .B(n2579), .C(n2580), .D(n10496), .Z(n4738) );
  AO4 U4026 ( .A(n10332), .B(n2580), .C(n2581), .D(n10496), .Z(n4739) );
  AO4 U4027 ( .A(n10332), .B(n2581), .C(n2582), .D(n10496), .Z(n4740) );
  AO4 U4028 ( .A(n10332), .B(n2582), .C(n2583), .D(n10496), .Z(n4741) );
  AO4 U4029 ( .A(n10332), .B(n2583), .C(n2584), .D(n10496), .Z(n4742) );
  AO4 U4030 ( .A(n10331), .B(n2584), .C(n2585), .D(n10496), .Z(n4743) );
  AO4 U4031 ( .A(n10331), .B(n2585), .C(n2586), .D(n10495), .Z(n4744) );
  AO4 U4032 ( .A(n10331), .B(n2586), .C(n2587), .D(n10495), .Z(n4745) );
  AO4 U4033 ( .A(n10331), .B(n2587), .C(n2588), .D(n10495), .Z(n4746) );
  AO4 U4034 ( .A(n10331), .B(n2588), .C(n2589), .D(n10495), .Z(n4747) );
  AO4 U4035 ( .A(n10331), .B(n2589), .C(n2590), .D(n10495), .Z(n4748) );
  AO4 U4036 ( .A(n10331), .B(n2590), .C(n2591), .D(n10495), .Z(n4749) );
  AO4 U4037 ( .A(n10331), .B(n2591), .C(n2592), .D(n10495), .Z(n4750) );
  AO4 U4038 ( .A(n10331), .B(n2592), .C(n2593), .D(n10495), .Z(n4751) );
  AO4 U4039 ( .A(n10331), .B(n2593), .C(n2594), .D(n10495), .Z(n4752) );
  AO4 U4040 ( .A(n10331), .B(n2594), .C(n2595), .D(n10495), .Z(n4753) );
  AO4 U4041 ( .A(n10331), .B(n2595), .C(n2596), .D(n10495), .Z(n4754) );
  AO4 U4042 ( .A(n10331), .B(n2596), .C(n2597), .D(n10495), .Z(n4755) );
  AO4 U4043 ( .A(n10331), .B(n2597), .C(n2598), .D(n10495), .Z(n4756) );
  AO4 U4044 ( .A(n10330), .B(n2598), .C(n2599), .D(n10495), .Z(n4757) );
  AO4 U4045 ( .A(n10330), .B(n2599), .C(n2600), .D(n10494), .Z(n4758) );
  AO4 U4046 ( .A(n10330), .B(n2600), .C(n2601), .D(n10494), .Z(n4759) );
  AO4 U4047 ( .A(n10330), .B(n2601), .C(n2602), .D(n10494), .Z(n4760) );
  AO4 U4048 ( .A(n10330), .B(n2602), .C(n2603), .D(n10494), .Z(n4761) );
  AO4 U4049 ( .A(n10330), .B(n2603), .C(n2604), .D(n10494), .Z(n4762) );
  AO4 U4050 ( .A(n10330), .B(n2604), .C(n2605), .D(n10494), .Z(n4763) );
  AO4 U4051 ( .A(n10330), .B(n2605), .C(n2606), .D(n10494), .Z(n4764) );
  AO4 U4052 ( .A(n10330), .B(n2606), .C(n2607), .D(n10494), .Z(n4765) );
  AO4 U4053 ( .A(n10330), .B(n2607), .C(n2608), .D(n10494), .Z(n4766) );
  AO4 U4054 ( .A(n10330), .B(n2608), .C(n2609), .D(n10494), .Z(n4767) );
  AO4 U4055 ( .A(n10330), .B(n2609), .C(n2610), .D(n10494), .Z(n4768) );
  AO4 U4056 ( .A(n10330), .B(n2610), .C(n2611), .D(n10494), .Z(n4769) );
  AO4 U4057 ( .A(n10330), .B(n2611), .C(n2612), .D(n10494), .Z(n4770) );
  AO4 U4058 ( .A(n10329), .B(n2612), .C(n2613), .D(n10494), .Z(n4771) );
  AO4 U4059 ( .A(n10329), .B(n2613), .C(n2614), .D(n10493), .Z(n4772) );
  AO4 U4060 ( .A(n10329), .B(n2614), .C(n2615), .D(n10493), .Z(n4773) );
  AO4 U4061 ( .A(n10329), .B(n2615), .C(n2616), .D(n10493), .Z(n4774) );
  AO4 U4062 ( .A(n10329), .B(n2616), .C(n2617), .D(n10493), .Z(n4775) );
  AO4 U4063 ( .A(n10329), .B(n2617), .C(n2618), .D(n10493), .Z(n4776) );
  AO4 U4064 ( .A(n10329), .B(n2618), .C(n2619), .D(n10493), .Z(n4777) );
  AO4 U4065 ( .A(n10329), .B(n2619), .C(n2620), .D(n10493), .Z(n4778) );
  AO4 U4066 ( .A(n10329), .B(n2620), .C(n2621), .D(n10493), .Z(n4779) );
  AO4 U4067 ( .A(n10329), .B(n2621), .C(n2622), .D(n10493), .Z(n4780) );
  AO4 U4068 ( .A(n10329), .B(n2622), .C(n2623), .D(n10493), .Z(n4781) );
  AO4 U4069 ( .A(n10329), .B(n2623), .C(n10493), .D(n1406), .Z(n4782) );
  AO4 U4070 ( .A(n10493), .B(n2559), .C(n10329), .D(n1406), .Z(n5854) );
  EN U4071 ( .A(n10252), .B(n10652), .Z(n2625) );
  EN U4072 ( .A(n10245), .B(n10652), .Z(n2626) );
  EN U4073 ( .A(n10242), .B(n10652), .Z(n2627) );
  EN U4074 ( .A(n10239), .B(n10652), .Z(n2628) );
  EN U4075 ( .A(n10236), .B(n10652), .Z(n2629) );
  EN U4076 ( .A(n10233), .B(n10652), .Z(n2630) );
  EN U4077 ( .A(n10230), .B(n10652), .Z(n2631) );
  EN U4078 ( .A(n10227), .B(n10652), .Z(n2632) );
  EN U4079 ( .A(n10224), .B(n10652), .Z(n2633) );
  EN U4080 ( .A(n10221), .B(n10651), .Z(n2634) );
  EN U4081 ( .A(n10218), .B(n10651), .Z(n2635) );
  EN U4082 ( .A(n10215), .B(n10651), .Z(n2636) );
  EN U4083 ( .A(n10212), .B(n10651), .Z(n2637) );
  EN U4084 ( .A(n10209), .B(n10651), .Z(n2638) );
  EN U4085 ( .A(n10206), .B(n10651), .Z(n2639) );
  EN U4086 ( .A(n10203), .B(n10651), .Z(n2640) );
  EN U4087 ( .A(n10200), .B(n10651), .Z(n2641) );
  EN U4088 ( .A(n10197), .B(n10651), .Z(n2642) );
  EN U4089 ( .A(n10194), .B(n10651), .Z(n2643) );
  EN U4090 ( .A(n10191), .B(n10651), .Z(n2644) );
  EN U4091 ( .A(n10188), .B(n10651), .Z(n2645) );
  EN U4092 ( .A(n10185), .B(n10651), .Z(n2646) );
  EN U4093 ( .A(n10182), .B(n10651), .Z(n2647) );
  EN U4094 ( .A(n10179), .B(n10650), .Z(n2648) );
  EN U4095 ( .A(n10176), .B(n10650), .Z(n2649) );
  EN U4096 ( .A(n10173), .B(n10650), .Z(n2650) );
  EN U4097 ( .A(n10170), .B(n10650), .Z(n2651) );
  EN U4098 ( .A(n10167), .B(n10650), .Z(n2652) );
  EN U4099 ( .A(n10164), .B(n10650), .Z(n2653) );
  EN U4100 ( .A(n10161), .B(n10650), .Z(n2654) );
  EN U4101 ( .A(n10158), .B(n10650), .Z(n2655) );
  EN U4102 ( .A(n10155), .B(n10650), .Z(n2656) );
  EN U4103 ( .A(n10152), .B(n10650), .Z(n2657) );
  EN U4104 ( .A(n10149), .B(n10650), .Z(n2658) );
  EN U4105 ( .A(n10146), .B(n10650), .Z(n2659) );
  EN U4106 ( .A(n10143), .B(n10650), .Z(n2660) );
  EN U4107 ( .A(n10140), .B(n10650), .Z(n2661) );
  EN U4108 ( .A(n10137), .B(n10649), .Z(n2662) );
  EN U4109 ( .A(n10134), .B(n10649), .Z(n2663) );
  EN U4110 ( .A(n10131), .B(n10649), .Z(n2664) );
  EN U4111 ( .A(n10128), .B(n10649), .Z(n2665) );
  EN U4112 ( .A(n10125), .B(n10649), .Z(n2666) );
  EN U4113 ( .A(n10122), .B(n10649), .Z(n2667) );
  EN U4114 ( .A(n10119), .B(n10649), .Z(n2668) );
  EN U4115 ( .A(n10116), .B(n10649), .Z(n2669) );
  EN U4116 ( .A(n10113), .B(n10649), .Z(n2670) );
  EN U4117 ( .A(n10110), .B(n10649), .Z(n2671) );
  EN U4118 ( .A(n10107), .B(n10649), .Z(n2672) );
  EN U4119 ( .A(n10104), .B(n10649), .Z(n2673) );
  EN U4120 ( .A(n10101), .B(n10649), .Z(n2674) );
  EN U4121 ( .A(n10098), .B(n10649), .Z(n2675) );
  EN U4122 ( .A(n10095), .B(n10648), .Z(n2676) );
  EN U4123 ( .A(n10092), .B(n10648), .Z(n2677) );
  EN U4124 ( .A(n10089), .B(n10648), .Z(n2678) );
  EN U4125 ( .A(n10086), .B(n10648), .Z(n2679) );
  EN U4126 ( .A(n10083), .B(n10648), .Z(n2680) );
  EN U4127 ( .A(n10080), .B(n10648), .Z(n2681) );
  EN U4128 ( .A(n10077), .B(n10648), .Z(n2682) );
  EN U4129 ( .A(n10074), .B(n10648), .Z(n2683) );
  EN U4130 ( .A(n10071), .B(n10648), .Z(n2684) );
  EN U4131 ( .A(n10068), .B(n10648), .Z(n2685) );
  EN U4132 ( .A(n10065), .B(n10648), .Z(n2686) );
  EN U4133 ( .A(n10062), .B(n10648), .Z(n2687) );
  EN U4134 ( .A(n10059), .B(n10648), .Z(n2688) );
  AO4 U4135 ( .A(n10328), .B(n2625), .C(n2626), .D(n10492), .Z(n4785) );
  AO4 U4136 ( .A(n10328), .B(n2626), .C(n2627), .D(n10492), .Z(n4786) );
  AO4 U4137 ( .A(n10328), .B(n2627), .C(n2628), .D(n10492), .Z(n4787) );
  AO4 U4138 ( .A(n10328), .B(n2628), .C(n2629), .D(n10492), .Z(n4788) );
  AO4 U4139 ( .A(n10328), .B(n2629), .C(n2630), .D(n10492), .Z(n4789) );
  AO4 U4140 ( .A(n10328), .B(n2630), .C(n2631), .D(n10492), .Z(n4790) );
  AO4 U4141 ( .A(n10328), .B(n2631), .C(n2632), .D(n10492), .Z(n4791) );
  AO4 U4142 ( .A(n10328), .B(n2632), .C(n2633), .D(n10492), .Z(n4792) );
  AO4 U4143 ( .A(n10328), .B(n2633), .C(n2634), .D(n10492), .Z(n4793) );
  AO4 U4144 ( .A(n10328), .B(n2634), .C(n2635), .D(n10492), .Z(n4794) );
  AO4 U4145 ( .A(n10327), .B(n2635), .C(n2636), .D(n10492), .Z(n4795) );
  AO4 U4146 ( .A(n10327), .B(n2636), .C(n2637), .D(n10491), .Z(n4796) );
  AO4 U4147 ( .A(n10327), .B(n2637), .C(n2638), .D(n10491), .Z(n4797) );
  AO4 U4148 ( .A(n10327), .B(n2638), .C(n2639), .D(n10491), .Z(n4798) );
  AO4 U4149 ( .A(n10327), .B(n2639), .C(n2640), .D(n10491), .Z(n4799) );
  AO4 U4150 ( .A(n10327), .B(n2640), .C(n2641), .D(n10491), .Z(n4800) );
  AO4 U4151 ( .A(n10327), .B(n2641), .C(n2642), .D(n10491), .Z(n4801) );
  AO4 U4152 ( .A(n10327), .B(n2642), .C(n2643), .D(n10491), .Z(n4802) );
  AO4 U4153 ( .A(n10327), .B(n2643), .C(n2644), .D(n10491), .Z(n4803) );
  AO4 U4154 ( .A(n10327), .B(n2644), .C(n2645), .D(n10491), .Z(n4804) );
  AO4 U4155 ( .A(n10327), .B(n2645), .C(n2646), .D(n10491), .Z(n4805) );
  AO4 U4156 ( .A(n10327), .B(n2646), .C(n2647), .D(n10491), .Z(n4806) );
  AO4 U4157 ( .A(n10327), .B(n2647), .C(n2648), .D(n10491), .Z(n4807) );
  AO4 U4158 ( .A(n10327), .B(n2648), .C(n2649), .D(n10491), .Z(n4808) );
  AO4 U4159 ( .A(n10326), .B(n2649), .C(n2650), .D(n10491), .Z(n4809) );
  AO4 U4160 ( .A(n10326), .B(n2650), .C(n2651), .D(n10490), .Z(n4810) );
  AO4 U4161 ( .A(n10326), .B(n2651), .C(n2652), .D(n10490), .Z(n4811) );
  AO4 U4162 ( .A(n10326), .B(n2652), .C(n2653), .D(n10490), .Z(n4812) );
  AO4 U4163 ( .A(n10326), .B(n2653), .C(n2654), .D(n10490), .Z(n4813) );
  AO4 U4164 ( .A(n10326), .B(n2654), .C(n2655), .D(n10490), .Z(n4814) );
  AO4 U4165 ( .A(n10326), .B(n2655), .C(n2656), .D(n10490), .Z(n4815) );
  AO4 U4166 ( .A(n10326), .B(n2656), .C(n2657), .D(n10490), .Z(n4816) );
  AO4 U4167 ( .A(n10326), .B(n2657), .C(n2658), .D(n10490), .Z(n4817) );
  AO4 U4168 ( .A(n10326), .B(n2658), .C(n2659), .D(n10490), .Z(n4818) );
  AO4 U4169 ( .A(n10326), .B(n2659), .C(n2660), .D(n10490), .Z(n4819) );
  AO4 U4170 ( .A(n10326), .B(n2660), .C(n2661), .D(n10490), .Z(n4820) );
  AO4 U4171 ( .A(n10326), .B(n2661), .C(n2662), .D(n10490), .Z(n4821) );
  AO4 U4172 ( .A(n10326), .B(n2662), .C(n2663), .D(n10490), .Z(n4822) );
  AO4 U4173 ( .A(n10325), .B(n2663), .C(n2664), .D(n10490), .Z(n4823) );
  AO4 U4174 ( .A(n10325), .B(n2664), .C(n2665), .D(n10489), .Z(n4824) );
  AO4 U4175 ( .A(n10325), .B(n2665), .C(n2666), .D(n10489), .Z(n4825) );
  AO4 U4176 ( .A(n10325), .B(n2666), .C(n2667), .D(n10489), .Z(n4826) );
  AO4 U4177 ( .A(n10325), .B(n2667), .C(n2668), .D(n10489), .Z(n4827) );
  AO4 U4178 ( .A(n10325), .B(n2668), .C(n2669), .D(n10489), .Z(n4828) );
  AO4 U4179 ( .A(n10325), .B(n2669), .C(n2670), .D(n10489), .Z(n4829) );
  AO4 U4180 ( .A(n10325), .B(n2670), .C(n2671), .D(n10489), .Z(n4830) );
  AO4 U4181 ( .A(n10325), .B(n2671), .C(n2672), .D(n10489), .Z(n4831) );
  AO4 U4182 ( .A(n10325), .B(n2672), .C(n2673), .D(n10489), .Z(n4832) );
  AO4 U4183 ( .A(n10325), .B(n2673), .C(n2674), .D(n10489), .Z(n4833) );
  AO4 U4184 ( .A(n10325), .B(n2674), .C(n2675), .D(n10489), .Z(n4834) );
  AO4 U4185 ( .A(n10325), .B(n2675), .C(n2676), .D(n10489), .Z(n4835) );
  AO4 U4186 ( .A(n10325), .B(n2676), .C(n2677), .D(n10489), .Z(n4836) );
  AO4 U4187 ( .A(n10324), .B(n2677), .C(n2678), .D(n10489), .Z(n4837) );
  AO4 U4188 ( .A(n10324), .B(n2678), .C(n2679), .D(n10488), .Z(n4838) );
  AO4 U4189 ( .A(n10324), .B(n2679), .C(n2680), .D(n10488), .Z(n4839) );
  AO4 U4190 ( .A(n10324), .B(n2680), .C(n2681), .D(n10488), .Z(n4840) );
  AO4 U4191 ( .A(n10324), .B(n2681), .C(n2682), .D(n10488), .Z(n4841) );
  AO4 U4192 ( .A(n10324), .B(n2682), .C(n2683), .D(n10488), .Z(n4842) );
  AO4 U4193 ( .A(n10324), .B(n2683), .C(n2684), .D(n10488), .Z(n4843) );
  AO4 U4194 ( .A(n10324), .B(n2684), .C(n2685), .D(n10488), .Z(n4844) );
  AO4 U4195 ( .A(n10324), .B(n2685), .C(n2686), .D(n10488), .Z(n4845) );
  AO4 U4196 ( .A(n10324), .B(n2686), .C(n2687), .D(n10488), .Z(n4846) );
  AO4 U4197 ( .A(n10324), .B(n2687), .C(n2688), .D(n10488), .Z(n4847) );
  AO4 U4198 ( .A(n10324), .B(n2688), .C(n10488), .D(n1407), .Z(n4848) );
  AO4 U4199 ( .A(n10488), .B(n2624), .C(n10324), .D(n1407), .Z(n5855) );
  EN U4200 ( .A(n10252), .B(n10647), .Z(n2690) );
  EN U4201 ( .A(n10245), .B(n10647), .Z(n2691) );
  EN U4202 ( .A(n10242), .B(n10647), .Z(n2692) );
  EN U4203 ( .A(n10239), .B(n10647), .Z(n2693) );
  EN U4204 ( .A(n10236), .B(n10647), .Z(n2694) );
  EN U4205 ( .A(n10233), .B(n10647), .Z(n2695) );
  EN U4206 ( .A(n10230), .B(n10647), .Z(n2696) );
  EN U4207 ( .A(n10227), .B(n10647), .Z(n2697) );
  EN U4208 ( .A(n10224), .B(n10647), .Z(n2698) );
  EN U4209 ( .A(n10221), .B(n10646), .Z(n2699) );
  EN U4210 ( .A(n10218), .B(n10646), .Z(n2700) );
  EN U4211 ( .A(n10215), .B(n10646), .Z(n2701) );
  EN U4212 ( .A(n10212), .B(n10646), .Z(n2702) );
  EN U4213 ( .A(n10209), .B(n10646), .Z(n2703) );
  EN U4214 ( .A(n10206), .B(n10646), .Z(n2704) );
  EN U4215 ( .A(n10203), .B(n10646), .Z(n2705) );
  EN U4216 ( .A(n10200), .B(n10646), .Z(n2706) );
  EN U4217 ( .A(n10197), .B(n10646), .Z(n2707) );
  EN U4218 ( .A(n10194), .B(n10646), .Z(n2708) );
  EN U4219 ( .A(n10191), .B(n10646), .Z(n2709) );
  EN U4220 ( .A(n10188), .B(n10646), .Z(n2710) );
  EN U4221 ( .A(n10185), .B(n10646), .Z(n2711) );
  EN U4222 ( .A(n10182), .B(n10646), .Z(n2712) );
  EN U4223 ( .A(n10179), .B(n10645), .Z(n2713) );
  EN U4224 ( .A(n10176), .B(n10645), .Z(n2714) );
  EN U4225 ( .A(n10173), .B(n10645), .Z(n2715) );
  EN U4226 ( .A(n10170), .B(n10645), .Z(n2716) );
  EN U4227 ( .A(n10167), .B(n10645), .Z(n2717) );
  EN U4228 ( .A(n10164), .B(n10645), .Z(n2718) );
  EN U4229 ( .A(n10161), .B(n10645), .Z(n2719) );
  EN U4230 ( .A(n10158), .B(n10645), .Z(n2720) );
  EN U4231 ( .A(n10155), .B(n10645), .Z(n2721) );
  EN U4232 ( .A(n10152), .B(n10645), .Z(n2722) );
  EN U4233 ( .A(n10149), .B(n10645), .Z(n2723) );
  EN U4234 ( .A(n10146), .B(n10645), .Z(n2724) );
  EN U4235 ( .A(n10143), .B(n10645), .Z(n2725) );
  EN U4236 ( .A(n10140), .B(n10645), .Z(n2726) );
  EN U4237 ( .A(n10137), .B(n10644), .Z(n2727) );
  EN U4238 ( .A(n10134), .B(n10644), .Z(n2728) );
  EN U4239 ( .A(n10131), .B(n10644), .Z(n2729) );
  EN U4240 ( .A(n10128), .B(n10644), .Z(n2730) );
  EN U4241 ( .A(n10125), .B(n10644), .Z(n2731) );
  EN U4242 ( .A(n10122), .B(n10644), .Z(n2732) );
  EN U4243 ( .A(n10119), .B(n10644), .Z(n2733) );
  EN U4244 ( .A(n10116), .B(n10644), .Z(n2734) );
  EN U4245 ( .A(n10113), .B(n10644), .Z(n2735) );
  EN U4246 ( .A(n10110), .B(n10644), .Z(n2736) );
  EN U4247 ( .A(n10107), .B(n10644), .Z(n2737) );
  EN U4248 ( .A(n10104), .B(n10644), .Z(n2738) );
  EN U4249 ( .A(n10101), .B(n10644), .Z(n2739) );
  EN U4250 ( .A(n10098), .B(n10644), .Z(n2740) );
  EN U4251 ( .A(n10095), .B(n10643), .Z(n2741) );
  EN U4252 ( .A(n10092), .B(n10643), .Z(n2742) );
  EN U4253 ( .A(n10089), .B(n10643), .Z(n2743) );
  EN U4254 ( .A(n10086), .B(n10643), .Z(n2744) );
  EN U4255 ( .A(n10083), .B(n10643), .Z(n2745) );
  EN U4256 ( .A(n10080), .B(n10643), .Z(n2746) );
  EN U4257 ( .A(n10077), .B(n10643), .Z(n2747) );
  EN U4258 ( .A(n10074), .B(n10643), .Z(n2748) );
  EN U4259 ( .A(n10071), .B(n10643), .Z(n2749) );
  EN U4260 ( .A(n10068), .B(n10643), .Z(n2750) );
  EN U4261 ( .A(n10065), .B(n10643), .Z(n2751) );
  EN U4262 ( .A(n10062), .B(n10643), .Z(n2752) );
  EN U4263 ( .A(n10059), .B(n10643), .Z(n2753) );
  AO4 U4264 ( .A(n10323), .B(n2690), .C(n2691), .D(n10487), .Z(n4851) );
  AO4 U4265 ( .A(n10323), .B(n2691), .C(n2692), .D(n10487), .Z(n4852) );
  AO4 U4266 ( .A(n10323), .B(n2692), .C(n2693), .D(n10487), .Z(n4853) );
  AO4 U4267 ( .A(n10323), .B(n2693), .C(n2694), .D(n10487), .Z(n4854) );
  AO4 U4268 ( .A(n10323), .B(n2694), .C(n2695), .D(n10487), .Z(n4855) );
  AO4 U4269 ( .A(n10323), .B(n2695), .C(n2696), .D(n10487), .Z(n4856) );
  AO4 U4270 ( .A(n10323), .B(n2696), .C(n2697), .D(n10487), .Z(n4857) );
  AO4 U4271 ( .A(n10323), .B(n2697), .C(n2698), .D(n10487), .Z(n4858) );
  AO4 U4272 ( .A(n10323), .B(n2698), .C(n2699), .D(n10487), .Z(n4859) );
  AO4 U4273 ( .A(n10323), .B(n2699), .C(n2700), .D(n10487), .Z(n4860) );
  AO4 U4274 ( .A(n10322), .B(n2700), .C(n2701), .D(n10487), .Z(n4861) );
  AO4 U4275 ( .A(n10322), .B(n2701), .C(n2702), .D(n10486), .Z(n4862) );
  AO4 U4276 ( .A(n10322), .B(n2702), .C(n2703), .D(n10486), .Z(n4863) );
  AO4 U4277 ( .A(n10322), .B(n2703), .C(n2704), .D(n10486), .Z(n4864) );
  AO4 U4278 ( .A(n10322), .B(n2704), .C(n2705), .D(n10486), .Z(n4865) );
  AO4 U4279 ( .A(n10322), .B(n2705), .C(n2706), .D(n10486), .Z(n4866) );
  AO4 U4280 ( .A(n10322), .B(n2706), .C(n2707), .D(n10486), .Z(n4867) );
  AO4 U4281 ( .A(n10322), .B(n2707), .C(n2708), .D(n10486), .Z(n4868) );
  AO4 U4282 ( .A(n10322), .B(n2708), .C(n2709), .D(n10486), .Z(n4869) );
  AO4 U4283 ( .A(n10322), .B(n2709), .C(n2710), .D(n10486), .Z(n4870) );
  AO4 U4284 ( .A(n10322), .B(n2710), .C(n2711), .D(n10486), .Z(n4871) );
  AO4 U4285 ( .A(n10322), .B(n2711), .C(n2712), .D(n10486), .Z(n4872) );
  AO4 U4286 ( .A(n10322), .B(n2712), .C(n2713), .D(n10486), .Z(n4873) );
  AO4 U4287 ( .A(n10322), .B(n2713), .C(n2714), .D(n10486), .Z(n4874) );
  AO4 U4288 ( .A(n10321), .B(n2714), .C(n2715), .D(n10486), .Z(n4875) );
  AO4 U4289 ( .A(n10321), .B(n2715), .C(n2716), .D(n10485), .Z(n4876) );
  AO4 U4290 ( .A(n10321), .B(n2716), .C(n2717), .D(n10485), .Z(n4877) );
  AO4 U4291 ( .A(n10321), .B(n2717), .C(n2718), .D(n10485), .Z(n4878) );
  AO4 U4292 ( .A(n10321), .B(n2718), .C(n2719), .D(n10485), .Z(n4879) );
  AO4 U4293 ( .A(n10321), .B(n2719), .C(n2720), .D(n10485), .Z(n4880) );
  AO4 U4294 ( .A(n10321), .B(n2720), .C(n2721), .D(n10485), .Z(n4881) );
  AO4 U4295 ( .A(n10321), .B(n2721), .C(n2722), .D(n10485), .Z(n4882) );
  AO4 U4296 ( .A(n10321), .B(n2722), .C(n2723), .D(n10485), .Z(n4883) );
  AO4 U4297 ( .A(n10321), .B(n2723), .C(n2724), .D(n10485), .Z(n4884) );
  AO4 U4298 ( .A(n10321), .B(n2724), .C(n2725), .D(n10485), .Z(n4885) );
  AO4 U4299 ( .A(n10321), .B(n2725), .C(n2726), .D(n10485), .Z(n4886) );
  AO4 U4300 ( .A(n10321), .B(n2726), .C(n2727), .D(n10485), .Z(n4887) );
  AO4 U4301 ( .A(n10321), .B(n2727), .C(n2728), .D(n10485), .Z(n4888) );
  AO4 U4302 ( .A(n10320), .B(n2728), .C(n2729), .D(n10485), .Z(n4889) );
  AO4 U4303 ( .A(n10320), .B(n2729), .C(n2730), .D(n10484), .Z(n4890) );
  AO4 U4304 ( .A(n10320), .B(n2730), .C(n2731), .D(n10484), .Z(n4891) );
  AO4 U4305 ( .A(n10320), .B(n2731), .C(n2732), .D(n10484), .Z(n4892) );
  AO4 U4306 ( .A(n10320), .B(n2732), .C(n2733), .D(n10484), .Z(n4893) );
  AO4 U4307 ( .A(n10320), .B(n2733), .C(n2734), .D(n10484), .Z(n4894) );
  AO4 U4308 ( .A(n10320), .B(n2734), .C(n2735), .D(n10484), .Z(n4895) );
  AO4 U4309 ( .A(n10320), .B(n2735), .C(n2736), .D(n10484), .Z(n4896) );
  AO4 U4310 ( .A(n10320), .B(n2736), .C(n2737), .D(n10484), .Z(n4897) );
  AO4 U4311 ( .A(n10320), .B(n2737), .C(n2738), .D(n10484), .Z(n4898) );
  AO4 U4312 ( .A(n10320), .B(n2738), .C(n2739), .D(n10484), .Z(n4899) );
  AO4 U4313 ( .A(n10320), .B(n2739), .C(n2740), .D(n10484), .Z(n4900) );
  AO4 U4314 ( .A(n10320), .B(n2740), .C(n2741), .D(n10484), .Z(n4901) );
  AO4 U4315 ( .A(n10320), .B(n2741), .C(n2742), .D(n10484), .Z(n4902) );
  AO4 U4316 ( .A(n10319), .B(n2742), .C(n2743), .D(n10484), .Z(n4903) );
  AO4 U4317 ( .A(n10319), .B(n2743), .C(n2744), .D(n10483), .Z(n4904) );
  AO4 U4318 ( .A(n10319), .B(n2744), .C(n2745), .D(n10483), .Z(n4905) );
  AO4 U4319 ( .A(n10319), .B(n2745), .C(n2746), .D(n10483), .Z(n4906) );
  AO4 U4320 ( .A(n10319), .B(n2746), .C(n2747), .D(n10483), .Z(n4907) );
  AO4 U4321 ( .A(n10319), .B(n2747), .C(n2748), .D(n10483), .Z(n4908) );
  AO4 U4322 ( .A(n10319), .B(n2748), .C(n2749), .D(n10483), .Z(n4909) );
  AO4 U4323 ( .A(n10319), .B(n2749), .C(n2750), .D(n10483), .Z(n4910) );
  AO4 U4324 ( .A(n10319), .B(n2750), .C(n2751), .D(n10483), .Z(n4911) );
  AO4 U4325 ( .A(n10319), .B(n2751), .C(n2752), .D(n10483), .Z(n4912) );
  AO4 U4326 ( .A(n10319), .B(n2752), .C(n2753), .D(n10483), .Z(n4913) );
  AO4 U4327 ( .A(n10319), .B(n2753), .C(n10483), .D(n1408), .Z(n4914) );
  AO4 U4328 ( .A(n10483), .B(n2689), .C(n10319), .D(n1408), .Z(n5856) );
  EN U4329 ( .A(n10252), .B(n10642), .Z(n2755) );
  EN U4330 ( .A(n10245), .B(n10642), .Z(n2756) );
  EN U4331 ( .A(n10242), .B(n10642), .Z(n2757) );
  EN U4332 ( .A(n10239), .B(n10642), .Z(n2758) );
  EN U4333 ( .A(n10236), .B(n10642), .Z(n2759) );
  EN U4334 ( .A(n10233), .B(n10642), .Z(n2760) );
  EN U4335 ( .A(n10230), .B(n10642), .Z(n2761) );
  EN U4336 ( .A(n10227), .B(n10642), .Z(n2762) );
  EN U4337 ( .A(n10224), .B(n10642), .Z(n2763) );
  EN U4338 ( .A(n10221), .B(n10641), .Z(n2764) );
  EN U4339 ( .A(n10218), .B(n10641), .Z(n2765) );
  EN U4340 ( .A(n10215), .B(n10641), .Z(n2766) );
  EN U4341 ( .A(n10212), .B(n10641), .Z(n2767) );
  EN U4342 ( .A(n10209), .B(n10641), .Z(n2768) );
  EN U4343 ( .A(n10206), .B(n10641), .Z(n2769) );
  EN U4344 ( .A(n10203), .B(n10641), .Z(n2770) );
  EN U4345 ( .A(n10200), .B(n10641), .Z(n2771) );
  EN U4346 ( .A(n10197), .B(n10641), .Z(n2772) );
  EN U4347 ( .A(n10194), .B(n10641), .Z(n2773) );
  EN U4348 ( .A(n10191), .B(n10641), .Z(n2774) );
  EN U4349 ( .A(n10188), .B(n10641), .Z(n2775) );
  EN U4350 ( .A(n10185), .B(n10641), .Z(n2776) );
  EN U4351 ( .A(n10182), .B(n10641), .Z(n2777) );
  EN U4352 ( .A(n10179), .B(n10640), .Z(n2778) );
  EN U4353 ( .A(n10176), .B(n10640), .Z(n2779) );
  EN U4354 ( .A(n10173), .B(n10640), .Z(n2780) );
  EN U4355 ( .A(n10170), .B(n10640), .Z(n2781) );
  EN U4356 ( .A(n10167), .B(n10640), .Z(n2782) );
  EN U4357 ( .A(n10164), .B(n10640), .Z(n2783) );
  EN U4358 ( .A(n10161), .B(n10640), .Z(n2784) );
  EN U4359 ( .A(n10158), .B(n10640), .Z(n2785) );
  EN U4360 ( .A(n10155), .B(n10640), .Z(n2786) );
  EN U4361 ( .A(n10152), .B(n10640), .Z(n2787) );
  EN U4362 ( .A(n10149), .B(n10640), .Z(n2788) );
  EN U4363 ( .A(n10146), .B(n10640), .Z(n2789) );
  EN U4364 ( .A(n10143), .B(n10640), .Z(n2790) );
  EN U4365 ( .A(n10140), .B(n10640), .Z(n2791) );
  EN U4366 ( .A(n10137), .B(n10639), .Z(n2792) );
  EN U4367 ( .A(n10134), .B(n10639), .Z(n2793) );
  EN U4368 ( .A(n10131), .B(n10639), .Z(n2794) );
  EN U4369 ( .A(n10128), .B(n10639), .Z(n2795) );
  EN U4370 ( .A(n10125), .B(n10639), .Z(n2796) );
  EN U4371 ( .A(n10122), .B(n10639), .Z(n2797) );
  EN U4372 ( .A(n10119), .B(n10639), .Z(n2798) );
  EN U4373 ( .A(n10116), .B(n10639), .Z(n2799) );
  EN U4374 ( .A(n10113), .B(n10639), .Z(n2800) );
  EN U4375 ( .A(n10110), .B(n10639), .Z(n2801) );
  EN U4376 ( .A(n10107), .B(n10639), .Z(n2802) );
  EN U4377 ( .A(n10104), .B(n10639), .Z(n2803) );
  EN U4378 ( .A(n10101), .B(n10639), .Z(n2804) );
  EN U4379 ( .A(n10098), .B(n10639), .Z(n2805) );
  EN U4380 ( .A(n10095), .B(n10638), .Z(n2806) );
  EN U4381 ( .A(n10092), .B(n10638), .Z(n2807) );
  EN U4382 ( .A(n10089), .B(n10638), .Z(n2808) );
  EN U4383 ( .A(n10086), .B(n10638), .Z(n2809) );
  EN U4384 ( .A(n10083), .B(n10638), .Z(n2810) );
  EN U4385 ( .A(n10080), .B(n10638), .Z(n2811) );
  EN U4386 ( .A(n10077), .B(n10638), .Z(n2812) );
  EN U4387 ( .A(n10074), .B(n10638), .Z(n2813) );
  EN U4388 ( .A(n10071), .B(n10638), .Z(n2814) );
  EN U4389 ( .A(n10068), .B(n10638), .Z(n2815) );
  EN U4390 ( .A(n10065), .B(n10638), .Z(n2816) );
  EN U4391 ( .A(n10062), .B(n10638), .Z(n2817) );
  EN U4392 ( .A(n10059), .B(n10638), .Z(n2818) );
  AO4 U4393 ( .A(n10318), .B(n2755), .C(n2756), .D(n10482), .Z(n4917) );
  AO4 U4394 ( .A(n10318), .B(n2756), .C(n2757), .D(n10482), .Z(n4918) );
  AO4 U4395 ( .A(n10318), .B(n2757), .C(n2758), .D(n10482), .Z(n4919) );
  AO4 U4396 ( .A(n10318), .B(n2758), .C(n2759), .D(n10482), .Z(n4920) );
  AO4 U4397 ( .A(n10318), .B(n2759), .C(n2760), .D(n10482), .Z(n4921) );
  AO4 U4398 ( .A(n10318), .B(n2760), .C(n2761), .D(n10482), .Z(n4922) );
  AO4 U4399 ( .A(n10318), .B(n2761), .C(n2762), .D(n10482), .Z(n4923) );
  AO4 U4400 ( .A(n10318), .B(n2762), .C(n2763), .D(n10482), .Z(n4924) );
  AO4 U4401 ( .A(n10318), .B(n2763), .C(n2764), .D(n10482), .Z(n4925) );
  AO4 U4402 ( .A(n10318), .B(n2764), .C(n2765), .D(n10482), .Z(n4926) );
  AO4 U4403 ( .A(n10317), .B(n2765), .C(n2766), .D(n10482), .Z(n4927) );
  AO4 U4404 ( .A(n10317), .B(n2766), .C(n2767), .D(n10481), .Z(n4928) );
  AO4 U4405 ( .A(n10317), .B(n2767), .C(n2768), .D(n10481), .Z(n4929) );
  AO4 U4406 ( .A(n10317), .B(n2768), .C(n2769), .D(n10481), .Z(n4930) );
  AO4 U4407 ( .A(n10317), .B(n2769), .C(n2770), .D(n10481), .Z(n4931) );
  AO4 U4408 ( .A(n10317), .B(n2770), .C(n2771), .D(n10481), .Z(n4932) );
  AO4 U4409 ( .A(n10317), .B(n2771), .C(n2772), .D(n10481), .Z(n4933) );
  AO4 U4410 ( .A(n10317), .B(n2772), .C(n2773), .D(n10481), .Z(n4934) );
  AO4 U4411 ( .A(n10317), .B(n2773), .C(n2774), .D(n10481), .Z(n4935) );
  AO4 U4412 ( .A(n10317), .B(n2774), .C(n2775), .D(n10481), .Z(n4936) );
  AO4 U4413 ( .A(n10317), .B(n2775), .C(n2776), .D(n10481), .Z(n4937) );
  AO4 U4414 ( .A(n10317), .B(n2776), .C(n2777), .D(n10481), .Z(n4938) );
  AO4 U4415 ( .A(n10317), .B(n2777), .C(n2778), .D(n10481), .Z(n4939) );
  AO4 U4416 ( .A(n10317), .B(n2778), .C(n2779), .D(n10481), .Z(n4940) );
  AO4 U4417 ( .A(n10316), .B(n2779), .C(n2780), .D(n10481), .Z(n4941) );
  AO4 U4418 ( .A(n10316), .B(n2780), .C(n2781), .D(n10480), .Z(n4942) );
  AO4 U4419 ( .A(n10316), .B(n2781), .C(n2782), .D(n10480), .Z(n4943) );
  AO4 U4420 ( .A(n10316), .B(n2782), .C(n2783), .D(n10480), .Z(n4944) );
  AO4 U4421 ( .A(n10316), .B(n2783), .C(n2784), .D(n10480), .Z(n4945) );
  AO4 U4422 ( .A(n10316), .B(n2784), .C(n2785), .D(n10480), .Z(n4946) );
  AO4 U4423 ( .A(n10316), .B(n2785), .C(n2786), .D(n10480), .Z(n4947) );
  AO4 U4424 ( .A(n10316), .B(n2786), .C(n2787), .D(n10480), .Z(n4948) );
  AO4 U4425 ( .A(n10316), .B(n2787), .C(n2788), .D(n10480), .Z(n4949) );
  AO4 U4426 ( .A(n10316), .B(n2788), .C(n2789), .D(n10480), .Z(n4950) );
  AO4 U4427 ( .A(n10316), .B(n2789), .C(n2790), .D(n10480), .Z(n4951) );
  AO4 U4428 ( .A(n10316), .B(n2790), .C(n2791), .D(n10480), .Z(n4952) );
  AO4 U4429 ( .A(n10316), .B(n2791), .C(n2792), .D(n10480), .Z(n4953) );
  AO4 U4430 ( .A(n10316), .B(n2792), .C(n2793), .D(n10480), .Z(n4954) );
  AO4 U4431 ( .A(n10315), .B(n2793), .C(n2794), .D(n10480), .Z(n4955) );
  AO4 U4432 ( .A(n10315), .B(n2794), .C(n2795), .D(n10479), .Z(n4956) );
  AO4 U4433 ( .A(n10315), .B(n2795), .C(n2796), .D(n10479), .Z(n4957) );
  AO4 U4434 ( .A(n10315), .B(n2796), .C(n2797), .D(n10479), .Z(n4958) );
  AO4 U4435 ( .A(n10315), .B(n2797), .C(n2798), .D(n10479), .Z(n4959) );
  AO4 U4436 ( .A(n10315), .B(n2798), .C(n2799), .D(n10479), .Z(n4960) );
  AO4 U4437 ( .A(n10315), .B(n2799), .C(n2800), .D(n10479), .Z(n4961) );
  AO4 U4438 ( .A(n10315), .B(n2800), .C(n2801), .D(n10479), .Z(n4962) );
  AO4 U4439 ( .A(n10315), .B(n2801), .C(n2802), .D(n10479), .Z(n4963) );
  AO4 U4440 ( .A(n10315), .B(n2802), .C(n2803), .D(n10479), .Z(n4964) );
  AO4 U4441 ( .A(n10315), .B(n2803), .C(n2804), .D(n10479), .Z(n4965) );
  AO4 U4442 ( .A(n10315), .B(n2804), .C(n2805), .D(n10479), .Z(n4966) );
  AO4 U4443 ( .A(n10315), .B(n2805), .C(n2806), .D(n10479), .Z(n4967) );
  AO4 U4444 ( .A(n10315), .B(n2806), .C(n2807), .D(n10479), .Z(n4968) );
  AO4 U4445 ( .A(n10314), .B(n2807), .C(n2808), .D(n10479), .Z(n4969) );
  AO4 U4446 ( .A(n10314), .B(n2808), .C(n2809), .D(n10478), .Z(n4970) );
  AO4 U4447 ( .A(n10314), .B(n2809), .C(n2810), .D(n10478), .Z(n4971) );
  AO4 U4448 ( .A(n10314), .B(n2810), .C(n2811), .D(n10478), .Z(n4972) );
  AO4 U4449 ( .A(n10314), .B(n2811), .C(n2812), .D(n10478), .Z(n4973) );
  AO4 U4450 ( .A(n10314), .B(n2812), .C(n2813), .D(n10478), .Z(n4974) );
  AO4 U4451 ( .A(n10314), .B(n2813), .C(n2814), .D(n10478), .Z(n4975) );
  AO4 U4452 ( .A(n10314), .B(n2814), .C(n2815), .D(n10478), .Z(n4976) );
  AO4 U4453 ( .A(n10314), .B(n2815), .C(n2816), .D(n10478), .Z(n4977) );
  AO4 U4454 ( .A(n10314), .B(n2816), .C(n2817), .D(n10478), .Z(n4978) );
  AO4 U4455 ( .A(n10314), .B(n2817), .C(n2818), .D(n10478), .Z(n4979) );
  AO4 U4456 ( .A(n10314), .B(n2818), .C(n10478), .D(n1409), .Z(n4980) );
  AO4 U4457 ( .A(n10478), .B(n2754), .C(n10314), .D(n1409), .Z(n5857) );
  EN U4458 ( .A(n10252), .B(n10637), .Z(n2820) );
  EN U4459 ( .A(n10245), .B(n10637), .Z(n2821) );
  EN U4460 ( .A(n10242), .B(n10637), .Z(n2822) );
  EN U4461 ( .A(n10239), .B(n10637), .Z(n2823) );
  EN U4462 ( .A(n10236), .B(n10637), .Z(n2824) );
  EN U4463 ( .A(n10233), .B(n10637), .Z(n2825) );
  EN U4464 ( .A(n10230), .B(n10637), .Z(n2826) );
  EN U4465 ( .A(n10227), .B(n10637), .Z(n2827) );
  EN U4466 ( .A(n10224), .B(n10637), .Z(n2828) );
  EN U4467 ( .A(n10221), .B(n10636), .Z(n2829) );
  EN U4468 ( .A(n10218), .B(n10636), .Z(n2830) );
  EN U4469 ( .A(n10215), .B(n10636), .Z(n2831) );
  EN U4470 ( .A(n10212), .B(n10636), .Z(n2832) );
  EN U4471 ( .A(n10209), .B(n10636), .Z(n2833) );
  EN U4472 ( .A(n10206), .B(n10636), .Z(n2834) );
  EN U4473 ( .A(n10203), .B(n10636), .Z(n2835) );
  EN U4474 ( .A(n10200), .B(n10636), .Z(n2836) );
  EN U4475 ( .A(n10197), .B(n10636), .Z(n2837) );
  EN U4476 ( .A(n10194), .B(n10636), .Z(n2838) );
  EN U4477 ( .A(n10191), .B(n10636), .Z(n2839) );
  EN U4478 ( .A(n10188), .B(n10636), .Z(n2840) );
  EN U4479 ( .A(n10185), .B(n10636), .Z(n2841) );
  EN U4480 ( .A(n10182), .B(n10636), .Z(n2842) );
  EN U4481 ( .A(n10179), .B(n10635), .Z(n2843) );
  EN U4482 ( .A(n10176), .B(n10635), .Z(n2844) );
  EN U4483 ( .A(n10173), .B(n10635), .Z(n2845) );
  EN U4484 ( .A(n10170), .B(n10635), .Z(n2846) );
  EN U4485 ( .A(n10167), .B(n10635), .Z(n2847) );
  EN U4486 ( .A(n10164), .B(n10635), .Z(n2848) );
  EN U4487 ( .A(n10161), .B(n10635), .Z(n2849) );
  EN U4488 ( .A(n10158), .B(n10635), .Z(n2850) );
  EN U4489 ( .A(n10155), .B(n10635), .Z(n2851) );
  EN U4490 ( .A(n10152), .B(n10635), .Z(n2852) );
  EN U4491 ( .A(n10149), .B(n10635), .Z(n2853) );
  EN U4492 ( .A(n10146), .B(n10635), .Z(n2854) );
  EN U4493 ( .A(n10143), .B(n10635), .Z(n2855) );
  EN U4494 ( .A(n10140), .B(n10635), .Z(n2856) );
  EN U4495 ( .A(n10137), .B(n10634), .Z(n2857) );
  EN U4496 ( .A(n10134), .B(n10634), .Z(n2858) );
  EN U4497 ( .A(n10131), .B(n10634), .Z(n2859) );
  EN U4498 ( .A(n10128), .B(n10634), .Z(n2860) );
  EN U4499 ( .A(n10125), .B(n10634), .Z(n2861) );
  EN U4500 ( .A(n10122), .B(n10634), .Z(n2862) );
  EN U4501 ( .A(n10119), .B(n10634), .Z(n2863) );
  EN U4502 ( .A(n10116), .B(n10634), .Z(n2864) );
  EN U4503 ( .A(n10113), .B(n10634), .Z(n2865) );
  EN U4504 ( .A(n10110), .B(n10634), .Z(n2866) );
  EN U4505 ( .A(n10107), .B(n10634), .Z(n2867) );
  EN U4506 ( .A(n10104), .B(n10634), .Z(n2868) );
  EN U4507 ( .A(n10101), .B(n10634), .Z(n2869) );
  EN U4508 ( .A(n10098), .B(n10634), .Z(n2870) );
  EN U4509 ( .A(n10095), .B(n10633), .Z(n2871) );
  EN U4510 ( .A(n10092), .B(n10633), .Z(n2872) );
  EN U4511 ( .A(n10089), .B(n10633), .Z(n2873) );
  EN U4512 ( .A(n10086), .B(n10633), .Z(n2874) );
  EN U4513 ( .A(n10083), .B(n10633), .Z(n2875) );
  EN U4514 ( .A(n10080), .B(n10633), .Z(n2876) );
  EN U4515 ( .A(n10077), .B(n10633), .Z(n2877) );
  EN U4516 ( .A(n10074), .B(n10633), .Z(n2878) );
  EN U4517 ( .A(n10071), .B(n10633), .Z(n2879) );
  EN U4518 ( .A(n10068), .B(n10633), .Z(n2880) );
  EN U4519 ( .A(n10065), .B(n10633), .Z(n2881) );
  EN U4520 ( .A(n10062), .B(n10633), .Z(n2882) );
  EN U4521 ( .A(n10059), .B(n10633), .Z(n2883) );
  AO4 U4522 ( .A(n10313), .B(n2820), .C(n2821), .D(n10477), .Z(n4983) );
  AO4 U4523 ( .A(n10313), .B(n2821), .C(n2822), .D(n10477), .Z(n4984) );
  AO4 U4524 ( .A(n10313), .B(n2822), .C(n2823), .D(n10477), .Z(n4985) );
  AO4 U4525 ( .A(n10313), .B(n2823), .C(n2824), .D(n10477), .Z(n4986) );
  AO4 U4526 ( .A(n10313), .B(n2824), .C(n2825), .D(n10477), .Z(n4987) );
  AO4 U4527 ( .A(n10313), .B(n2825), .C(n2826), .D(n10477), .Z(n4988) );
  AO4 U4528 ( .A(n10313), .B(n2826), .C(n2827), .D(n10477), .Z(n4989) );
  AO4 U4529 ( .A(n10313), .B(n2827), .C(n2828), .D(n10477), .Z(n4990) );
  AO4 U4530 ( .A(n10313), .B(n2828), .C(n2829), .D(n10477), .Z(n4991) );
  AO4 U4531 ( .A(n10313), .B(n2829), .C(n2830), .D(n10477), .Z(n4992) );
  AO4 U4532 ( .A(n10312), .B(n2830), .C(n2831), .D(n10477), .Z(n4993) );
  AO4 U4533 ( .A(n10312), .B(n2831), .C(n2832), .D(n10476), .Z(n4994) );
  AO4 U4534 ( .A(n10312), .B(n2832), .C(n2833), .D(n10476), .Z(n4995) );
  AO4 U4535 ( .A(n10312), .B(n2833), .C(n2834), .D(n10476), .Z(n4996) );
  AO4 U4536 ( .A(n10312), .B(n2834), .C(n2835), .D(n10476), .Z(n4997) );
  AO4 U4537 ( .A(n10312), .B(n2835), .C(n2836), .D(n10476), .Z(n4998) );
  AO4 U4538 ( .A(n10312), .B(n2836), .C(n2837), .D(n10476), .Z(n4999) );
  AO4 U4539 ( .A(n10312), .B(n2837), .C(n2838), .D(n10476), .Z(n5000) );
  AO4 U4540 ( .A(n10312), .B(n2838), .C(n2839), .D(n10476), .Z(n5001) );
  AO4 U4541 ( .A(n10312), .B(n2839), .C(n2840), .D(n10476), .Z(n5002) );
  AO4 U4542 ( .A(n10312), .B(n2840), .C(n2841), .D(n10476), .Z(n5003) );
  AO4 U4543 ( .A(n10312), .B(n2841), .C(n2842), .D(n10476), .Z(n5004) );
  AO4 U4544 ( .A(n10312), .B(n2842), .C(n2843), .D(n10476), .Z(n5005) );
  AO4 U4545 ( .A(n10312), .B(n2843), .C(n2844), .D(n10476), .Z(n5006) );
  AO4 U4546 ( .A(n10311), .B(n2844), .C(n2845), .D(n10476), .Z(n5007) );
  AO4 U4547 ( .A(n10311), .B(n2845), .C(n2846), .D(n10475), .Z(n5008) );
  AO4 U4548 ( .A(n10311), .B(n2846), .C(n2847), .D(n10475), .Z(n5009) );
  AO4 U4549 ( .A(n10311), .B(n2847), .C(n2848), .D(n10475), .Z(n5010) );
  AO4 U4550 ( .A(n10311), .B(n2848), .C(n2849), .D(n10475), .Z(n5011) );
  AO4 U4551 ( .A(n10311), .B(n2849), .C(n2850), .D(n10475), .Z(n5012) );
  AO4 U4552 ( .A(n10311), .B(n2850), .C(n2851), .D(n10475), .Z(n5013) );
  AO4 U4553 ( .A(n10311), .B(n2851), .C(n2852), .D(n10475), .Z(n5014) );
  AO4 U4554 ( .A(n10311), .B(n2852), .C(n2853), .D(n10475), .Z(n5015) );
  AO4 U4555 ( .A(n10311), .B(n2853), .C(n2854), .D(n10475), .Z(n5016) );
  AO4 U4556 ( .A(n10311), .B(n2854), .C(n2855), .D(n10475), .Z(n5017) );
  AO4 U4557 ( .A(n10311), .B(n2855), .C(n2856), .D(n10475), .Z(n5018) );
  AO4 U4558 ( .A(n10311), .B(n2856), .C(n2857), .D(n10475), .Z(n5019) );
  AO4 U4559 ( .A(n10311), .B(n2857), .C(n2858), .D(n10475), .Z(n5020) );
  AO4 U4560 ( .A(n10310), .B(n2858), .C(n2859), .D(n10475), .Z(n5021) );
  AO4 U4561 ( .A(n10310), .B(n2859), .C(n2860), .D(n10474), .Z(n5022) );
  AO4 U4562 ( .A(n10310), .B(n2860), .C(n2861), .D(n10474), .Z(n5023) );
  AO4 U4563 ( .A(n10310), .B(n2861), .C(n2862), .D(n10474), .Z(n5024) );
  AO4 U4564 ( .A(n10310), .B(n2862), .C(n2863), .D(n10474), .Z(n5025) );
  AO4 U4565 ( .A(n10310), .B(n2863), .C(n2864), .D(n10474), .Z(n5026) );
  AO4 U4566 ( .A(n10310), .B(n2864), .C(n2865), .D(n10474), .Z(n5027) );
  AO4 U4567 ( .A(n10310), .B(n2865), .C(n2866), .D(n10474), .Z(n5028) );
  AO4 U4568 ( .A(n10310), .B(n2866), .C(n2867), .D(n10474), .Z(n5029) );
  AO4 U4569 ( .A(n10310), .B(n2867), .C(n2868), .D(n10474), .Z(n5030) );
  AO4 U4570 ( .A(n10310), .B(n2868), .C(n2869), .D(n10474), .Z(n5031) );
  AO4 U4571 ( .A(n10310), .B(n2869), .C(n2870), .D(n10474), .Z(n5032) );
  AO4 U4572 ( .A(n10310), .B(n2870), .C(n2871), .D(n10474), .Z(n5033) );
  AO4 U4573 ( .A(n10310), .B(n2871), .C(n2872), .D(n10474), .Z(n5034) );
  AO4 U4574 ( .A(n10309), .B(n2872), .C(n2873), .D(n10474), .Z(n5035) );
  AO4 U4575 ( .A(n10309), .B(n2873), .C(n2874), .D(n10473), .Z(n5036) );
  AO4 U4576 ( .A(n10309), .B(n2874), .C(n2875), .D(n10473), .Z(n5037) );
  AO4 U4577 ( .A(n10309), .B(n2875), .C(n2876), .D(n10473), .Z(n5038) );
  AO4 U4578 ( .A(n10309), .B(n2876), .C(n2877), .D(n10473), .Z(n5039) );
  AO4 U4579 ( .A(n10309), .B(n2877), .C(n2878), .D(n10473), .Z(n5040) );
  AO4 U4580 ( .A(n10309), .B(n2878), .C(n2879), .D(n10473), .Z(n5041) );
  AO4 U4581 ( .A(n10309), .B(n2879), .C(n2880), .D(n10473), .Z(n5042) );
  AO4 U4582 ( .A(n10309), .B(n2880), .C(n2881), .D(n10473), .Z(n5043) );
  AO4 U4583 ( .A(n10309), .B(n2881), .C(n2882), .D(n10473), .Z(n5044) );
  AO4 U4584 ( .A(n10309), .B(n2882), .C(n2883), .D(n10473), .Z(n5045) );
  AO4 U4585 ( .A(n10309), .B(n2883), .C(n10473), .D(n1410), .Z(n5046) );
  AO4 U4586 ( .A(n10473), .B(n2819), .C(n10309), .D(n1410), .Z(n5858) );
  EN U4587 ( .A(n10252), .B(n10632), .Z(n2885) );
  EN U4588 ( .A(n10245), .B(n10632), .Z(n2886) );
  EN U4589 ( .A(n10242), .B(n10632), .Z(n2887) );
  EN U4590 ( .A(n10239), .B(n10632), .Z(n2888) );
  EN U4591 ( .A(n10236), .B(n10632), .Z(n2889) );
  EN U4592 ( .A(n10233), .B(n10632), .Z(n2890) );
  EN U4593 ( .A(n10230), .B(n10632), .Z(n2891) );
  EN U4594 ( .A(n10227), .B(n10632), .Z(n2892) );
  EN U4595 ( .A(n10224), .B(n10632), .Z(n2893) );
  EN U4596 ( .A(n10221), .B(n10631), .Z(n2894) );
  EN U4597 ( .A(n10218), .B(n10631), .Z(n2895) );
  EN U4598 ( .A(n10215), .B(n10631), .Z(n2896) );
  EN U4599 ( .A(n10212), .B(n10631), .Z(n2897) );
  EN U4600 ( .A(n10209), .B(n10631), .Z(n2898) );
  EN U4601 ( .A(n10206), .B(n10631), .Z(n2899) );
  EN U4602 ( .A(n10203), .B(n10631), .Z(n2900) );
  EN U4603 ( .A(n10200), .B(n10631), .Z(n2901) );
  EN U4604 ( .A(n10197), .B(n10631), .Z(n2902) );
  EN U4605 ( .A(n10194), .B(n10631), .Z(n2903) );
  EN U4606 ( .A(n10191), .B(n10631), .Z(n2904) );
  EN U4607 ( .A(n10188), .B(n10631), .Z(n2905) );
  EN U4608 ( .A(n10185), .B(n10631), .Z(n2906) );
  EN U4609 ( .A(n10182), .B(n10631), .Z(n2907) );
  EN U4610 ( .A(n10179), .B(n10630), .Z(n2908) );
  EN U4611 ( .A(n10176), .B(n10630), .Z(n2909) );
  EN U4612 ( .A(n10173), .B(n10630), .Z(n2910) );
  EN U4613 ( .A(n10170), .B(n10630), .Z(n2911) );
  EN U4614 ( .A(n10167), .B(n10630), .Z(n2912) );
  EN U4615 ( .A(n10164), .B(n10630), .Z(n2913) );
  EN U4616 ( .A(n10161), .B(n10630), .Z(n2914) );
  EN U4617 ( .A(n10158), .B(n10630), .Z(n2915) );
  EN U4618 ( .A(n10155), .B(n10630), .Z(n2916) );
  EN U4619 ( .A(n10152), .B(n10630), .Z(n2917) );
  EN U4620 ( .A(n10149), .B(n10630), .Z(n2918) );
  EN U4621 ( .A(n10146), .B(n10630), .Z(n2919) );
  EN U4622 ( .A(n10143), .B(n10630), .Z(n2920) );
  EN U4623 ( .A(n10140), .B(n10630), .Z(n2921) );
  EN U4624 ( .A(n10137), .B(n10629), .Z(n2922) );
  EN U4625 ( .A(n10134), .B(n10629), .Z(n2923) );
  EN U4626 ( .A(n10131), .B(n10629), .Z(n2924) );
  EN U4627 ( .A(n10128), .B(n10629), .Z(n2925) );
  EN U4628 ( .A(n10125), .B(n10629), .Z(n2926) );
  EN U4629 ( .A(n10122), .B(n10629), .Z(n2927) );
  EN U4630 ( .A(n10119), .B(n10629), .Z(n2928) );
  EN U4631 ( .A(n10116), .B(n10629), .Z(n2929) );
  EN U4632 ( .A(n10113), .B(n10629), .Z(n2930) );
  EN U4633 ( .A(n10110), .B(n10629), .Z(n2931) );
  EN U4634 ( .A(n10107), .B(n10629), .Z(n2932) );
  EN U4635 ( .A(n10104), .B(n10629), .Z(n2933) );
  EN U4636 ( .A(n10101), .B(n10629), .Z(n2934) );
  EN U4637 ( .A(n10098), .B(n10629), .Z(n2935) );
  EN U4638 ( .A(n10095), .B(n10628), .Z(n2936) );
  EN U4639 ( .A(n10092), .B(n10628), .Z(n2937) );
  EN U4640 ( .A(n10089), .B(n10628), .Z(n2938) );
  EN U4641 ( .A(n10086), .B(n10628), .Z(n2939) );
  EN U4642 ( .A(n10083), .B(n10628), .Z(n2940) );
  EN U4643 ( .A(n10080), .B(n10628), .Z(n2941) );
  EN U4644 ( .A(n10077), .B(n10628), .Z(n2942) );
  EN U4645 ( .A(n10074), .B(n10628), .Z(n2943) );
  EN U4646 ( .A(n10071), .B(n10628), .Z(n2944) );
  EN U4647 ( .A(n10068), .B(n10628), .Z(n2945) );
  EN U4648 ( .A(n10065), .B(n10628), .Z(n2946) );
  EN U4649 ( .A(n10062), .B(n10628), .Z(n2947) );
  EN U4650 ( .A(n10059), .B(n10628), .Z(n2948) );
  AO4 U4651 ( .A(n10308), .B(n2885), .C(n2886), .D(n10472), .Z(n5049) );
  AO4 U4652 ( .A(n10308), .B(n2886), .C(n2887), .D(n10472), .Z(n5050) );
  AO4 U4653 ( .A(n10308), .B(n2887), .C(n2888), .D(n10472), .Z(n5051) );
  AO4 U4654 ( .A(n10308), .B(n2888), .C(n2889), .D(n10472), .Z(n5052) );
  AO4 U4655 ( .A(n10308), .B(n2889), .C(n2890), .D(n10472), .Z(n5053) );
  AO4 U4656 ( .A(n10308), .B(n2890), .C(n2891), .D(n10472), .Z(n5054) );
  AO4 U4657 ( .A(n10308), .B(n2891), .C(n2892), .D(n10472), .Z(n5055) );
  AO4 U4658 ( .A(n10308), .B(n2892), .C(n2893), .D(n10472), .Z(n5056) );
  AO4 U4659 ( .A(n10308), .B(n2893), .C(n2894), .D(n10472), .Z(n5057) );
  AO4 U4660 ( .A(n10308), .B(n2894), .C(n2895), .D(n10472), .Z(n5058) );
  AO4 U4661 ( .A(n10307), .B(n2895), .C(n2896), .D(n10472), .Z(n5059) );
  AO4 U4662 ( .A(n10307), .B(n2896), .C(n2897), .D(n10471), .Z(n5060) );
  AO4 U4663 ( .A(n10307), .B(n2897), .C(n2898), .D(n10471), .Z(n5061) );
  AO4 U4664 ( .A(n10307), .B(n2898), .C(n2899), .D(n10471), .Z(n5062) );
  AO4 U4665 ( .A(n10307), .B(n2899), .C(n2900), .D(n10471), .Z(n5063) );
  AO4 U4666 ( .A(n10307), .B(n2900), .C(n2901), .D(n10471), .Z(n5064) );
  AO4 U4667 ( .A(n10307), .B(n2901), .C(n2902), .D(n10471), .Z(n5065) );
  AO4 U4668 ( .A(n10307), .B(n2902), .C(n2903), .D(n10471), .Z(n5066) );
  AO4 U4669 ( .A(n10307), .B(n2903), .C(n2904), .D(n10471), .Z(n5067) );
  AO4 U4670 ( .A(n10307), .B(n2904), .C(n2905), .D(n10471), .Z(n5068) );
  AO4 U4671 ( .A(n10307), .B(n2905), .C(n2906), .D(n10471), .Z(n5069) );
  AO4 U4672 ( .A(n10307), .B(n2906), .C(n2907), .D(n10471), .Z(n5070) );
  AO4 U4673 ( .A(n10307), .B(n2907), .C(n2908), .D(n10471), .Z(n5071) );
  AO4 U4674 ( .A(n10307), .B(n2908), .C(n2909), .D(n10471), .Z(n5072) );
  AO4 U4675 ( .A(n10306), .B(n2909), .C(n2910), .D(n10471), .Z(n5073) );
  AO4 U4676 ( .A(n10306), .B(n2910), .C(n2911), .D(n10470), .Z(n5074) );
  AO4 U4677 ( .A(n10306), .B(n2911), .C(n2912), .D(n10470), .Z(n5075) );
  AO4 U4678 ( .A(n10306), .B(n2912), .C(n2913), .D(n10470), .Z(n5076) );
  AO4 U4679 ( .A(n10306), .B(n2913), .C(n2914), .D(n10470), .Z(n5077) );
  AO4 U4680 ( .A(n10306), .B(n2914), .C(n2915), .D(n10470), .Z(n5078) );
  AO4 U4681 ( .A(n10306), .B(n2915), .C(n2916), .D(n10470), .Z(n5079) );
  AO4 U4682 ( .A(n10306), .B(n2916), .C(n2917), .D(n10470), .Z(n5080) );
  AO4 U4683 ( .A(n10306), .B(n2917), .C(n2918), .D(n10470), .Z(n5081) );
  AO4 U4684 ( .A(n10306), .B(n2918), .C(n2919), .D(n10470), .Z(n5082) );
  AO4 U4685 ( .A(n10306), .B(n2919), .C(n2920), .D(n10470), .Z(n5083) );
  AO4 U4686 ( .A(n10306), .B(n2920), .C(n2921), .D(n10470), .Z(n5084) );
  AO4 U4687 ( .A(n10306), .B(n2921), .C(n2922), .D(n10470), .Z(n5085) );
  AO4 U4688 ( .A(n10306), .B(n2922), .C(n2923), .D(n10470), .Z(n5086) );
  AO4 U4689 ( .A(n10305), .B(n2923), .C(n2924), .D(n10470), .Z(n5087) );
  AO4 U4690 ( .A(n10305), .B(n2924), .C(n2925), .D(n10469), .Z(n5088) );
  AO4 U4691 ( .A(n10305), .B(n2925), .C(n2926), .D(n10469), .Z(n5089) );
  AO4 U4692 ( .A(n10305), .B(n2926), .C(n2927), .D(n10469), .Z(n5090) );
  AO4 U4693 ( .A(n10305), .B(n2927), .C(n2928), .D(n10469), .Z(n5091) );
  AO4 U4694 ( .A(n10305), .B(n2928), .C(n2929), .D(n10469), .Z(n5092) );
  AO4 U4695 ( .A(n10305), .B(n2929), .C(n2930), .D(n10469), .Z(n5093) );
  AO4 U4696 ( .A(n10305), .B(n2930), .C(n2931), .D(n10469), .Z(n5094) );
  AO4 U4697 ( .A(n10305), .B(n2931), .C(n2932), .D(n10469), .Z(n5095) );
  AO4 U4698 ( .A(n10305), .B(n2932), .C(n2933), .D(n10469), .Z(n5096) );
  AO4 U4699 ( .A(n10305), .B(n2933), .C(n2934), .D(n10469), .Z(n5097) );
  AO4 U4700 ( .A(n10305), .B(n2934), .C(n2935), .D(n10469), .Z(n5098) );
  AO4 U4701 ( .A(n10305), .B(n2935), .C(n2936), .D(n10469), .Z(n5099) );
  AO4 U4702 ( .A(n10305), .B(n2936), .C(n2937), .D(n10469), .Z(n5100) );
  AO4 U4703 ( .A(n10304), .B(n2937), .C(n2938), .D(n10469), .Z(n5101) );
  AO4 U4704 ( .A(n10304), .B(n2938), .C(n2939), .D(n10468), .Z(n5102) );
  AO4 U4705 ( .A(n10304), .B(n2939), .C(n2940), .D(n10468), .Z(n5103) );
  AO4 U4706 ( .A(n10304), .B(n2940), .C(n2941), .D(n10468), .Z(n5104) );
  AO4 U4707 ( .A(n10304), .B(n2941), .C(n2942), .D(n10468), .Z(n5105) );
  AO4 U4708 ( .A(n10304), .B(n2942), .C(n2943), .D(n10468), .Z(n5106) );
  AO4 U4709 ( .A(n10304), .B(n2943), .C(n2944), .D(n10468), .Z(n5107) );
  AO4 U4710 ( .A(n10304), .B(n2944), .C(n2945), .D(n10468), .Z(n5108) );
  AO4 U4711 ( .A(n10304), .B(n2945), .C(n2946), .D(n10468), .Z(n5109) );
  AO4 U4712 ( .A(n10304), .B(n2946), .C(n2947), .D(n10468), .Z(n5110) );
  AO4 U4713 ( .A(n10304), .B(n2947), .C(n2948), .D(n10468), .Z(n5111) );
  AO4 U4714 ( .A(n10304), .B(n2948), .C(n10468), .D(n1411), .Z(n5112) );
  AO4 U4715 ( .A(n10468), .B(n2884), .C(n10304), .D(n1411), .Z(n5859) );
  EN U4716 ( .A(n10252), .B(n10627), .Z(n2950) );
  EN U4717 ( .A(n10244), .B(n10627), .Z(n2951) );
  EN U4718 ( .A(n10241), .B(n10627), .Z(n2952) );
  EN U4719 ( .A(n10238), .B(n10627), .Z(n2953) );
  EN U4720 ( .A(n10235), .B(n10627), .Z(n2954) );
  EN U4721 ( .A(n10232), .B(n10627), .Z(n2955) );
  EN U4722 ( .A(n10229), .B(n10627), .Z(n2956) );
  EN U4723 ( .A(n10226), .B(n10627), .Z(n2957) );
  EN U4724 ( .A(n10223), .B(n10627), .Z(n2958) );
  EN U4725 ( .A(n10220), .B(n10626), .Z(n2959) );
  EN U4726 ( .A(n10217), .B(n10626), .Z(n2960) );
  EN U4727 ( .A(n10214), .B(n10626), .Z(n2961) );
  EN U4728 ( .A(n10211), .B(n10626), .Z(n2962) );
  EN U4729 ( .A(n10208), .B(n10626), .Z(n2963) );
  EN U4730 ( .A(n10205), .B(n10626), .Z(n2964) );
  EN U4731 ( .A(n10202), .B(n10626), .Z(n2965) );
  EN U4732 ( .A(n10199), .B(n10626), .Z(n2966) );
  EN U4733 ( .A(n10196), .B(n10626), .Z(n2967) );
  EN U4734 ( .A(n10193), .B(n10626), .Z(n2968) );
  EN U4735 ( .A(n10190), .B(n10626), .Z(n2969) );
  EN U4736 ( .A(n10187), .B(n10626), .Z(n2970) );
  EN U4737 ( .A(n10184), .B(n10626), .Z(n2971) );
  EN U4738 ( .A(n10181), .B(n10626), .Z(n2972) );
  EN U4739 ( .A(n10178), .B(n10625), .Z(n2973) );
  EN U4740 ( .A(n10175), .B(n10625), .Z(n2974) );
  EN U4741 ( .A(n10172), .B(n10625), .Z(n2975) );
  EN U4742 ( .A(n10169), .B(n10625), .Z(n2976) );
  EN U4743 ( .A(n10166), .B(n10625), .Z(n2977) );
  EN U4744 ( .A(n10163), .B(n10625), .Z(n2978) );
  EN U4745 ( .A(n10160), .B(n10625), .Z(n2979) );
  EN U4746 ( .A(n10157), .B(n10625), .Z(n2980) );
  EN U4747 ( .A(n10154), .B(n10625), .Z(n2981) );
  EN U4748 ( .A(n10151), .B(n10625), .Z(n2982) );
  EN U4749 ( .A(n10148), .B(n10625), .Z(n2983) );
  EN U4750 ( .A(n10145), .B(n10625), .Z(n2984) );
  EN U4751 ( .A(n10142), .B(n10625), .Z(n2985) );
  EN U4752 ( .A(n10139), .B(n10625), .Z(n2986) );
  EN U4753 ( .A(n10136), .B(n10624), .Z(n2987) );
  EN U4754 ( .A(n10133), .B(n10624), .Z(n2988) );
  EN U4755 ( .A(n10130), .B(n10624), .Z(n2989) );
  EN U4756 ( .A(n10127), .B(n10624), .Z(n2990) );
  EN U4757 ( .A(n10124), .B(n10624), .Z(n2991) );
  EN U4758 ( .A(n10121), .B(n10624), .Z(n2992) );
  EN U4759 ( .A(n10118), .B(n10624), .Z(n2993) );
  EN U4760 ( .A(n10115), .B(n10624), .Z(n2994) );
  EN U4761 ( .A(n10112), .B(n10624), .Z(n2995) );
  EN U4762 ( .A(n10109), .B(n10624), .Z(n2996) );
  EN U4763 ( .A(n10106), .B(n10624), .Z(n2997) );
  EN U4764 ( .A(n10103), .B(n10624), .Z(n2998) );
  EN U4765 ( .A(n10100), .B(n10624), .Z(n2999) );
  EN U4766 ( .A(n10097), .B(n10624), .Z(n3000) );
  EN U4767 ( .A(n10094), .B(n10623), .Z(n3001) );
  EN U4768 ( .A(n10091), .B(n10623), .Z(n3002) );
  EN U4769 ( .A(n10088), .B(n10623), .Z(n3003) );
  EN U4770 ( .A(n10085), .B(n10623), .Z(n3004) );
  EN U4771 ( .A(n10082), .B(n10623), .Z(n3005) );
  EN U4772 ( .A(n10079), .B(n10623), .Z(n3006) );
  EN U4773 ( .A(n10076), .B(n10623), .Z(n3007) );
  EN U4774 ( .A(n10073), .B(n10623), .Z(n3008) );
  EN U4775 ( .A(n10070), .B(n10623), .Z(n3009) );
  EN U4776 ( .A(n10067), .B(n10623), .Z(n3010) );
  EN U4777 ( .A(n10064), .B(n10623), .Z(n3011) );
  EN U4778 ( .A(n10061), .B(n10623), .Z(n3012) );
  EN U4779 ( .A(n10058), .B(n10623), .Z(n3013) );
  AO4 U4780 ( .A(n10303), .B(n2950), .C(n2951), .D(n10467), .Z(n5115) );
  AO4 U4781 ( .A(n10303), .B(n2951), .C(n2952), .D(n10467), .Z(n5116) );
  AO4 U4782 ( .A(n10303), .B(n2952), .C(n2953), .D(n10467), .Z(n5117) );
  AO4 U4783 ( .A(n10303), .B(n2953), .C(n2954), .D(n10467), .Z(n5118) );
  AO4 U4784 ( .A(n10303), .B(n2954), .C(n2955), .D(n10467), .Z(n5119) );
  AO4 U4785 ( .A(n10303), .B(n2955), .C(n2956), .D(n10467), .Z(n5120) );
  AO4 U4786 ( .A(n10303), .B(n2956), .C(n2957), .D(n10467), .Z(n5121) );
  AO4 U4787 ( .A(n10303), .B(n2957), .C(n2958), .D(n10467), .Z(n5122) );
  AO4 U4788 ( .A(n10303), .B(n2958), .C(n2959), .D(n10467), .Z(n5123) );
  AO4 U4789 ( .A(n10303), .B(n2959), .C(n2960), .D(n10467), .Z(n5124) );
  AO4 U4790 ( .A(n10302), .B(n2960), .C(n2961), .D(n10467), .Z(n5125) );
  AO4 U4791 ( .A(n10302), .B(n2961), .C(n2962), .D(n10466), .Z(n5126) );
  AO4 U4792 ( .A(n10302), .B(n2962), .C(n2963), .D(n10466), .Z(n5127) );
  AO4 U4793 ( .A(n10302), .B(n2963), .C(n2964), .D(n10466), .Z(n5128) );
  AO4 U4794 ( .A(n10302), .B(n2964), .C(n2965), .D(n10466), .Z(n5129) );
  AO4 U4795 ( .A(n10302), .B(n2965), .C(n2966), .D(n10466), .Z(n5130) );
  AO4 U4796 ( .A(n10302), .B(n2966), .C(n2967), .D(n10466), .Z(n5131) );
  AO4 U4797 ( .A(n10302), .B(n2967), .C(n2968), .D(n10466), .Z(n5132) );
  AO4 U4798 ( .A(n10302), .B(n2968), .C(n2969), .D(n10466), .Z(n5133) );
  AO4 U4799 ( .A(n10302), .B(n2969), .C(n2970), .D(n10466), .Z(n5134) );
  AO4 U4800 ( .A(n10302), .B(n2970), .C(n2971), .D(n10466), .Z(n5135) );
  AO4 U4801 ( .A(n10302), .B(n2971), .C(n2972), .D(n10466), .Z(n5136) );
  AO4 U4802 ( .A(n10302), .B(n2972), .C(n2973), .D(n10466), .Z(n5137) );
  AO4 U4803 ( .A(n10302), .B(n2973), .C(n2974), .D(n10466), .Z(n5138) );
  AO4 U4804 ( .A(n10301), .B(n2974), .C(n2975), .D(n10466), .Z(n5139) );
  AO4 U4805 ( .A(n10301), .B(n2975), .C(n2976), .D(n10465), .Z(n5140) );
  AO4 U4806 ( .A(n10301), .B(n2976), .C(n2977), .D(n10465), .Z(n5141) );
  AO4 U4807 ( .A(n10301), .B(n2977), .C(n2978), .D(n10465), .Z(n5142) );
  AO4 U4808 ( .A(n10301), .B(n2978), .C(n2979), .D(n10465), .Z(n5143) );
  AO4 U4809 ( .A(n10301), .B(n2979), .C(n2980), .D(n10465), .Z(n5144) );
  AO4 U4810 ( .A(n10301), .B(n2980), .C(n2981), .D(n10465), .Z(n5145) );
  AO4 U4811 ( .A(n10301), .B(n2981), .C(n2982), .D(n10465), .Z(n5146) );
  AO4 U4812 ( .A(n10301), .B(n2982), .C(n2983), .D(n10465), .Z(n5147) );
  AO4 U4813 ( .A(n10301), .B(n2983), .C(n2984), .D(n10465), .Z(n5148) );
  AO4 U4814 ( .A(n10301), .B(n2984), .C(n2985), .D(n10465), .Z(n5149) );
  AO4 U4815 ( .A(n10301), .B(n2985), .C(n2986), .D(n10465), .Z(n5150) );
  AO4 U4816 ( .A(n10301), .B(n2986), .C(n2987), .D(n10465), .Z(n5151) );
  AO4 U4817 ( .A(n10301), .B(n2987), .C(n2988), .D(n10465), .Z(n5152) );
  AO4 U4818 ( .A(n10300), .B(n2988), .C(n2989), .D(n10465), .Z(n5153) );
  AO4 U4819 ( .A(n10300), .B(n2989), .C(n2990), .D(n10464), .Z(n5154) );
  AO4 U4820 ( .A(n10300), .B(n2990), .C(n2991), .D(n10464), .Z(n5155) );
  AO4 U4821 ( .A(n10300), .B(n2991), .C(n2992), .D(n10464), .Z(n5156) );
  AO4 U4822 ( .A(n10300), .B(n2992), .C(n2993), .D(n10464), .Z(n5157) );
  AO4 U4823 ( .A(n10300), .B(n2993), .C(n2994), .D(n10464), .Z(n5158) );
  AO4 U4824 ( .A(n10300), .B(n2994), .C(n2995), .D(n10464), .Z(n5159) );
  AO4 U4825 ( .A(n10300), .B(n2995), .C(n2996), .D(n10464), .Z(n5160) );
  AO4 U4826 ( .A(n10300), .B(n2996), .C(n2997), .D(n10464), .Z(n5161) );
  AO4 U4827 ( .A(n10300), .B(n2997), .C(n2998), .D(n10464), .Z(n5162) );
  AO4 U4828 ( .A(n10300), .B(n2998), .C(n2999), .D(n10464), .Z(n5163) );
  AO4 U4829 ( .A(n10300), .B(n2999), .C(n3000), .D(n10464), .Z(n5164) );
  AO4 U4830 ( .A(n10300), .B(n3000), .C(n3001), .D(n10464), .Z(n5165) );
  AO4 U4831 ( .A(n10300), .B(n3001), .C(n3002), .D(n10464), .Z(n5166) );
  AO4 U4832 ( .A(n10299), .B(n3002), .C(n3003), .D(n10464), .Z(n5167) );
  AO4 U4833 ( .A(n10299), .B(n3003), .C(n3004), .D(n10463), .Z(n5168) );
  AO4 U4834 ( .A(n10299), .B(n3004), .C(n3005), .D(n10463), .Z(n5169) );
  AO4 U4835 ( .A(n10299), .B(n3005), .C(n3006), .D(n10463), .Z(n5170) );
  AO4 U4836 ( .A(n10299), .B(n3006), .C(n3007), .D(n10463), .Z(n5171) );
  AO4 U4837 ( .A(n10299), .B(n3007), .C(n3008), .D(n10463), .Z(n5172) );
  AO4 U4838 ( .A(n10299), .B(n3008), .C(n3009), .D(n10463), .Z(n5173) );
  AO4 U4839 ( .A(n10299), .B(n3009), .C(n3010), .D(n10463), .Z(n5174) );
  AO4 U4840 ( .A(n10299), .B(n3010), .C(n3011), .D(n10463), .Z(n5175) );
  AO4 U4841 ( .A(n10299), .B(n3011), .C(n3012), .D(n10463), .Z(n5176) );
  AO4 U4842 ( .A(n10299), .B(n3012), .C(n3013), .D(n10463), .Z(n5177) );
  AO4 U4843 ( .A(n10299), .B(n3013), .C(n10463), .D(n1412), .Z(n5178) );
  AO4 U4844 ( .A(n10463), .B(n2949), .C(n10299), .D(n1412), .Z(n5860) );
  EN U4845 ( .A(n10252), .B(n10622), .Z(n3015) );
  EN U4846 ( .A(n10244), .B(n10622), .Z(n3016) );
  EN U4847 ( .A(n10241), .B(n10622), .Z(n3017) );
  EN U4848 ( .A(n10238), .B(n10622), .Z(n3018) );
  EN U4849 ( .A(n10235), .B(n10622), .Z(n3019) );
  EN U4850 ( .A(n10232), .B(n10622), .Z(n3020) );
  EN U4851 ( .A(n10229), .B(n10622), .Z(n3021) );
  EN U4852 ( .A(n10226), .B(n10622), .Z(n3022) );
  EN U4853 ( .A(n10223), .B(n10622), .Z(n3023) );
  EN U4854 ( .A(n10220), .B(n10621), .Z(n3024) );
  EN U4855 ( .A(n10217), .B(n10621), .Z(n3025) );
  EN U4856 ( .A(n10214), .B(n10621), .Z(n3026) );
  EN U4857 ( .A(n10211), .B(n10621), .Z(n3027) );
  EN U4858 ( .A(n10208), .B(n10621), .Z(n3028) );
  EN U4859 ( .A(n10205), .B(n10621), .Z(n3029) );
  EN U4860 ( .A(n10202), .B(n10621), .Z(n3030) );
  EN U4861 ( .A(n10199), .B(n10621), .Z(n3031) );
  EN U4862 ( .A(n10196), .B(n10621), .Z(n3032) );
  EN U4863 ( .A(n10193), .B(n10621), .Z(n3033) );
  EN U4864 ( .A(n10190), .B(n10621), .Z(n3034) );
  EN U4865 ( .A(n10187), .B(n10621), .Z(n3035) );
  EN U4866 ( .A(n10184), .B(n10621), .Z(n3036) );
  EN U4867 ( .A(n10181), .B(n10621), .Z(n3037) );
  EN U4868 ( .A(n10178), .B(n10620), .Z(n3038) );
  EN U4869 ( .A(n10175), .B(n10620), .Z(n3039) );
  EN U4870 ( .A(n10172), .B(n10620), .Z(n3040) );
  EN U4871 ( .A(n10169), .B(n10620), .Z(n3041) );
  EN U4872 ( .A(n10166), .B(n10620), .Z(n3042) );
  EN U4873 ( .A(n10163), .B(n10620), .Z(n3043) );
  EN U4874 ( .A(n10160), .B(n10620), .Z(n3044) );
  EN U4875 ( .A(n10157), .B(n10620), .Z(n3045) );
  EN U4876 ( .A(n10154), .B(n10620), .Z(n3046) );
  EN U4877 ( .A(n10151), .B(n10620), .Z(n3047) );
  EN U4878 ( .A(n10148), .B(n10620), .Z(n3048) );
  EN U4879 ( .A(n10145), .B(n10620), .Z(n3049) );
  EN U4880 ( .A(n10142), .B(n10620), .Z(n3050) );
  EN U4881 ( .A(n10139), .B(n10620), .Z(n3051) );
  EN U4882 ( .A(n10136), .B(n10619), .Z(n3052) );
  EN U4883 ( .A(n10133), .B(n10619), .Z(n3053) );
  EN U4884 ( .A(n10130), .B(n10619), .Z(n3054) );
  EN U4885 ( .A(n10127), .B(n10619), .Z(n3055) );
  EN U4886 ( .A(n10124), .B(n10619), .Z(n3056) );
  EN U4887 ( .A(n10121), .B(n10619), .Z(n3057) );
  EN U4888 ( .A(n10118), .B(n10619), .Z(n3058) );
  EN U4889 ( .A(n10115), .B(n10619), .Z(n3059) );
  EN U4890 ( .A(n10112), .B(n10619), .Z(n3060) );
  EN U4891 ( .A(n10109), .B(n10619), .Z(n3061) );
  EN U4892 ( .A(n10106), .B(n10619), .Z(n3062) );
  EN U4893 ( .A(n10103), .B(n10619), .Z(n3063) );
  EN U4894 ( .A(n10100), .B(n10619), .Z(n3064) );
  EN U4895 ( .A(n10097), .B(n10619), .Z(n3065) );
  EN U4896 ( .A(n10094), .B(n10618), .Z(n3066) );
  EN U4897 ( .A(n10091), .B(n10618), .Z(n3067) );
  EN U4898 ( .A(n10088), .B(n10618), .Z(n3068) );
  EN U4899 ( .A(n10085), .B(n10618), .Z(n3069) );
  EN U4900 ( .A(n10082), .B(n10618), .Z(n3070) );
  EN U4901 ( .A(n10079), .B(n10618), .Z(n3071) );
  EN U4902 ( .A(n10076), .B(n10618), .Z(n3072) );
  EN U4903 ( .A(n10073), .B(n10618), .Z(n3073) );
  EN U4904 ( .A(n10070), .B(n10618), .Z(n3074) );
  EN U4905 ( .A(n10067), .B(n10618), .Z(n3075) );
  EN U4906 ( .A(n10064), .B(n10618), .Z(n3076) );
  EN U4907 ( .A(n10061), .B(n10618), .Z(n3077) );
  EN U4908 ( .A(n10058), .B(n10618), .Z(n3078) );
  AO4 U4909 ( .A(n10298), .B(n3015), .C(n3016), .D(n10462), .Z(n5181) );
  AO4 U4910 ( .A(n10298), .B(n3016), .C(n3017), .D(n10462), .Z(n5182) );
  AO4 U4911 ( .A(n10298), .B(n3017), .C(n3018), .D(n10462), .Z(n5183) );
  AO4 U4912 ( .A(n10298), .B(n3018), .C(n3019), .D(n10462), .Z(n5184) );
  AO4 U4913 ( .A(n10298), .B(n3019), .C(n3020), .D(n10462), .Z(n5185) );
  AO4 U4914 ( .A(n10298), .B(n3020), .C(n3021), .D(n10462), .Z(n5186) );
  AO4 U4915 ( .A(n10298), .B(n3021), .C(n3022), .D(n10462), .Z(n5187) );
  AO4 U4916 ( .A(n10298), .B(n3022), .C(n3023), .D(n10462), .Z(n5188) );
  AO4 U4917 ( .A(n10298), .B(n3023), .C(n3024), .D(n10462), .Z(n5189) );
  AO4 U4918 ( .A(n10298), .B(n3024), .C(n3025), .D(n10462), .Z(n5190) );
  AO4 U4919 ( .A(n10297), .B(n3025), .C(n3026), .D(n10462), .Z(n5191) );
  AO4 U4920 ( .A(n10297), .B(n3026), .C(n3027), .D(n10461), .Z(n5192) );
  AO4 U4921 ( .A(n10297), .B(n3027), .C(n3028), .D(n10461), .Z(n5193) );
  AO4 U4922 ( .A(n10297), .B(n3028), .C(n3029), .D(n10461), .Z(n5194) );
  AO4 U4923 ( .A(n10297), .B(n3029), .C(n3030), .D(n10461), .Z(n5195) );
  AO4 U4924 ( .A(n10297), .B(n3030), .C(n3031), .D(n10461), .Z(n5196) );
  AO4 U4925 ( .A(n10297), .B(n3031), .C(n3032), .D(n10461), .Z(n5197) );
  AO4 U4926 ( .A(n10297), .B(n3032), .C(n3033), .D(n10461), .Z(n5198) );
  AO4 U4927 ( .A(n10297), .B(n3033), .C(n3034), .D(n10461), .Z(n5199) );
  AO4 U4928 ( .A(n10297), .B(n3034), .C(n3035), .D(n10461), .Z(n5200) );
  AO4 U4929 ( .A(n10297), .B(n3035), .C(n3036), .D(n10461), .Z(n5201) );
  AO4 U4930 ( .A(n10297), .B(n3036), .C(n3037), .D(n10461), .Z(n5202) );
  AO4 U4931 ( .A(n10297), .B(n3037), .C(n3038), .D(n10461), .Z(n5203) );
  AO4 U4932 ( .A(n10297), .B(n3038), .C(n3039), .D(n10461), .Z(n5204) );
  AO4 U4933 ( .A(n10296), .B(n3039), .C(n3040), .D(n10461), .Z(n5205) );
  AO4 U4934 ( .A(n10296), .B(n3040), .C(n3041), .D(n10460), .Z(n5206) );
  AO4 U4935 ( .A(n10296), .B(n3041), .C(n3042), .D(n10460), .Z(n5207) );
  AO4 U4936 ( .A(n10296), .B(n3042), .C(n3043), .D(n10460), .Z(n5208) );
  AO4 U4937 ( .A(n10296), .B(n3043), .C(n3044), .D(n10460), .Z(n5209) );
  AO4 U4938 ( .A(n10296), .B(n3044), .C(n3045), .D(n10460), .Z(n5210) );
  AO4 U4939 ( .A(n10296), .B(n3045), .C(n3046), .D(n10460), .Z(n5211) );
  AO4 U4940 ( .A(n10296), .B(n3046), .C(n3047), .D(n10460), .Z(n5212) );
  AO4 U4941 ( .A(n10296), .B(n3047), .C(n3048), .D(n10460), .Z(n5213) );
  AO4 U4942 ( .A(n10296), .B(n3048), .C(n3049), .D(n10460), .Z(n5214) );
  AO4 U4943 ( .A(n10296), .B(n3049), .C(n3050), .D(n10460), .Z(n5215) );
  AO4 U4944 ( .A(n10296), .B(n3050), .C(n3051), .D(n10460), .Z(n5216) );
  AO4 U4945 ( .A(n10296), .B(n3051), .C(n3052), .D(n10460), .Z(n5217) );
  AO4 U4946 ( .A(n10296), .B(n3052), .C(n3053), .D(n10460), .Z(n5218) );
  AO4 U4947 ( .A(n10295), .B(n3053), .C(n3054), .D(n10460), .Z(n5219) );
  AO4 U4948 ( .A(n10295), .B(n3054), .C(n3055), .D(n10459), .Z(n5220) );
  AO4 U4949 ( .A(n10295), .B(n3055), .C(n3056), .D(n10459), .Z(n5221) );
  AO4 U4950 ( .A(n10295), .B(n3056), .C(n3057), .D(n10459), .Z(n5222) );
  AO4 U4951 ( .A(n10295), .B(n3057), .C(n3058), .D(n10459), .Z(n5223) );
  AO4 U4952 ( .A(n10295), .B(n3058), .C(n3059), .D(n10459), .Z(n5224) );
  AO4 U4953 ( .A(n10295), .B(n3059), .C(n3060), .D(n10459), .Z(n5225) );
  AO4 U4954 ( .A(n10295), .B(n3060), .C(n3061), .D(n10459), .Z(n5226) );
  AO4 U4955 ( .A(n10295), .B(n3061), .C(n3062), .D(n10459), .Z(n5227) );
  AO4 U4956 ( .A(n10295), .B(n3062), .C(n3063), .D(n10459), .Z(n5228) );
  AO4 U4957 ( .A(n10295), .B(n3063), .C(n3064), .D(n10459), .Z(n5229) );
  AO4 U4958 ( .A(n10295), .B(n3064), .C(n3065), .D(n10459), .Z(n5230) );
  AO4 U4959 ( .A(n10295), .B(n3065), .C(n3066), .D(n10459), .Z(n5231) );
  AO4 U4960 ( .A(n10295), .B(n3066), .C(n3067), .D(n10459), .Z(n5232) );
  AO4 U4961 ( .A(n10294), .B(n3067), .C(n3068), .D(n10459), .Z(n5233) );
  AO4 U4962 ( .A(n10294), .B(n3068), .C(n3069), .D(n10458), .Z(n5234) );
  AO4 U4963 ( .A(n10294), .B(n3069), .C(n3070), .D(n10458), .Z(n5235) );
  AO4 U4964 ( .A(n10294), .B(n3070), .C(n3071), .D(n10458), .Z(n5236) );
  AO4 U4965 ( .A(n10294), .B(n3071), .C(n3072), .D(n10458), .Z(n5237) );
  AO4 U4966 ( .A(n10294), .B(n3072), .C(n3073), .D(n10458), .Z(n5238) );
  AO4 U4967 ( .A(n10294), .B(n3073), .C(n3074), .D(n10458), .Z(n5239) );
  AO4 U4968 ( .A(n10294), .B(n3074), .C(n3075), .D(n10458), .Z(n5240) );
  AO4 U4969 ( .A(n10294), .B(n3075), .C(n3076), .D(n10458), .Z(n5241) );
  AO4 U4970 ( .A(n10294), .B(n3076), .C(n3077), .D(n10458), .Z(n5242) );
  AO4 U4971 ( .A(n10294), .B(n3077), .C(n3078), .D(n10458), .Z(n5243) );
  AO4 U4972 ( .A(n10294), .B(n3078), .C(n10458), .D(n1413), .Z(n5244) );
  AO4 U4973 ( .A(n10458), .B(n3014), .C(n10294), .D(n1413), .Z(n5861) );
  EN U4974 ( .A(n10252), .B(n10617), .Z(n3080) );
  EN U4975 ( .A(n10244), .B(n10617), .Z(n3081) );
  EN U4976 ( .A(n10241), .B(n10617), .Z(n3082) );
  EN U4977 ( .A(n10238), .B(n10617), .Z(n3083) );
  EN U4978 ( .A(n10235), .B(n10617), .Z(n3084) );
  EN U4979 ( .A(n10232), .B(n10617), .Z(n3085) );
  EN U4980 ( .A(n10229), .B(n10617), .Z(n3086) );
  EN U4981 ( .A(n10226), .B(n10617), .Z(n3087) );
  EN U4982 ( .A(n10223), .B(n10617), .Z(n3088) );
  EN U4983 ( .A(n10220), .B(n10616), .Z(n3089) );
  EN U4984 ( .A(n10217), .B(n10616), .Z(n3090) );
  EN U4985 ( .A(n10214), .B(n10616), .Z(n3091) );
  EN U4986 ( .A(n10211), .B(n10616), .Z(n3092) );
  EN U4987 ( .A(n10208), .B(n10616), .Z(n3093) );
  EN U4988 ( .A(n10205), .B(n10616), .Z(n3094) );
  EN U4989 ( .A(n10202), .B(n10616), .Z(n3095) );
  EN U4990 ( .A(n10199), .B(n10616), .Z(n3096) );
  EN U4991 ( .A(n10196), .B(n10616), .Z(n3097) );
  EN U4992 ( .A(n10193), .B(n10616), .Z(n3098) );
  EN U4993 ( .A(n10190), .B(n10616), .Z(n3099) );
  EN U4994 ( .A(n10187), .B(n10616), .Z(n3100) );
  EN U4995 ( .A(n10184), .B(n10616), .Z(n3101) );
  EN U4996 ( .A(n10181), .B(n10616), .Z(n3102) );
  EN U4997 ( .A(n10178), .B(n10615), .Z(n3103) );
  EN U4998 ( .A(n10175), .B(n10615), .Z(n3104) );
  EN U4999 ( .A(n10172), .B(n10615), .Z(n3105) );
  EN U5000 ( .A(n10169), .B(n10615), .Z(n3106) );
  EN U5001 ( .A(n10166), .B(n10615), .Z(n3107) );
  EN U5002 ( .A(n10163), .B(n10615), .Z(n3108) );
  EN U5003 ( .A(n10160), .B(n10615), .Z(n3109) );
  EN U5004 ( .A(n10157), .B(n10615), .Z(n3110) );
  EN U5005 ( .A(n10154), .B(n10615), .Z(n3111) );
  EN U5006 ( .A(n10151), .B(n10615), .Z(n3112) );
  EN U5007 ( .A(n10148), .B(n10615), .Z(n3113) );
  EN U5008 ( .A(n10145), .B(n10615), .Z(n3114) );
  EN U5009 ( .A(n10142), .B(n10615), .Z(n3115) );
  EN U5010 ( .A(n10139), .B(n10615), .Z(n3116) );
  EN U5011 ( .A(n10136), .B(n10614), .Z(n3117) );
  EN U5012 ( .A(n10133), .B(n10614), .Z(n3118) );
  EN U5013 ( .A(n10130), .B(n10614), .Z(n3119) );
  EN U5014 ( .A(n10127), .B(n10614), .Z(n3120) );
  EN U5015 ( .A(n10124), .B(n10614), .Z(n3121) );
  EN U5016 ( .A(n10121), .B(n10614), .Z(n3122) );
  EN U5017 ( .A(n10118), .B(n10614), .Z(n3123) );
  EN U5018 ( .A(n10115), .B(n10614), .Z(n3124) );
  EN U5019 ( .A(n10112), .B(n10614), .Z(n3125) );
  EN U5020 ( .A(n10109), .B(n10614), .Z(n3126) );
  EN U5021 ( .A(n10106), .B(n10614), .Z(n3127) );
  EN U5022 ( .A(n10103), .B(n10614), .Z(n3128) );
  EN U5023 ( .A(n10100), .B(n10614), .Z(n3129) );
  EN U5024 ( .A(n10097), .B(n10614), .Z(n3130) );
  EN U5025 ( .A(n10094), .B(n10613), .Z(n3131) );
  EN U5026 ( .A(n10091), .B(n10613), .Z(n3132) );
  EN U5027 ( .A(n10088), .B(n10613), .Z(n3133) );
  EN U5028 ( .A(n10085), .B(n10613), .Z(n3134) );
  EN U5029 ( .A(n10082), .B(n10613), .Z(n3135) );
  EN U5030 ( .A(n10079), .B(n10613), .Z(n3136) );
  EN U5031 ( .A(n10076), .B(n10613), .Z(n3137) );
  EN U5032 ( .A(n10073), .B(n10613), .Z(n3138) );
  EN U5033 ( .A(n10070), .B(n10613), .Z(n3139) );
  EN U5034 ( .A(n10067), .B(n10613), .Z(n3140) );
  EN U5035 ( .A(n10064), .B(n10613), .Z(n3141) );
  EN U5036 ( .A(n10061), .B(n10613), .Z(n3142) );
  EN U5037 ( .A(n10058), .B(n10613), .Z(n3143) );
  AO4 U5038 ( .A(n10293), .B(n3080), .C(n3081), .D(n10457), .Z(n5247) );
  AO4 U5039 ( .A(n10293), .B(n3081), .C(n3082), .D(n10457), .Z(n5248) );
  AO4 U5040 ( .A(n10293), .B(n3082), .C(n3083), .D(n10457), .Z(n5249) );
  AO4 U5041 ( .A(n10293), .B(n3083), .C(n3084), .D(n10457), .Z(n5250) );
  AO4 U5042 ( .A(n10293), .B(n3084), .C(n3085), .D(n10457), .Z(n5251) );
  AO4 U5043 ( .A(n10293), .B(n3085), .C(n3086), .D(n10457), .Z(n5252) );
  AO4 U5044 ( .A(n10293), .B(n3086), .C(n3087), .D(n10457), .Z(n5253) );
  AO4 U5045 ( .A(n10293), .B(n3087), .C(n3088), .D(n10457), .Z(n5254) );
  AO4 U5046 ( .A(n10293), .B(n3088), .C(n3089), .D(n10457), .Z(n5255) );
  AO4 U5047 ( .A(n10293), .B(n3089), .C(n3090), .D(n10457), .Z(n5256) );
  AO4 U5048 ( .A(n10292), .B(n3090), .C(n3091), .D(n10457), .Z(n5257) );
  AO4 U5049 ( .A(n10292), .B(n3091), .C(n3092), .D(n10456), .Z(n5258) );
  AO4 U5050 ( .A(n10292), .B(n3092), .C(n3093), .D(n10456), .Z(n5259) );
  AO4 U5051 ( .A(n10292), .B(n3093), .C(n3094), .D(n10456), .Z(n5260) );
  AO4 U5052 ( .A(n10292), .B(n3094), .C(n3095), .D(n10456), .Z(n5261) );
  AO4 U5053 ( .A(n10292), .B(n3095), .C(n3096), .D(n10456), .Z(n5262) );
  AO4 U5054 ( .A(n10292), .B(n3096), .C(n3097), .D(n10456), .Z(n5263) );
  AO4 U5055 ( .A(n10292), .B(n3097), .C(n3098), .D(n10456), .Z(n5264) );
  AO4 U5056 ( .A(n10292), .B(n3098), .C(n3099), .D(n10456), .Z(n5265) );
  AO4 U5057 ( .A(n10292), .B(n3099), .C(n3100), .D(n10456), .Z(n5266) );
  AO4 U5058 ( .A(n10292), .B(n3100), .C(n3101), .D(n10456), .Z(n5267) );
  AO4 U5059 ( .A(n10292), .B(n3101), .C(n3102), .D(n10456), .Z(n5268) );
  AO4 U5060 ( .A(n10292), .B(n3102), .C(n3103), .D(n10456), .Z(n5269) );
  AO4 U5061 ( .A(n10292), .B(n3103), .C(n3104), .D(n10456), .Z(n5270) );
  AO4 U5062 ( .A(n10291), .B(n3104), .C(n3105), .D(n10456), .Z(n5271) );
  AO4 U5063 ( .A(n10291), .B(n3105), .C(n3106), .D(n10455), .Z(n5272) );
  AO4 U5064 ( .A(n10291), .B(n3106), .C(n3107), .D(n10455), .Z(n5273) );
  AO4 U5065 ( .A(n10291), .B(n3107), .C(n3108), .D(n10455), .Z(n5274) );
  AO4 U5066 ( .A(n10291), .B(n3108), .C(n3109), .D(n10455), .Z(n5275) );
  AO4 U5067 ( .A(n10291), .B(n3109), .C(n3110), .D(n10455), .Z(n5276) );
  AO4 U5068 ( .A(n10291), .B(n3110), .C(n3111), .D(n10455), .Z(n5277) );
  AO4 U5069 ( .A(n10291), .B(n3111), .C(n3112), .D(n10455), .Z(n5278) );
  AO4 U5070 ( .A(n10291), .B(n3112), .C(n3113), .D(n10455), .Z(n5279) );
  AO4 U5071 ( .A(n10291), .B(n3113), .C(n3114), .D(n10455), .Z(n5280) );
  AO4 U5072 ( .A(n10291), .B(n3114), .C(n3115), .D(n10455), .Z(n5281) );
  AO4 U5073 ( .A(n10291), .B(n3115), .C(n3116), .D(n10455), .Z(n5282) );
  AO4 U5074 ( .A(n10291), .B(n3116), .C(n3117), .D(n10455), .Z(n5283) );
  AO4 U5075 ( .A(n10291), .B(n3117), .C(n3118), .D(n10455), .Z(n5284) );
  AO4 U5076 ( .A(n10290), .B(n3118), .C(n3119), .D(n10455), .Z(n5285) );
  AO4 U5077 ( .A(n10290), .B(n3119), .C(n3120), .D(n10454), .Z(n5286) );
  AO4 U5078 ( .A(n10290), .B(n3120), .C(n3121), .D(n10454), .Z(n5287) );
  AO4 U5079 ( .A(n10290), .B(n3121), .C(n3122), .D(n10454), .Z(n5288) );
  AO4 U5080 ( .A(n10290), .B(n3122), .C(n3123), .D(n10454), .Z(n5289) );
  AO4 U5081 ( .A(n10290), .B(n3123), .C(n3124), .D(n10454), .Z(n5290) );
  AO4 U5082 ( .A(n10290), .B(n3124), .C(n3125), .D(n10454), .Z(n5291) );
  AO4 U5083 ( .A(n10290), .B(n3125), .C(n3126), .D(n10454), .Z(n5292) );
  AO4 U5084 ( .A(n10290), .B(n3126), .C(n3127), .D(n10454), .Z(n5293) );
  AO4 U5085 ( .A(n10290), .B(n3127), .C(n3128), .D(n10454), .Z(n5294) );
  AO4 U5086 ( .A(n10290), .B(n3128), .C(n3129), .D(n10454), .Z(n5295) );
  AO4 U5087 ( .A(n10290), .B(n3129), .C(n3130), .D(n10454), .Z(n5296) );
  AO4 U5088 ( .A(n10290), .B(n3130), .C(n3131), .D(n10454), .Z(n5297) );
  AO4 U5089 ( .A(n10290), .B(n3131), .C(n3132), .D(n10454), .Z(n5298) );
  AO4 U5090 ( .A(n10289), .B(n3132), .C(n3133), .D(n10454), .Z(n5299) );
  AO4 U5091 ( .A(n10289), .B(n3133), .C(n3134), .D(n10453), .Z(n5300) );
  AO4 U5092 ( .A(n10289), .B(n3134), .C(n3135), .D(n10453), .Z(n5301) );
  AO4 U5093 ( .A(n10289), .B(n3135), .C(n3136), .D(n10453), .Z(n5302) );
  AO4 U5094 ( .A(n10289), .B(n3136), .C(n3137), .D(n10453), .Z(n5303) );
  AO4 U5095 ( .A(n10289), .B(n3137), .C(n3138), .D(n10453), .Z(n5304) );
  AO4 U5096 ( .A(n10289), .B(n3138), .C(n3139), .D(n10453), .Z(n5305) );
  AO4 U5097 ( .A(n10289), .B(n3139), .C(n3140), .D(n10453), .Z(n5306) );
  AO4 U5098 ( .A(n10289), .B(n3140), .C(n3141), .D(n10453), .Z(n5307) );
  AO4 U5099 ( .A(n10289), .B(n3141), .C(n3142), .D(n10453), .Z(n5308) );
  AO4 U5100 ( .A(n10289), .B(n3142), .C(n3143), .D(n10453), .Z(n5309) );
  AO4 U5101 ( .A(n10289), .B(n3143), .C(n10453), .D(n1414), .Z(n5310) );
  AO4 U5102 ( .A(n10453), .B(n3079), .C(n10289), .D(n1414), .Z(n5862) );
  EN U5103 ( .A(n10252), .B(n10612), .Z(n3145) );
  EN U5104 ( .A(n10244), .B(n10612), .Z(n3146) );
  EN U5105 ( .A(n10241), .B(n10612), .Z(n3147) );
  EN U5106 ( .A(n10238), .B(n10612), .Z(n3148) );
  EN U5107 ( .A(n10235), .B(n10612), .Z(n3149) );
  EN U5108 ( .A(n10232), .B(n10612), .Z(n3150) );
  EN U5109 ( .A(n10229), .B(n10612), .Z(n3151) );
  EN U5110 ( .A(n10226), .B(n10612), .Z(n3152) );
  EN U5111 ( .A(n10223), .B(n10612), .Z(n3153) );
  EN U5112 ( .A(n10220), .B(n10611), .Z(n3154) );
  EN U5113 ( .A(n10217), .B(n10611), .Z(n3155) );
  EN U5114 ( .A(n10214), .B(n10611), .Z(n3156) );
  EN U5115 ( .A(n10211), .B(n10611), .Z(n3157) );
  EN U5116 ( .A(n10208), .B(n10611), .Z(n3158) );
  EN U5117 ( .A(n10205), .B(n10611), .Z(n3159) );
  EN U5118 ( .A(n10202), .B(n10611), .Z(n3160) );
  EN U5119 ( .A(n10199), .B(n10611), .Z(n3161) );
  EN U5120 ( .A(n10196), .B(n10611), .Z(n3162) );
  EN U5121 ( .A(n10193), .B(n10611), .Z(n3163) );
  EN U5122 ( .A(n10190), .B(n10611), .Z(n3164) );
  EN U5123 ( .A(n10187), .B(n10611), .Z(n3165) );
  EN U5124 ( .A(n10184), .B(n10611), .Z(n3166) );
  EN U5125 ( .A(n10181), .B(n10611), .Z(n3167) );
  EN U5126 ( .A(n10178), .B(n10610), .Z(n3168) );
  EN U5127 ( .A(n10175), .B(n10610), .Z(n3169) );
  EN U5128 ( .A(n10172), .B(n10610), .Z(n3170) );
  EN U5129 ( .A(n10169), .B(n10610), .Z(n3171) );
  EN U5130 ( .A(n10166), .B(n10610), .Z(n3172) );
  EN U5131 ( .A(n10163), .B(n10610), .Z(n3173) );
  EN U5132 ( .A(n10160), .B(n10610), .Z(n3174) );
  EN U5133 ( .A(n10157), .B(n10610), .Z(n3175) );
  EN U5134 ( .A(n10154), .B(n10610), .Z(n3176) );
  EN U5135 ( .A(n10151), .B(n10610), .Z(n3177) );
  EN U5136 ( .A(n10148), .B(n10610), .Z(n3178) );
  EN U5137 ( .A(n10145), .B(n10610), .Z(n3179) );
  EN U5138 ( .A(n10142), .B(n10610), .Z(n3180) );
  EN U5139 ( .A(n10139), .B(n10610), .Z(n3181) );
  EN U5140 ( .A(n10136), .B(n10609), .Z(n3182) );
  EN U5141 ( .A(n10133), .B(n10609), .Z(n3183) );
  EN U5142 ( .A(n10130), .B(n10609), .Z(n3184) );
  EN U5143 ( .A(n10127), .B(n10609), .Z(n3185) );
  EN U5144 ( .A(n10124), .B(n10609), .Z(n3186) );
  EN U5145 ( .A(n10121), .B(n10609), .Z(n3187) );
  EN U5146 ( .A(n10118), .B(n10609), .Z(n3188) );
  EN U5147 ( .A(n10115), .B(n10609), .Z(n3189) );
  EN U5148 ( .A(n10112), .B(n10609), .Z(n3190) );
  EN U5149 ( .A(n10109), .B(n10609), .Z(n3191) );
  EN U5150 ( .A(n10106), .B(n10609), .Z(n3192) );
  EN U5151 ( .A(n10103), .B(n10609), .Z(n3193) );
  EN U5152 ( .A(n10100), .B(n10609), .Z(n3194) );
  EN U5153 ( .A(n10097), .B(n10609), .Z(n3195) );
  EN U5154 ( .A(n10094), .B(n10608), .Z(n3196) );
  EN U5155 ( .A(n10091), .B(n10608), .Z(n3197) );
  EN U5156 ( .A(n10088), .B(n10608), .Z(n3198) );
  EN U5157 ( .A(n10085), .B(n10608), .Z(n3199) );
  EN U5158 ( .A(n10082), .B(n10608), .Z(n3200) );
  EN U5159 ( .A(n10079), .B(n10608), .Z(n3201) );
  EN U5160 ( .A(n10076), .B(n10608), .Z(n3202) );
  EN U5161 ( .A(n10073), .B(n10608), .Z(n3203) );
  EN U5162 ( .A(n10070), .B(n10608), .Z(n3204) );
  EN U5163 ( .A(n10067), .B(n10608), .Z(n3205) );
  EN U5164 ( .A(n10064), .B(n10608), .Z(n3206) );
  EN U5165 ( .A(n10061), .B(n10608), .Z(n3207) );
  EN U5166 ( .A(n10058), .B(n10608), .Z(n3208) );
  AO4 U5167 ( .A(n10288), .B(n3145), .C(n3146), .D(n10452), .Z(n5313) );
  AO4 U5168 ( .A(n10288), .B(n3146), .C(n3147), .D(n10452), .Z(n5314) );
  AO4 U5169 ( .A(n10288), .B(n3147), .C(n3148), .D(n10452), .Z(n5315) );
  AO4 U5170 ( .A(n10288), .B(n3148), .C(n3149), .D(n10452), .Z(n5316) );
  AO4 U5171 ( .A(n10288), .B(n3149), .C(n3150), .D(n10452), .Z(n5317) );
  AO4 U5172 ( .A(n10288), .B(n3150), .C(n3151), .D(n10452), .Z(n5318) );
  AO4 U5173 ( .A(n10288), .B(n3151), .C(n3152), .D(n10452), .Z(n5319) );
  AO4 U5174 ( .A(n10288), .B(n3152), .C(n3153), .D(n10452), .Z(n5320) );
  AO4 U5175 ( .A(n10288), .B(n3153), .C(n3154), .D(n10452), .Z(n5321) );
  AO4 U5176 ( .A(n10288), .B(n3154), .C(n3155), .D(n10452), .Z(n5322) );
  AO4 U5177 ( .A(n10287), .B(n3155), .C(n3156), .D(n10452), .Z(n5323) );
  AO4 U5178 ( .A(n10287), .B(n3156), .C(n3157), .D(n10451), .Z(n5324) );
  AO4 U5179 ( .A(n10287), .B(n3157), .C(n3158), .D(n10451), .Z(n5325) );
  AO4 U5180 ( .A(n10287), .B(n3158), .C(n3159), .D(n10451), .Z(n5326) );
  AO4 U5181 ( .A(n10287), .B(n3159), .C(n3160), .D(n10451), .Z(n5327) );
  AO4 U5182 ( .A(n10287), .B(n3160), .C(n3161), .D(n10451), .Z(n5328) );
  AO4 U5183 ( .A(n10287), .B(n3161), .C(n3162), .D(n10451), .Z(n5329) );
  AO4 U5184 ( .A(n10287), .B(n3162), .C(n3163), .D(n10451), .Z(n5330) );
  AO4 U5185 ( .A(n10287), .B(n3163), .C(n3164), .D(n10451), .Z(n5331) );
  AO4 U5186 ( .A(n10287), .B(n3164), .C(n3165), .D(n10451), .Z(n5332) );
  AO4 U5187 ( .A(n10287), .B(n3165), .C(n3166), .D(n10451), .Z(n5333) );
  AO4 U5188 ( .A(n10287), .B(n3166), .C(n3167), .D(n10451), .Z(n5334) );
  AO4 U5189 ( .A(n10287), .B(n3167), .C(n3168), .D(n10451), .Z(n5335) );
  AO4 U5190 ( .A(n10287), .B(n3168), .C(n3169), .D(n10451), .Z(n5336) );
  AO4 U5191 ( .A(n10286), .B(n3169), .C(n3170), .D(n10451), .Z(n5337) );
  AO4 U5192 ( .A(n10286), .B(n3170), .C(n3171), .D(n10450), .Z(n5338) );
  AO4 U5193 ( .A(n10286), .B(n3171), .C(n3172), .D(n10450), .Z(n5339) );
  AO4 U5194 ( .A(n10286), .B(n3172), .C(n3173), .D(n10450), .Z(n5340) );
  AO4 U5195 ( .A(n10286), .B(n3173), .C(n3174), .D(n10450), .Z(n5341) );
  AO4 U5196 ( .A(n10286), .B(n3174), .C(n3175), .D(n10450), .Z(n5342) );
  AO4 U5197 ( .A(n10286), .B(n3175), .C(n3176), .D(n10450), .Z(n5343) );
  AO4 U5198 ( .A(n10286), .B(n3176), .C(n3177), .D(n10450), .Z(n5344) );
  AO4 U5199 ( .A(n10286), .B(n3177), .C(n3178), .D(n10450), .Z(n5345) );
  AO4 U5200 ( .A(n10286), .B(n3178), .C(n3179), .D(n10450), .Z(n5346) );
  AO4 U5201 ( .A(n10286), .B(n3179), .C(n3180), .D(n10450), .Z(n5347) );
  AO4 U5202 ( .A(n10286), .B(n3180), .C(n3181), .D(n10450), .Z(n5348) );
  AO4 U5203 ( .A(n10286), .B(n3181), .C(n3182), .D(n10450), .Z(n5349) );
  AO4 U5204 ( .A(n10286), .B(n3182), .C(n3183), .D(n10450), .Z(n5350) );
  AO4 U5205 ( .A(n10285), .B(n3183), .C(n3184), .D(n10450), .Z(n5351) );
  AO4 U5206 ( .A(n10285), .B(n3184), .C(n3185), .D(n10449), .Z(n5352) );
  AO4 U5207 ( .A(n10285), .B(n3185), .C(n3186), .D(n10449), .Z(n5353) );
  AO4 U5208 ( .A(n10285), .B(n3186), .C(n3187), .D(n10449), .Z(n5354) );
  AO4 U5209 ( .A(n10285), .B(n3187), .C(n3188), .D(n10449), .Z(n5355) );
  AO4 U5210 ( .A(n10285), .B(n3188), .C(n3189), .D(n10449), .Z(n5356) );
  AO4 U5211 ( .A(n10285), .B(n3189), .C(n3190), .D(n10449), .Z(n5357) );
  AO4 U5212 ( .A(n10285), .B(n3190), .C(n3191), .D(n10449), .Z(n5358) );
  AO4 U5213 ( .A(n10285), .B(n3191), .C(n3192), .D(n10449), .Z(n5359) );
  AO4 U5214 ( .A(n10285), .B(n3192), .C(n3193), .D(n10449), .Z(n5360) );
  AO4 U5215 ( .A(n10285), .B(n3193), .C(n3194), .D(n10449), .Z(n5361) );
  AO4 U5216 ( .A(n10285), .B(n3194), .C(n3195), .D(n10449), .Z(n5362) );
  AO4 U5217 ( .A(n10285), .B(n3195), .C(n3196), .D(n10449), .Z(n5363) );
  AO4 U5218 ( .A(n10285), .B(n3196), .C(n3197), .D(n10449), .Z(n5364) );
  AO4 U5219 ( .A(n10284), .B(n3197), .C(n3198), .D(n10449), .Z(n5365) );
  AO4 U5220 ( .A(n10284), .B(n3198), .C(n3199), .D(n10448), .Z(n5366) );
  AO4 U5221 ( .A(n10284), .B(n3199), .C(n3200), .D(n10448), .Z(n5367) );
  AO4 U5222 ( .A(n10284), .B(n3200), .C(n3201), .D(n10448), .Z(n5368) );
  AO4 U5223 ( .A(n10284), .B(n3201), .C(n3202), .D(n10448), .Z(n5369) );
  AO4 U5224 ( .A(n10284), .B(n3202), .C(n3203), .D(n10448), .Z(n5370) );
  AO4 U5225 ( .A(n10284), .B(n3203), .C(n3204), .D(n10448), .Z(n5371) );
  AO4 U5226 ( .A(n10284), .B(n3204), .C(n3205), .D(n10448), .Z(n5372) );
  AO4 U5227 ( .A(n10284), .B(n3205), .C(n3206), .D(n10448), .Z(n5373) );
  AO4 U5228 ( .A(n10284), .B(n3206), .C(n3207), .D(n10448), .Z(n5374) );
  AO4 U5229 ( .A(n10284), .B(n3207), .C(n3208), .D(n10448), .Z(n5375) );
  AO4 U5230 ( .A(n10284), .B(n3208), .C(n10448), .D(n1415), .Z(n5376) );
  AO4 U5231 ( .A(n10448), .B(n3144), .C(n10284), .D(n1415), .Z(n5863) );
  EN U5232 ( .A(n10252), .B(n10607), .Z(n3210) );
  EN U5233 ( .A(n10244), .B(n10607), .Z(n3211) );
  EN U5234 ( .A(n10241), .B(n10607), .Z(n3212) );
  EN U5235 ( .A(n10238), .B(n10607), .Z(n3213) );
  EN U5236 ( .A(n10235), .B(n10607), .Z(n3214) );
  EN U5237 ( .A(n10232), .B(n10607), .Z(n3215) );
  EN U5238 ( .A(n10229), .B(n10607), .Z(n3216) );
  EN U5239 ( .A(n10226), .B(n10607), .Z(n3217) );
  EN U5240 ( .A(n10223), .B(n10607), .Z(n3218) );
  EN U5241 ( .A(n10220), .B(n10606), .Z(n3219) );
  EN U5242 ( .A(n10217), .B(n10606), .Z(n3220) );
  EN U5243 ( .A(n10214), .B(n10606), .Z(n3221) );
  EN U5244 ( .A(n10211), .B(n10606), .Z(n3222) );
  EN U5245 ( .A(n10208), .B(n10606), .Z(n3223) );
  EN U5246 ( .A(n10205), .B(n10606), .Z(n3224) );
  EN U5247 ( .A(n10202), .B(n10606), .Z(n3225) );
  EN U5248 ( .A(n10199), .B(n10606), .Z(n3226) );
  EN U5249 ( .A(n10196), .B(n10606), .Z(n3227) );
  EN U5250 ( .A(n10193), .B(n10606), .Z(n3228) );
  EN U5251 ( .A(n10190), .B(n10606), .Z(n3229) );
  EN U5252 ( .A(n10187), .B(n10606), .Z(n3230) );
  EN U5253 ( .A(n10184), .B(n10606), .Z(n3231) );
  EN U5254 ( .A(n10181), .B(n10606), .Z(n3232) );
  EN U5255 ( .A(n10178), .B(n10605), .Z(n3233) );
  EN U5256 ( .A(n10175), .B(n10605), .Z(n3234) );
  EN U5257 ( .A(n10172), .B(n10605), .Z(n3235) );
  EN U5258 ( .A(n10169), .B(n10605), .Z(n3236) );
  EN U5259 ( .A(n10166), .B(n10605), .Z(n3237) );
  EN U5260 ( .A(n10163), .B(n10605), .Z(n3238) );
  EN U5261 ( .A(n10160), .B(n10605), .Z(n3239) );
  EN U5262 ( .A(n10157), .B(n10605), .Z(n3240) );
  EN U5263 ( .A(n10154), .B(n10605), .Z(n3241) );
  EN U5264 ( .A(n10151), .B(n10605), .Z(n3242) );
  EN U5265 ( .A(n10148), .B(n10605), .Z(n3243) );
  EN U5266 ( .A(n10145), .B(n10605), .Z(n3244) );
  EN U5267 ( .A(n10142), .B(n10605), .Z(n3245) );
  EN U5268 ( .A(n10139), .B(n10605), .Z(n3246) );
  EN U5269 ( .A(n10136), .B(n10604), .Z(n3247) );
  EN U5270 ( .A(n10133), .B(n10604), .Z(n3248) );
  EN U5271 ( .A(n10130), .B(n10604), .Z(n3249) );
  EN U5272 ( .A(n10127), .B(n10604), .Z(n3250) );
  EN U5273 ( .A(n10124), .B(n10604), .Z(n3251) );
  EN U5274 ( .A(n10121), .B(n10604), .Z(n3252) );
  EN U5275 ( .A(n10118), .B(n10604), .Z(n3253) );
  EN U5276 ( .A(n10115), .B(n10604), .Z(n3254) );
  EN U5277 ( .A(n10112), .B(n10604), .Z(n3255) );
  EN U5278 ( .A(n10109), .B(n10604), .Z(n3256) );
  EN U5279 ( .A(n10106), .B(n10604), .Z(n3257) );
  EN U5280 ( .A(n10103), .B(n10604), .Z(n3258) );
  EN U5281 ( .A(n10100), .B(n10604), .Z(n3259) );
  EN U5282 ( .A(n10097), .B(n10604), .Z(n3260) );
  EN U5283 ( .A(n10094), .B(n10603), .Z(n3261) );
  EN U5284 ( .A(n10091), .B(n10603), .Z(n3262) );
  EN U5285 ( .A(n10088), .B(n10603), .Z(n3263) );
  EN U5286 ( .A(n10085), .B(n10603), .Z(n3264) );
  EN U5287 ( .A(n10082), .B(n10603), .Z(n3265) );
  EN U5288 ( .A(n10079), .B(n10603), .Z(n3266) );
  EN U5289 ( .A(n10076), .B(n10603), .Z(n3267) );
  EN U5290 ( .A(n10073), .B(n10603), .Z(n3268) );
  EN U5291 ( .A(n10070), .B(n10603), .Z(n3269) );
  EN U5292 ( .A(n10067), .B(n10603), .Z(n3270) );
  EN U5293 ( .A(n10064), .B(n10603), .Z(n3271) );
  EN U5294 ( .A(n10061), .B(n10603), .Z(n3272) );
  EN U5295 ( .A(n10058), .B(n10603), .Z(n3273) );
  AO4 U5296 ( .A(n10283), .B(n3210), .C(n3211), .D(n10447), .Z(n5379) );
  AO4 U5297 ( .A(n10283), .B(n3211), .C(n3212), .D(n10447), .Z(n5380) );
  AO4 U5298 ( .A(n10283), .B(n3212), .C(n3213), .D(n10447), .Z(n5381) );
  AO4 U5299 ( .A(n10283), .B(n3213), .C(n3214), .D(n10447), .Z(n5382) );
  AO4 U5300 ( .A(n10283), .B(n3214), .C(n3215), .D(n10447), .Z(n5383) );
  AO4 U5301 ( .A(n10283), .B(n3215), .C(n3216), .D(n10447), .Z(n5384) );
  AO4 U5302 ( .A(n10283), .B(n3216), .C(n3217), .D(n10447), .Z(n5385) );
  AO4 U5303 ( .A(n10283), .B(n3217), .C(n3218), .D(n10447), .Z(n5386) );
  AO4 U5304 ( .A(n10283), .B(n3218), .C(n3219), .D(n10447), .Z(n5387) );
  AO4 U5305 ( .A(n10283), .B(n3219), .C(n3220), .D(n10447), .Z(n5388) );
  AO4 U5306 ( .A(n10282), .B(n3220), .C(n3221), .D(n10447), .Z(n5389) );
  AO4 U5307 ( .A(n10282), .B(n3221), .C(n3222), .D(n10446), .Z(n5390) );
  AO4 U5308 ( .A(n10282), .B(n3222), .C(n3223), .D(n10446), .Z(n5391) );
  AO4 U5309 ( .A(n10282), .B(n3223), .C(n3224), .D(n10446), .Z(n5392) );
  AO4 U5310 ( .A(n10282), .B(n3224), .C(n3225), .D(n10446), .Z(n5393) );
  AO4 U5311 ( .A(n10282), .B(n3225), .C(n3226), .D(n10446), .Z(n5394) );
  AO4 U5312 ( .A(n10282), .B(n3226), .C(n3227), .D(n10446), .Z(n5395) );
  AO4 U5313 ( .A(n10282), .B(n3227), .C(n3228), .D(n10446), .Z(n5396) );
  AO4 U5314 ( .A(n10282), .B(n3228), .C(n3229), .D(n10446), .Z(n5397) );
  AO4 U5315 ( .A(n10282), .B(n3229), .C(n3230), .D(n10446), .Z(n5398) );
  AO4 U5316 ( .A(n10282), .B(n3230), .C(n3231), .D(n10446), .Z(n5399) );
  AO4 U5317 ( .A(n10282), .B(n3231), .C(n3232), .D(n10446), .Z(n5400) );
  AO4 U5318 ( .A(n10282), .B(n3232), .C(n3233), .D(n10446), .Z(n5401) );
  AO4 U5319 ( .A(n10282), .B(n3233), .C(n3234), .D(n10446), .Z(n5402) );
  AO4 U5320 ( .A(n10281), .B(n3234), .C(n3235), .D(n10446), .Z(n5403) );
  AO4 U5321 ( .A(n10281), .B(n3235), .C(n3236), .D(n10445), .Z(n5404) );
  AO4 U5322 ( .A(n10281), .B(n3236), .C(n3237), .D(n10445), .Z(n5405) );
  AO4 U5323 ( .A(n10281), .B(n3237), .C(n3238), .D(n10445), .Z(n5406) );
  AO4 U5324 ( .A(n10281), .B(n3238), .C(n3239), .D(n10445), .Z(n5407) );
  AO4 U5325 ( .A(n10281), .B(n3239), .C(n3240), .D(n10445), .Z(n5408) );
  AO4 U5326 ( .A(n10281), .B(n3240), .C(n3241), .D(n10445), .Z(n5409) );
  AO4 U5327 ( .A(n10281), .B(n3241), .C(n3242), .D(n10445), .Z(n5410) );
  AO4 U5328 ( .A(n10281), .B(n3242), .C(n3243), .D(n10445), .Z(n5411) );
  AO4 U5329 ( .A(n10281), .B(n3243), .C(n3244), .D(n10445), .Z(n5412) );
  AO4 U5330 ( .A(n10281), .B(n3244), .C(n3245), .D(n10445), .Z(n5413) );
  AO4 U5331 ( .A(n10281), .B(n3245), .C(n3246), .D(n10445), .Z(n5414) );
  AO4 U5332 ( .A(n10281), .B(n3246), .C(n3247), .D(n10445), .Z(n5415) );
  AO4 U5333 ( .A(n10281), .B(n3247), .C(n3248), .D(n10445), .Z(n5416) );
  AO4 U5334 ( .A(n10280), .B(n3248), .C(n3249), .D(n10445), .Z(n5417) );
  AO4 U5335 ( .A(n10280), .B(n3249), .C(n3250), .D(n10444), .Z(n5418) );
  AO4 U5336 ( .A(n10280), .B(n3250), .C(n3251), .D(n10444), .Z(n5419) );
  AO4 U5337 ( .A(n10280), .B(n3251), .C(n3252), .D(n10444), .Z(n5420) );
  AO4 U5338 ( .A(n10280), .B(n3252), .C(n3253), .D(n10444), .Z(n5421) );
  AO4 U5339 ( .A(n10280), .B(n3253), .C(n3254), .D(n10444), .Z(n5422) );
  AO4 U5340 ( .A(n10280), .B(n3254), .C(n3255), .D(n10444), .Z(n5423) );
  AO4 U5341 ( .A(n10280), .B(n3255), .C(n3256), .D(n10444), .Z(n5424) );
  AO4 U5342 ( .A(n10280), .B(n3256), .C(n3257), .D(n10444), .Z(n5425) );
  AO4 U5343 ( .A(n10280), .B(n3257), .C(n3258), .D(n10444), .Z(n5426) );
  AO4 U5344 ( .A(n10280), .B(n3258), .C(n3259), .D(n10444), .Z(n5427) );
  AO4 U5345 ( .A(n10280), .B(n3259), .C(n3260), .D(n10444), .Z(n5428) );
  AO4 U5346 ( .A(n10280), .B(n3260), .C(n3261), .D(n10444), .Z(n5429) );
  AO4 U5347 ( .A(n10280), .B(n3261), .C(n3262), .D(n10444), .Z(n5430) );
  AO4 U5348 ( .A(n10279), .B(n3262), .C(n3263), .D(n10444), .Z(n5431) );
  AO4 U5349 ( .A(n10279), .B(n3263), .C(n3264), .D(n10443), .Z(n5432) );
  AO4 U5350 ( .A(n10279), .B(n3264), .C(n3265), .D(n10443), .Z(n5433) );
  AO4 U5351 ( .A(n10279), .B(n3265), .C(n3266), .D(n10443), .Z(n5434) );
  AO4 U5352 ( .A(n10279), .B(n3266), .C(n3267), .D(n10443), .Z(n5435) );
  AO4 U5353 ( .A(n10279), .B(n3267), .C(n3268), .D(n10443), .Z(n5436) );
  AO4 U5354 ( .A(n10279), .B(n3268), .C(n3269), .D(n10443), .Z(n5437) );
  AO4 U5355 ( .A(n10279), .B(n3269), .C(n3270), .D(n10443), .Z(n5438) );
  AO4 U5356 ( .A(n10279), .B(n3270), .C(n3271), .D(n10443), .Z(n5439) );
  AO4 U5357 ( .A(n10279), .B(n3271), .C(n3272), .D(n10443), .Z(n5440) );
  AO4 U5358 ( .A(n10279), .B(n3272), .C(n3273), .D(n10443), .Z(n5441) );
  AO4 U5359 ( .A(n10279), .B(n3273), .C(n10443), .D(n1416), .Z(n5442) );
  AO4 U5360 ( .A(n10443), .B(n3209), .C(n10279), .D(n1416), .Z(n5864) );
  EN U5361 ( .A(n10252), .B(n10602), .Z(n3275) );
  EN U5362 ( .A(n10244), .B(n10602), .Z(n3276) );
  EN U5363 ( .A(n10241), .B(n10602), .Z(n3277) );
  EN U5364 ( .A(n10238), .B(n10602), .Z(n3278) );
  EN U5365 ( .A(n10235), .B(n10602), .Z(n3279) );
  EN U5366 ( .A(n10232), .B(n10602), .Z(n3280) );
  EN U5367 ( .A(n10229), .B(n10602), .Z(n3281) );
  EN U5368 ( .A(n10226), .B(n10602), .Z(n3282) );
  EN U5369 ( .A(n10223), .B(n10602), .Z(n3283) );
  EN U5370 ( .A(n10220), .B(n10601), .Z(n3284) );
  EN U5371 ( .A(n10217), .B(n10601), .Z(n3285) );
  EN U5372 ( .A(n10214), .B(n10601), .Z(n3286) );
  EN U5373 ( .A(n10211), .B(n10601), .Z(n3287) );
  EN U5374 ( .A(n10208), .B(n10601), .Z(n3288) );
  EN U5375 ( .A(n10205), .B(n10601), .Z(n3289) );
  EN U5376 ( .A(n10202), .B(n10601), .Z(n3290) );
  EN U5377 ( .A(n10199), .B(n10601), .Z(n3291) );
  EN U5378 ( .A(n10196), .B(n10601), .Z(n3292) );
  EN U5379 ( .A(n10193), .B(n10601), .Z(n3293) );
  EN U5380 ( .A(n10190), .B(n10601), .Z(n3294) );
  EN U5381 ( .A(n10187), .B(n10601), .Z(n3295) );
  EN U5382 ( .A(n10184), .B(n10601), .Z(n3296) );
  EN U5383 ( .A(n10181), .B(n10601), .Z(n3297) );
  EN U5384 ( .A(n10178), .B(n10600), .Z(n3298) );
  EN U5385 ( .A(n10175), .B(n10600), .Z(n3299) );
  EN U5386 ( .A(n10172), .B(n10600), .Z(n3300) );
  EN U5387 ( .A(n10169), .B(n10600), .Z(n3301) );
  EN U5388 ( .A(n10166), .B(n10600), .Z(n3302) );
  EN U5389 ( .A(n10163), .B(n10600), .Z(n3303) );
  EN U5390 ( .A(n10160), .B(n10600), .Z(n3304) );
  EN U5391 ( .A(n10157), .B(n10600), .Z(n3305) );
  EN U5392 ( .A(n10154), .B(n10600), .Z(n3306) );
  EN U5393 ( .A(n10151), .B(n10600), .Z(n3307) );
  EN U5394 ( .A(n10148), .B(n10600), .Z(n3308) );
  EN U5395 ( .A(n10145), .B(n10600), .Z(n3309) );
  EN U5396 ( .A(n10142), .B(n10600), .Z(n3310) );
  EN U5397 ( .A(n10139), .B(n10600), .Z(n3311) );
  EN U5398 ( .A(n10136), .B(n10599), .Z(n3312) );
  EN U5399 ( .A(n10133), .B(n10599), .Z(n3313) );
  EN U5400 ( .A(n10130), .B(n10599), .Z(n3314) );
  EN U5401 ( .A(n10127), .B(n10599), .Z(n3315) );
  EN U5402 ( .A(n10124), .B(n10599), .Z(n3316) );
  EN U5403 ( .A(n10121), .B(n10599), .Z(n3317) );
  EN U5404 ( .A(n10118), .B(n10599), .Z(n3318) );
  EN U5405 ( .A(n10115), .B(n10599), .Z(n3319) );
  EN U5406 ( .A(n10112), .B(n10599), .Z(n3320) );
  EN U5407 ( .A(n10109), .B(n10599), .Z(n3321) );
  EN U5408 ( .A(n10106), .B(n10599), .Z(n3322) );
  EN U5409 ( .A(n10103), .B(n10599), .Z(n3323) );
  EN U5410 ( .A(n10100), .B(n10599), .Z(n3324) );
  EN U5411 ( .A(n10097), .B(n10599), .Z(n3325) );
  EN U5412 ( .A(n10094), .B(n10598), .Z(n3326) );
  EN U5413 ( .A(n10091), .B(n10598), .Z(n3327) );
  EN U5414 ( .A(n10088), .B(n10598), .Z(n3328) );
  EN U5415 ( .A(n10085), .B(n10598), .Z(n3329) );
  EN U5416 ( .A(n10082), .B(n10598), .Z(n3330) );
  EN U5417 ( .A(n10079), .B(n10598), .Z(n3331) );
  EN U5418 ( .A(n10076), .B(n10598), .Z(n3332) );
  EN U5419 ( .A(n10073), .B(n10598), .Z(n3333) );
  EN U5420 ( .A(n10070), .B(n10598), .Z(n3334) );
  EN U5421 ( .A(n10067), .B(n10598), .Z(n3335) );
  EN U5422 ( .A(n10064), .B(n10598), .Z(n3336) );
  EN U5423 ( .A(n10061), .B(n10598), .Z(n3337) );
  EN U5424 ( .A(n10058), .B(n10598), .Z(n3338) );
  AO4 U5425 ( .A(n10278), .B(n3275), .C(n3276), .D(n10442), .Z(n5445) );
  AO4 U5426 ( .A(n10278), .B(n3276), .C(n3277), .D(n10442), .Z(n5446) );
  AO4 U5427 ( .A(n10278), .B(n3277), .C(n3278), .D(n10442), .Z(n5447) );
  AO4 U5428 ( .A(n10278), .B(n3278), .C(n3279), .D(n10442), .Z(n5448) );
  AO4 U5429 ( .A(n10278), .B(n3279), .C(n3280), .D(n10442), .Z(n5449) );
  AO4 U5430 ( .A(n10278), .B(n3280), .C(n3281), .D(n10442), .Z(n5450) );
  AO4 U5431 ( .A(n10278), .B(n3281), .C(n3282), .D(n10442), .Z(n5451) );
  AO4 U5432 ( .A(n10278), .B(n3282), .C(n3283), .D(n10442), .Z(n5452) );
  AO4 U5433 ( .A(n10278), .B(n3283), .C(n3284), .D(n10442), .Z(n5453) );
  AO4 U5434 ( .A(n10278), .B(n3284), .C(n3285), .D(n10442), .Z(n5454) );
  AO4 U5435 ( .A(n10277), .B(n3285), .C(n3286), .D(n10442), .Z(n5455) );
  AO4 U5436 ( .A(n10277), .B(n3286), .C(n3287), .D(n10441), .Z(n5456) );
  AO4 U5437 ( .A(n10277), .B(n3287), .C(n3288), .D(n10441), .Z(n5457) );
  AO4 U5438 ( .A(n10277), .B(n3288), .C(n3289), .D(n10441), .Z(n5458) );
  AO4 U5439 ( .A(n10277), .B(n3289), .C(n3290), .D(n10441), .Z(n5459) );
  AO4 U5440 ( .A(n10277), .B(n3290), .C(n3291), .D(n10441), .Z(n5460) );
  AO4 U5441 ( .A(n10277), .B(n3291), .C(n3292), .D(n10441), .Z(n5461) );
  AO4 U5442 ( .A(n10277), .B(n3292), .C(n3293), .D(n10441), .Z(n5462) );
  AO4 U5443 ( .A(n10277), .B(n3293), .C(n3294), .D(n10441), .Z(n5463) );
  AO4 U5444 ( .A(n10277), .B(n3294), .C(n3295), .D(n10441), .Z(n5464) );
  AO4 U5445 ( .A(n10277), .B(n3295), .C(n3296), .D(n10441), .Z(n5465) );
  AO4 U5446 ( .A(n10277), .B(n3296), .C(n3297), .D(n10441), .Z(n5466) );
  AO4 U5447 ( .A(n10277), .B(n3297), .C(n3298), .D(n10441), .Z(n5467) );
  AO4 U5448 ( .A(n10277), .B(n3298), .C(n3299), .D(n10441), .Z(n5468) );
  AO4 U5449 ( .A(n10276), .B(n3299), .C(n3300), .D(n10441), .Z(n5469) );
  AO4 U5450 ( .A(n10276), .B(n3300), .C(n3301), .D(n10440), .Z(n5470) );
  AO4 U5451 ( .A(n10276), .B(n3301), .C(n3302), .D(n10440), .Z(n5471) );
  AO4 U5452 ( .A(n10276), .B(n3302), .C(n3303), .D(n10440), .Z(n5472) );
  AO4 U5453 ( .A(n10276), .B(n3303), .C(n3304), .D(n10440), .Z(n5473) );
  AO4 U5454 ( .A(n10276), .B(n3304), .C(n3305), .D(n10440), .Z(n5474) );
  AO4 U5455 ( .A(n10276), .B(n3305), .C(n3306), .D(n10440), .Z(n5475) );
  AO4 U5456 ( .A(n10276), .B(n3306), .C(n3307), .D(n10440), .Z(n5476) );
  AO4 U5457 ( .A(n10276), .B(n3307), .C(n3308), .D(n10440), .Z(n5477) );
  AO4 U5458 ( .A(n10276), .B(n3308), .C(n3309), .D(n10440), .Z(n5478) );
  AO4 U5459 ( .A(n10276), .B(n3309), .C(n3310), .D(n10440), .Z(n5479) );
  AO4 U5460 ( .A(n10276), .B(n3310), .C(n3311), .D(n10440), .Z(n5480) );
  AO4 U5461 ( .A(n10276), .B(n3311), .C(n3312), .D(n10440), .Z(n5481) );
  AO4 U5462 ( .A(n10276), .B(n3312), .C(n3313), .D(n10440), .Z(n5482) );
  AO4 U5463 ( .A(n10275), .B(n3313), .C(n3314), .D(n10440), .Z(n5483) );
  AO4 U5464 ( .A(n10275), .B(n3314), .C(n3315), .D(n10439), .Z(n5484) );
  AO4 U5465 ( .A(n10275), .B(n3315), .C(n3316), .D(n10439), .Z(n5485) );
  AO4 U5466 ( .A(n10275), .B(n3316), .C(n3317), .D(n10439), .Z(n5486) );
  AO4 U5467 ( .A(n10275), .B(n3317), .C(n3318), .D(n10439), .Z(n5487) );
  AO4 U5468 ( .A(n10275), .B(n3318), .C(n3319), .D(n10439), .Z(n5488) );
  AO4 U5469 ( .A(n10275), .B(n3319), .C(n3320), .D(n10439), .Z(n5489) );
  AO4 U5470 ( .A(n10275), .B(n3320), .C(n3321), .D(n10439), .Z(n5490) );
  AO4 U5471 ( .A(n10275), .B(n3321), .C(n3322), .D(n10439), .Z(n5491) );
  AO4 U5472 ( .A(n10275), .B(n3322), .C(n3323), .D(n10439), .Z(n5492) );
  AO4 U5473 ( .A(n10275), .B(n3323), .C(n3324), .D(n10439), .Z(n5493) );
  AO4 U5474 ( .A(n10275), .B(n3324), .C(n3325), .D(n10439), .Z(n5494) );
  AO4 U5475 ( .A(n10275), .B(n3325), .C(n3326), .D(n10439), .Z(n5495) );
  AO4 U5476 ( .A(n10275), .B(n3326), .C(n3327), .D(n10439), .Z(n5496) );
  AO4 U5477 ( .A(n10274), .B(n3327), .C(n3328), .D(n10439), .Z(n5497) );
  AO4 U5478 ( .A(n10274), .B(n3328), .C(n3329), .D(n10438), .Z(n5498) );
  AO4 U5479 ( .A(n10274), .B(n3329), .C(n3330), .D(n10438), .Z(n5499) );
  AO4 U5480 ( .A(n10274), .B(n3330), .C(n3331), .D(n10438), .Z(n5500) );
  AO4 U5481 ( .A(n10274), .B(n3331), .C(n3332), .D(n10438), .Z(n5501) );
  AO4 U5482 ( .A(n10274), .B(n3332), .C(n3333), .D(n10438), .Z(n5502) );
  AO4 U5483 ( .A(n10274), .B(n3333), .C(n3334), .D(n10438), .Z(n5503) );
  AO4 U5484 ( .A(n10274), .B(n3334), .C(n3335), .D(n10438), .Z(n5504) );
  AO4 U5485 ( .A(n10274), .B(n3335), .C(n3336), .D(n10438), .Z(n5505) );
  AO4 U5486 ( .A(n10274), .B(n3336), .C(n3337), .D(n10438), .Z(n5506) );
  AO4 U5487 ( .A(n10274), .B(n3337), .C(n3338), .D(n10438), .Z(n5507) );
  AO4 U5488 ( .A(n10274), .B(n3338), .C(n10438), .D(n1417), .Z(n5508) );
  AO4 U5489 ( .A(n10438), .B(n3274), .C(n10274), .D(n1417), .Z(n5865) );
  EN U5490 ( .A(n10251), .B(n10597), .Z(n3340) );
  EN U5491 ( .A(n10244), .B(n10597), .Z(n3341) );
  EN U5492 ( .A(n10241), .B(n10597), .Z(n3342) );
  EN U5493 ( .A(n10238), .B(n10597), .Z(n3343) );
  EN U5494 ( .A(n10235), .B(n10597), .Z(n3344) );
  EN U5495 ( .A(n10232), .B(n10597), .Z(n3345) );
  EN U5496 ( .A(n10229), .B(n10597), .Z(n3346) );
  EN U5497 ( .A(n10226), .B(n10597), .Z(n3347) );
  EN U5498 ( .A(n10223), .B(n10597), .Z(n3348) );
  EN U5499 ( .A(n10220), .B(n10596), .Z(n3349) );
  EN U5500 ( .A(n10217), .B(n10596), .Z(n3350) );
  EN U5501 ( .A(n10214), .B(n10596), .Z(n3351) );
  EN U5502 ( .A(n10211), .B(n10596), .Z(n3352) );
  EN U5503 ( .A(n10208), .B(n10596), .Z(n3353) );
  EN U5504 ( .A(n10205), .B(n10596), .Z(n3354) );
  EN U5505 ( .A(n10202), .B(n10596), .Z(n3355) );
  EN U5506 ( .A(n10199), .B(n10596), .Z(n3356) );
  EN U5507 ( .A(n10196), .B(n10596), .Z(n3357) );
  EN U5508 ( .A(n10193), .B(n10596), .Z(n3358) );
  EN U5509 ( .A(n10190), .B(n10596), .Z(n3359) );
  EN U5510 ( .A(n10187), .B(n10596), .Z(n3360) );
  EN U5511 ( .A(n10184), .B(n10596), .Z(n3361) );
  EN U5512 ( .A(n10181), .B(n10596), .Z(n3362) );
  EN U5513 ( .A(n10178), .B(n10595), .Z(n3363) );
  EN U5514 ( .A(n10175), .B(n10595), .Z(n3364) );
  EN U5515 ( .A(n10172), .B(n10595), .Z(n3365) );
  EN U5516 ( .A(n10169), .B(n10595), .Z(n3366) );
  EN U5517 ( .A(n10166), .B(n10595), .Z(n3367) );
  EN U5518 ( .A(n10163), .B(n10595), .Z(n3368) );
  EN U5519 ( .A(n10160), .B(n10595), .Z(n3369) );
  EN U5520 ( .A(n10157), .B(n10595), .Z(n3370) );
  EN U5521 ( .A(n10154), .B(n10595), .Z(n3371) );
  EN U5522 ( .A(n10151), .B(n10595), .Z(n3372) );
  EN U5523 ( .A(n10148), .B(n10595), .Z(n3373) );
  EN U5524 ( .A(n10145), .B(n10595), .Z(n3374) );
  EN U5525 ( .A(n10142), .B(n10595), .Z(n3375) );
  EN U5526 ( .A(n10139), .B(n10595), .Z(n3376) );
  EN U5527 ( .A(n10136), .B(n10594), .Z(n3377) );
  EN U5528 ( .A(n10133), .B(n10594), .Z(n3378) );
  EN U5529 ( .A(n10130), .B(n10594), .Z(n3379) );
  EN U5530 ( .A(n10127), .B(n10594), .Z(n3380) );
  EN U5531 ( .A(n10124), .B(n10594), .Z(n3381) );
  EN U5532 ( .A(n10121), .B(n10594), .Z(n3382) );
  EN U5533 ( .A(n10118), .B(n10594), .Z(n3383) );
  EN U5534 ( .A(n10115), .B(n10594), .Z(n3384) );
  EN U5535 ( .A(n10112), .B(n10594), .Z(n3385) );
  EN U5536 ( .A(n10109), .B(n10594), .Z(n3386) );
  EN U5537 ( .A(n10106), .B(n10594), .Z(n3387) );
  EN U5538 ( .A(n10103), .B(n10594), .Z(n3388) );
  EN U5539 ( .A(n10100), .B(n10594), .Z(n3389) );
  EN U5540 ( .A(n10097), .B(n10594), .Z(n3390) );
  EN U5541 ( .A(n10094), .B(n10593), .Z(n3391) );
  EN U5542 ( .A(n10091), .B(n10593), .Z(n3392) );
  EN U5543 ( .A(n10088), .B(n10593), .Z(n3393) );
  EN U5544 ( .A(n10085), .B(n10593), .Z(n3394) );
  EN U5545 ( .A(n10082), .B(n10593), .Z(n3395) );
  EN U5546 ( .A(n10079), .B(n10593), .Z(n3396) );
  EN U5547 ( .A(n10076), .B(n10593), .Z(n3397) );
  EN U5548 ( .A(n10073), .B(n10593), .Z(n3398) );
  EN U5549 ( .A(n10070), .B(n10593), .Z(n3399) );
  EN U5550 ( .A(n10067), .B(n10593), .Z(n3400) );
  EN U5551 ( .A(n10064), .B(n10593), .Z(n3401) );
  EN U5552 ( .A(n10061), .B(n10593), .Z(n3402) );
  EN U5553 ( .A(n10058), .B(n10593), .Z(n3403) );
  AO4 U5554 ( .A(n10273), .B(n3340), .C(n3341), .D(n10437), .Z(n5511) );
  AO4 U5555 ( .A(n10273), .B(n3341), .C(n3342), .D(n10437), .Z(n5512) );
  AO4 U5556 ( .A(n10273), .B(n3342), .C(n3343), .D(n10437), .Z(n5513) );
  AO4 U5557 ( .A(n10273), .B(n3343), .C(n3344), .D(n10437), .Z(n5514) );
  AO4 U5558 ( .A(n10273), .B(n3344), .C(n3345), .D(n10437), .Z(n5515) );
  AO4 U5559 ( .A(n10273), .B(n3345), .C(n3346), .D(n10437), .Z(n5516) );
  AO4 U5560 ( .A(n10273), .B(n3346), .C(n3347), .D(n10437), .Z(n5517) );
  AO4 U5561 ( .A(n10273), .B(n3347), .C(n3348), .D(n10437), .Z(n5518) );
  AO4 U5562 ( .A(n10273), .B(n3348), .C(n3349), .D(n10437), .Z(n5519) );
  AO4 U5563 ( .A(n10273), .B(n3349), .C(n3350), .D(n10437), .Z(n5520) );
  AO4 U5564 ( .A(n10272), .B(n3350), .C(n3351), .D(n10437), .Z(n5521) );
  AO4 U5565 ( .A(n10272), .B(n3351), .C(n3352), .D(n10436), .Z(n5522) );
  AO4 U5566 ( .A(n10272), .B(n3352), .C(n3353), .D(n10436), .Z(n5523) );
  AO4 U5567 ( .A(n10272), .B(n3353), .C(n3354), .D(n10436), .Z(n5524) );
  AO4 U5568 ( .A(n10272), .B(n3354), .C(n3355), .D(n10436), .Z(n5525) );
  AO4 U5569 ( .A(n10272), .B(n3355), .C(n3356), .D(n10436), .Z(n5526) );
  AO4 U5570 ( .A(n10272), .B(n3356), .C(n3357), .D(n10436), .Z(n5527) );
  AO4 U5571 ( .A(n10272), .B(n3357), .C(n3358), .D(n10436), .Z(n5528) );
  AO4 U5572 ( .A(n10272), .B(n3358), .C(n3359), .D(n10436), .Z(n5529) );
  AO4 U5573 ( .A(n10272), .B(n3359), .C(n3360), .D(n10436), .Z(n5530) );
  AO4 U5574 ( .A(n10272), .B(n3360), .C(n3361), .D(n10436), .Z(n5531) );
  AO4 U5575 ( .A(n10272), .B(n3361), .C(n3362), .D(n10436), .Z(n5532) );
  AO4 U5576 ( .A(n10272), .B(n3362), .C(n3363), .D(n10436), .Z(n5533) );
  AO4 U5577 ( .A(n10272), .B(n3363), .C(n3364), .D(n10436), .Z(n5534) );
  AO4 U5578 ( .A(n10271), .B(n3364), .C(n3365), .D(n10436), .Z(n5535) );
  AO4 U5579 ( .A(n10271), .B(n3365), .C(n3366), .D(n10435), .Z(n5536) );
  AO4 U5580 ( .A(n10271), .B(n3366), .C(n3367), .D(n10435), .Z(n5537) );
  AO4 U5581 ( .A(n10271), .B(n3367), .C(n3368), .D(n10435), .Z(n5538) );
  AO4 U5582 ( .A(n10271), .B(n3368), .C(n3369), .D(n10435), .Z(n5539) );
  AO4 U5583 ( .A(n10271), .B(n3369), .C(n3370), .D(n10435), .Z(n5540) );
  AO4 U5584 ( .A(n10271), .B(n3370), .C(n3371), .D(n10435), .Z(n5541) );
  AO4 U5585 ( .A(n10271), .B(n3371), .C(n3372), .D(n10435), .Z(n5542) );
  AO4 U5586 ( .A(n10271), .B(n3372), .C(n3373), .D(n10435), .Z(n5543) );
  AO4 U5587 ( .A(n10271), .B(n3373), .C(n3374), .D(n10435), .Z(n5544) );
  AO4 U5588 ( .A(n10271), .B(n3374), .C(n3375), .D(n10435), .Z(n5545) );
  AO4 U5589 ( .A(n10271), .B(n3375), .C(n3376), .D(n10435), .Z(n5546) );
  AO4 U5590 ( .A(n10271), .B(n3376), .C(n3377), .D(n10435), .Z(n5547) );
  AO4 U5591 ( .A(n10271), .B(n3377), .C(n3378), .D(n10435), .Z(n5548) );
  AO4 U5592 ( .A(n10270), .B(n3378), .C(n3379), .D(n10435), .Z(n5549) );
  AO4 U5593 ( .A(n10270), .B(n3379), .C(n3380), .D(n10434), .Z(n5550) );
  AO4 U5594 ( .A(n10270), .B(n3380), .C(n3381), .D(n10434), .Z(n5551) );
  AO4 U5595 ( .A(n10270), .B(n3381), .C(n3382), .D(n10434), .Z(n5552) );
  AO4 U5596 ( .A(n10270), .B(n3382), .C(n3383), .D(n10434), .Z(n5553) );
  AO4 U5597 ( .A(n10270), .B(n3383), .C(n3384), .D(n10434), .Z(n5554) );
  AO4 U5598 ( .A(n10270), .B(n3384), .C(n3385), .D(n10434), .Z(n5555) );
  AO4 U5599 ( .A(n10270), .B(n3385), .C(n3386), .D(n10434), .Z(n5556) );
  AO4 U5600 ( .A(n10270), .B(n3386), .C(n3387), .D(n10434), .Z(n5557) );
  AO4 U5601 ( .A(n10270), .B(n3387), .C(n3388), .D(n10434), .Z(n5558) );
  AO4 U5602 ( .A(n10270), .B(n3388), .C(n3389), .D(n10434), .Z(n5559) );
  AO4 U5603 ( .A(n10270), .B(n3389), .C(n3390), .D(n10434), .Z(n5560) );
  AO4 U5604 ( .A(n10270), .B(n3390), .C(n3391), .D(n10434), .Z(n5561) );
  AO4 U5605 ( .A(n10270), .B(n3391), .C(n3392), .D(n10434), .Z(n5562) );
  AO4 U5606 ( .A(n10269), .B(n3392), .C(n3393), .D(n10434), .Z(n5563) );
  AO4 U5607 ( .A(n10269), .B(n3393), .C(n3394), .D(n10433), .Z(n5564) );
  AO4 U5608 ( .A(n10269), .B(n3394), .C(n3395), .D(n10433), .Z(n5565) );
  AO4 U5609 ( .A(n10269), .B(n3395), .C(n3396), .D(n10433), .Z(n5566) );
  AO4 U5610 ( .A(n10269), .B(n3396), .C(n3397), .D(n10433), .Z(n5567) );
  AO4 U5611 ( .A(n10269), .B(n3397), .C(n3398), .D(n10433), .Z(n5568) );
  AO4 U5612 ( .A(n10269), .B(n3398), .C(n3399), .D(n10433), .Z(n5569) );
  AO4 U5613 ( .A(n10269), .B(n3399), .C(n3400), .D(n10433), .Z(n5570) );
  AO4 U5614 ( .A(n10269), .B(n3400), .C(n3401), .D(n10433), .Z(n5571) );
  AO4 U5615 ( .A(n10269), .B(n3401), .C(n3402), .D(n10433), .Z(n5572) );
  AO4 U5616 ( .A(n10269), .B(n3402), .C(n3403), .D(n10433), .Z(n5573) );
  AO4 U5617 ( .A(n10269), .B(n3403), .C(n10433), .D(n1418), .Z(n5574) );
  AO4 U5618 ( .A(n10433), .B(n3339), .C(n10269), .D(n1418), .Z(n5866) );
  EN U5619 ( .A(n10251), .B(n10592), .Z(n3405) );
  EN U5620 ( .A(n10244), .B(n10592), .Z(n3406) );
  EN U5621 ( .A(n10241), .B(n10592), .Z(n3407) );
  EN U5622 ( .A(n10238), .B(n10592), .Z(n3408) );
  EN U5623 ( .A(n10235), .B(n10592), .Z(n3409) );
  EN U5624 ( .A(n10232), .B(n10592), .Z(n3410) );
  EN U5625 ( .A(n10229), .B(n10592), .Z(n3411) );
  EN U5626 ( .A(n10226), .B(n10592), .Z(n3412) );
  EN U5627 ( .A(n10223), .B(n10592), .Z(n3413) );
  EN U5628 ( .A(n10220), .B(n10591), .Z(n3414) );
  EN U5629 ( .A(n10217), .B(n10591), .Z(n3415) );
  EN U5630 ( .A(n10214), .B(n10591), .Z(n3416) );
  EN U5631 ( .A(n10211), .B(n10591), .Z(n3417) );
  EN U5632 ( .A(n10208), .B(n10591), .Z(n3418) );
  EN U5633 ( .A(n10205), .B(n10591), .Z(n3419) );
  EN U5634 ( .A(n10202), .B(n10591), .Z(n3420) );
  EN U5635 ( .A(n10199), .B(n10591), .Z(n3421) );
  EN U5636 ( .A(n10196), .B(n10591), .Z(n3422) );
  EN U5637 ( .A(n10193), .B(n10591), .Z(n3423) );
  EN U5638 ( .A(n10190), .B(n10591), .Z(n3424) );
  EN U5639 ( .A(n10187), .B(n10591), .Z(n3425) );
  EN U5640 ( .A(n10184), .B(n10591), .Z(n3426) );
  EN U5641 ( .A(n10181), .B(n10591), .Z(n3427) );
  EN U5642 ( .A(n10178), .B(n10590), .Z(n3428) );
  EN U5643 ( .A(n10175), .B(n10590), .Z(n3429) );
  EN U5644 ( .A(n10172), .B(n10590), .Z(n3430) );
  EN U5645 ( .A(n10169), .B(n10590), .Z(n3431) );
  EN U5646 ( .A(n10166), .B(n10590), .Z(n3432) );
  EN U5647 ( .A(n10163), .B(n10590), .Z(n3433) );
  EN U5648 ( .A(n10160), .B(n10590), .Z(n3434) );
  EN U5649 ( .A(n10157), .B(n10590), .Z(n3435) );
  EN U5650 ( .A(n10154), .B(n10590), .Z(n3436) );
  EN U5651 ( .A(n10151), .B(n10590), .Z(n3437) );
  EN U5652 ( .A(n10148), .B(n10590), .Z(n3438) );
  EN U5653 ( .A(n10145), .B(n10590), .Z(n3439) );
  EN U5654 ( .A(n10142), .B(n10590), .Z(n3440) );
  EN U5655 ( .A(n10139), .B(n10590), .Z(n3441) );
  EN U5656 ( .A(n10136), .B(n10589), .Z(n3442) );
  EN U5657 ( .A(n10133), .B(n10589), .Z(n3443) );
  EN U5658 ( .A(n10130), .B(n10589), .Z(n3444) );
  EN U5659 ( .A(n10127), .B(n10589), .Z(n3445) );
  EN U5660 ( .A(n10124), .B(n10589), .Z(n3446) );
  EN U5661 ( .A(n10121), .B(n10589), .Z(n3447) );
  EN U5662 ( .A(n10118), .B(n10589), .Z(n3448) );
  EN U5663 ( .A(n10115), .B(n10589), .Z(n3449) );
  EN U5664 ( .A(n10112), .B(n10589), .Z(n3450) );
  EN U5665 ( .A(n10109), .B(n10589), .Z(n3451) );
  EN U5666 ( .A(n10106), .B(n10589), .Z(n3452) );
  EN U5667 ( .A(n10103), .B(n10589), .Z(n3453) );
  EN U5668 ( .A(n10100), .B(n10589), .Z(n3454) );
  EN U5669 ( .A(n10097), .B(n10589), .Z(n3455) );
  EN U5670 ( .A(n10094), .B(n10588), .Z(n3456) );
  EN U5671 ( .A(n10091), .B(n10588), .Z(n3457) );
  EN U5672 ( .A(n10088), .B(n10588), .Z(n3458) );
  EN U5673 ( .A(n10085), .B(n10588), .Z(n3459) );
  EN U5674 ( .A(n10082), .B(n10588), .Z(n3460) );
  EN U5675 ( .A(n10079), .B(n10588), .Z(n3461) );
  EN U5676 ( .A(n10076), .B(n10588), .Z(n3462) );
  EN U5677 ( .A(n10073), .B(n10588), .Z(n3463) );
  EN U5678 ( .A(n10070), .B(n10588), .Z(n3464) );
  EN U5679 ( .A(n10067), .B(n10588), .Z(n3465) );
  EN U5680 ( .A(n10064), .B(n10588), .Z(n3466) );
  EN U5681 ( .A(n10061), .B(n10588), .Z(n3467) );
  EN U5682 ( .A(n10058), .B(n10588), .Z(n3468) );
  AO4 U5683 ( .A(n10268), .B(n3405), .C(n3406), .D(n10432), .Z(n5577) );
  AO4 U5684 ( .A(n10268), .B(n3406), .C(n3407), .D(n10432), .Z(n5578) );
  AO4 U5685 ( .A(n10268), .B(n3407), .C(n3408), .D(n10432), .Z(n5579) );
  AO4 U5686 ( .A(n10268), .B(n3408), .C(n3409), .D(n10432), .Z(n5580) );
  AO4 U5687 ( .A(n10268), .B(n3409), .C(n3410), .D(n10432), .Z(n5581) );
  AO4 U5688 ( .A(n10268), .B(n3410), .C(n3411), .D(n10432), .Z(n5582) );
  AO4 U5689 ( .A(n10268), .B(n3411), .C(n3412), .D(n10432), .Z(n5583) );
  AO4 U5690 ( .A(n10268), .B(n3412), .C(n3413), .D(n10432), .Z(n5584) );
  AO4 U5691 ( .A(n10268), .B(n3413), .C(n3414), .D(n10432), .Z(n5585) );
  AO4 U5692 ( .A(n10268), .B(n3414), .C(n3415), .D(n10432), .Z(n5586) );
  AO4 U5693 ( .A(n10267), .B(n3415), .C(n3416), .D(n10432), .Z(n5587) );
  AO4 U5694 ( .A(n10267), .B(n3416), .C(n3417), .D(n10431), .Z(n5588) );
  AO4 U5695 ( .A(n10267), .B(n3417), .C(n3418), .D(n10431), .Z(n5589) );
  AO4 U5696 ( .A(n10267), .B(n3418), .C(n3419), .D(n10431), .Z(n5590) );
  AO4 U5697 ( .A(n10267), .B(n3419), .C(n3420), .D(n10431), .Z(n5591) );
  AO4 U5698 ( .A(n10267), .B(n3420), .C(n3421), .D(n10431), .Z(n5592) );
  AO4 U5699 ( .A(n10267), .B(n3421), .C(n3422), .D(n10431), .Z(n5593) );
  AO4 U5700 ( .A(n10267), .B(n3422), .C(n3423), .D(n10431), .Z(n5594) );
  AO4 U5701 ( .A(n10267), .B(n3423), .C(n3424), .D(n10431), .Z(n5595) );
  AO4 U5702 ( .A(n10267), .B(n3424), .C(n3425), .D(n10431), .Z(n5596) );
  AO4 U5703 ( .A(n10267), .B(n3425), .C(n3426), .D(n10431), .Z(n5597) );
  AO4 U5704 ( .A(n10267), .B(n3426), .C(n3427), .D(n10431), .Z(n5598) );
  AO4 U5705 ( .A(n10267), .B(n3427), .C(n3428), .D(n10431), .Z(n5599) );
  AO4 U5706 ( .A(n10267), .B(n3428), .C(n3429), .D(n10431), .Z(n5600) );
  AO4 U5707 ( .A(n10266), .B(n3429), .C(n3430), .D(n10431), .Z(n5601) );
  AO4 U5708 ( .A(n10266), .B(n3430), .C(n3431), .D(n10430), .Z(n5602) );
  AO4 U5709 ( .A(n10266), .B(n3431), .C(n3432), .D(n10430), .Z(n5603) );
  AO4 U5710 ( .A(n10266), .B(n3432), .C(n3433), .D(n10430), .Z(n5604) );
  AO4 U5711 ( .A(n10266), .B(n3433), .C(n3434), .D(n10430), .Z(n5605) );
  AO4 U5712 ( .A(n10266), .B(n3434), .C(n3435), .D(n10430), .Z(n5606) );
  AO4 U5713 ( .A(n10266), .B(n3435), .C(n3436), .D(n10430), .Z(n5607) );
  AO4 U5714 ( .A(n10266), .B(n3436), .C(n3437), .D(n10430), .Z(n5608) );
  AO4 U5715 ( .A(n10266), .B(n3437), .C(n3438), .D(n10430), .Z(n5609) );
  AO4 U5716 ( .A(n10266), .B(n3438), .C(n3439), .D(n10430), .Z(n5610) );
  AO4 U5717 ( .A(n10266), .B(n3439), .C(n3440), .D(n10430), .Z(n5611) );
  AO4 U5718 ( .A(n10266), .B(n3440), .C(n3441), .D(n10430), .Z(n5612) );
  AO4 U5719 ( .A(n10266), .B(n3441), .C(n3442), .D(n10430), .Z(n5613) );
  AO4 U5720 ( .A(n10266), .B(n3442), .C(n3443), .D(n10430), .Z(n5614) );
  AO4 U5721 ( .A(n10265), .B(n3443), .C(n3444), .D(n10430), .Z(n5615) );
  AO4 U5722 ( .A(n10265), .B(n3444), .C(n3445), .D(n10429), .Z(n5616) );
  AO4 U5723 ( .A(n10265), .B(n3445), .C(n3446), .D(n10429), .Z(n5617) );
  AO4 U5724 ( .A(n10265), .B(n3446), .C(n3447), .D(n10429), .Z(n5618) );
  AO4 U5725 ( .A(n10265), .B(n3447), .C(n3448), .D(n10429), .Z(n5619) );
  AO4 U5726 ( .A(n10265), .B(n3448), .C(n3449), .D(n10429), .Z(n5620) );
  AO4 U5727 ( .A(n10265), .B(n3449), .C(n3450), .D(n10429), .Z(n5621) );
  AO4 U5728 ( .A(n10265), .B(n3450), .C(n3451), .D(n10429), .Z(n5622) );
  AO4 U5729 ( .A(n10265), .B(n3451), .C(n3452), .D(n10429), .Z(n5623) );
  AO4 U5730 ( .A(n10265), .B(n3452), .C(n3453), .D(n10429), .Z(n5624) );
  AO4 U5731 ( .A(n10265), .B(n3453), .C(n3454), .D(n10429), .Z(n5625) );
  AO4 U5732 ( .A(n10265), .B(n3454), .C(n3455), .D(n10429), .Z(n5626) );
  AO4 U5733 ( .A(n10265), .B(n3455), .C(n3456), .D(n10429), .Z(n5627) );
  AO4 U5734 ( .A(n10265), .B(n3456), .C(n3457), .D(n10429), .Z(n5628) );
  AO4 U5735 ( .A(n10264), .B(n3457), .C(n3458), .D(n10429), .Z(n5629) );
  AO4 U5736 ( .A(n10264), .B(n3458), .C(n3459), .D(n10428), .Z(n5630) );
  AO4 U5737 ( .A(n10264), .B(n3459), .C(n3460), .D(n10428), .Z(n5631) );
  AO4 U5738 ( .A(n10264), .B(n3460), .C(n3461), .D(n10428), .Z(n5632) );
  AO4 U5739 ( .A(n10264), .B(n3461), .C(n3462), .D(n10428), .Z(n5633) );
  AO4 U5740 ( .A(n10264), .B(n3462), .C(n3463), .D(n10428), .Z(n5634) );
  AO4 U5741 ( .A(n10264), .B(n3463), .C(n3464), .D(n10428), .Z(n5635) );
  AO4 U5742 ( .A(n10264), .B(n3464), .C(n3465), .D(n10428), .Z(n5636) );
  AO4 U5743 ( .A(n10264), .B(n3465), .C(n3466), .D(n10428), .Z(n5637) );
  AO4 U5744 ( .A(n10264), .B(n3466), .C(n3467), .D(n10428), .Z(n5638) );
  AO4 U5745 ( .A(n10264), .B(n3467), .C(n3468), .D(n10428), .Z(n5639) );
  AO4 U5746 ( .A(n10264), .B(n3468), .C(n10428), .D(n1419), .Z(n5640) );
  AO4 U5747 ( .A(n10428), .B(n3404), .C(n10264), .D(n1419), .Z(n5867) );
  EN U5748 ( .A(n10251), .B(n10587), .Z(n3470) );
  EN U5749 ( .A(n10244), .B(n10587), .Z(n3471) );
  EN U5750 ( .A(n10241), .B(n10587), .Z(n3472) );
  EN U5751 ( .A(n10238), .B(n10587), .Z(n3473) );
  EN U5752 ( .A(n10235), .B(n10587), .Z(n3474) );
  EN U5753 ( .A(n10232), .B(n10587), .Z(n3475) );
  EN U5754 ( .A(n10229), .B(n10587), .Z(n3476) );
  EN U5755 ( .A(n10226), .B(n10587), .Z(n3477) );
  EN U5756 ( .A(n10223), .B(n10587), .Z(n3478) );
  EN U5757 ( .A(n10220), .B(n10586), .Z(n3479) );
  EN U5758 ( .A(n10217), .B(n10586), .Z(n3480) );
  EN U5759 ( .A(n10214), .B(n10586), .Z(n3481) );
  EN U5760 ( .A(n10211), .B(n10586), .Z(n3482) );
  EN U5761 ( .A(n10208), .B(n10586), .Z(n3483) );
  EN U5762 ( .A(n10205), .B(n10586), .Z(n3484) );
  EN U5763 ( .A(n10202), .B(n10586), .Z(n3485) );
  EN U5764 ( .A(n10199), .B(n10586), .Z(n3486) );
  EN U5765 ( .A(n10196), .B(n10586), .Z(n3487) );
  EN U5766 ( .A(n10193), .B(n10586), .Z(n3488) );
  EN U5767 ( .A(n10190), .B(n10586), .Z(n3489) );
  EN U5768 ( .A(n10187), .B(n10586), .Z(n3490) );
  EN U5769 ( .A(n10184), .B(n10586), .Z(n3491) );
  EN U5770 ( .A(n10181), .B(n10586), .Z(n3492) );
  EN U5771 ( .A(n10178), .B(n10585), .Z(n3493) );
  EN U5772 ( .A(n10175), .B(n10585), .Z(n3494) );
  EN U5773 ( .A(n10172), .B(n10585), .Z(n3495) );
  EN U5774 ( .A(n10169), .B(n10585), .Z(n3496) );
  EN U5775 ( .A(n10166), .B(n10585), .Z(n3497) );
  EN U5776 ( .A(n10163), .B(n10585), .Z(n3498) );
  EN U5777 ( .A(n10160), .B(n10585), .Z(n3499) );
  EN U5778 ( .A(n10157), .B(n10585), .Z(n3500) );
  EN U5779 ( .A(n10154), .B(n10585), .Z(n3501) );
  EN U5780 ( .A(n10151), .B(n10585), .Z(n3502) );
  EN U5781 ( .A(n10148), .B(n10585), .Z(n3503) );
  EN U5782 ( .A(n10145), .B(n10585), .Z(n3504) );
  EN U5783 ( .A(n10142), .B(n10585), .Z(n3505) );
  EN U5784 ( .A(n10139), .B(n10585), .Z(n3506) );
  EN U5785 ( .A(n10136), .B(n10584), .Z(n3507) );
  EN U5786 ( .A(n10133), .B(n10584), .Z(n3508) );
  EN U5787 ( .A(n10130), .B(n10584), .Z(n3509) );
  EN U5788 ( .A(n10127), .B(n10584), .Z(n3510) );
  EN U5789 ( .A(n10124), .B(n10584), .Z(n3511) );
  EN U5790 ( .A(n10121), .B(n10584), .Z(n3512) );
  EN U5791 ( .A(n10118), .B(n10584), .Z(n3513) );
  EN U5792 ( .A(n10115), .B(n10584), .Z(n3514) );
  EN U5793 ( .A(n10112), .B(n10584), .Z(n3515) );
  EN U5794 ( .A(n10109), .B(n10584), .Z(n3516) );
  EN U5795 ( .A(n10106), .B(n10584), .Z(n3517) );
  EN U5796 ( .A(n10103), .B(n10584), .Z(n3518) );
  EN U5797 ( .A(n10100), .B(n10584), .Z(n3519) );
  EN U5798 ( .A(n10097), .B(n10584), .Z(n3520) );
  EN U5799 ( .A(n10094), .B(n10583), .Z(n3521) );
  EN U5800 ( .A(n10091), .B(n10583), .Z(n3522) );
  EN U5801 ( .A(n10088), .B(n10583), .Z(n3523) );
  EN U5802 ( .A(n10085), .B(n10583), .Z(n3524) );
  EN U5803 ( .A(n10082), .B(n10583), .Z(n3525) );
  EN U5804 ( .A(n10079), .B(n10583), .Z(n3526) );
  EN U5805 ( .A(n10076), .B(n10583), .Z(n3527) );
  EN U5806 ( .A(n10073), .B(n10583), .Z(n3528) );
  EN U5807 ( .A(n10070), .B(n10583), .Z(n3529) );
  EN U5808 ( .A(n10067), .B(n10583), .Z(n3530) );
  EN U5809 ( .A(n10064), .B(n10583), .Z(n3531) );
  EN U5810 ( .A(n10061), .B(n10583), .Z(n3532) );
  EN U5811 ( .A(n10058), .B(n10583), .Z(n3533) );
  AO4 U5812 ( .A(n10263), .B(n3470), .C(n3471), .D(n10427), .Z(n5643) );
  AO4 U5813 ( .A(n10263), .B(n3471), .C(n3472), .D(n10427), .Z(n5644) );
  AO4 U5814 ( .A(n10263), .B(n3472), .C(n3473), .D(n10427), .Z(n5645) );
  AO4 U5815 ( .A(n10263), .B(n3473), .C(n3474), .D(n10427), .Z(n5646) );
  AO4 U5816 ( .A(n10263), .B(n3474), .C(n3475), .D(n10427), .Z(n5647) );
  AO4 U5817 ( .A(n10263), .B(n3475), .C(n3476), .D(n10427), .Z(n5648) );
  AO4 U5818 ( .A(n10263), .B(n3476), .C(n3477), .D(n10427), .Z(n5649) );
  AO4 U5819 ( .A(n10263), .B(n3477), .C(n3478), .D(n10427), .Z(n5650) );
  AO4 U5820 ( .A(n10263), .B(n3478), .C(n3479), .D(n10427), .Z(n5651) );
  AO4 U5821 ( .A(n10263), .B(n3479), .C(n3480), .D(n10427), .Z(n5652) );
  AO4 U5822 ( .A(n10262), .B(n3480), .C(n3481), .D(n10427), .Z(n5653) );
  AO4 U5823 ( .A(n10262), .B(n3481), .C(n3482), .D(n10426), .Z(n5654) );
  AO4 U5824 ( .A(n10262), .B(n3482), .C(n3483), .D(n10426), .Z(n5655) );
  AO4 U5825 ( .A(n10262), .B(n3483), .C(n3484), .D(n10426), .Z(n5656) );
  AO4 U5826 ( .A(n10262), .B(n3484), .C(n3485), .D(n10426), .Z(n5657) );
  AO4 U5827 ( .A(n10262), .B(n3485), .C(n3486), .D(n10426), .Z(n5658) );
  AO4 U5828 ( .A(n10262), .B(n3486), .C(n3487), .D(n10426), .Z(n5659) );
  AO4 U5829 ( .A(n10262), .B(n3487), .C(n3488), .D(n10426), .Z(n5660) );
  AO4 U5830 ( .A(n10262), .B(n3488), .C(n3489), .D(n10426), .Z(n5661) );
  AO4 U5831 ( .A(n10262), .B(n3489), .C(n3490), .D(n10426), .Z(n5662) );
  AO4 U5832 ( .A(n10262), .B(n3490), .C(n3491), .D(n10426), .Z(n5663) );
  AO4 U5833 ( .A(n10262), .B(n3491), .C(n3492), .D(n10426), .Z(n5664) );
  AO4 U5834 ( .A(n10262), .B(n3492), .C(n3493), .D(n10426), .Z(n5665) );
  AO4 U5835 ( .A(n10262), .B(n3493), .C(n3494), .D(n10426), .Z(n5666) );
  AO4 U5836 ( .A(n10261), .B(n3494), .C(n3495), .D(n10426), .Z(n5667) );
  AO4 U5837 ( .A(n10261), .B(n3495), .C(n3496), .D(n10425), .Z(n5668) );
  AO4 U5838 ( .A(n10261), .B(n3496), .C(n3497), .D(n10425), .Z(n5669) );
  AO4 U5839 ( .A(n10261), .B(n3497), .C(n3498), .D(n10425), .Z(n5670) );
  AO4 U5840 ( .A(n10261), .B(n3498), .C(n3499), .D(n10425), .Z(n5671) );
  AO4 U5841 ( .A(n10261), .B(n3499), .C(n3500), .D(n10425), .Z(n5672) );
  AO4 U5842 ( .A(n10261), .B(n3500), .C(n3501), .D(n10425), .Z(n5673) );
  AO4 U5843 ( .A(n10261), .B(n3501), .C(n3502), .D(n10425), .Z(n5674) );
  AO4 U5844 ( .A(n10261), .B(n3502), .C(n3503), .D(n10425), .Z(n5675) );
  AO4 U5845 ( .A(n10261), .B(n3503), .C(n3504), .D(n10425), .Z(n5676) );
  AO4 U5846 ( .A(n10261), .B(n3504), .C(n3505), .D(n10425), .Z(n5677) );
  AO4 U5847 ( .A(n10261), .B(n3505), .C(n3506), .D(n10425), .Z(n5678) );
  AO4 U5848 ( .A(n10261), .B(n3506), .C(n3507), .D(n10425), .Z(n5679) );
  AO4 U5849 ( .A(n10261), .B(n3507), .C(n3508), .D(n10425), .Z(n5680) );
  AO4 U5850 ( .A(n10260), .B(n3508), .C(n3509), .D(n10425), .Z(n5681) );
  AO4 U5851 ( .A(n10260), .B(n3509), .C(n3510), .D(n10424), .Z(n5682) );
  AO4 U5852 ( .A(n10260), .B(n3510), .C(n3511), .D(n10424), .Z(n5683) );
  AO4 U5853 ( .A(n10260), .B(n3511), .C(n3512), .D(n10424), .Z(n5684) );
  AO4 U5854 ( .A(n10260), .B(n3512), .C(n3513), .D(n10424), .Z(n5685) );
  AO4 U5855 ( .A(n10260), .B(n3513), .C(n3514), .D(n10424), .Z(n5686) );
  AO4 U5856 ( .A(n10260), .B(n3514), .C(n3515), .D(n10424), .Z(n5687) );
  AO4 U5857 ( .A(n10260), .B(n3515), .C(n3516), .D(n10424), .Z(n5688) );
  AO4 U5858 ( .A(n10260), .B(n3516), .C(n3517), .D(n10424), .Z(n5689) );
  AO4 U5859 ( .A(n10260), .B(n3517), .C(n3518), .D(n10424), .Z(n5690) );
  AO4 U5860 ( .A(n10260), .B(n3518), .C(n3519), .D(n10424), .Z(n5691) );
  AO4 U5861 ( .A(n10260), .B(n3519), .C(n3520), .D(n10424), .Z(n5692) );
  AO4 U5862 ( .A(n10260), .B(n3520), .C(n3521), .D(n10424), .Z(n5693) );
  AO4 U5863 ( .A(n10260), .B(n3521), .C(n3522), .D(n10424), .Z(n5694) );
  AO4 U5864 ( .A(n10259), .B(n3522), .C(n3523), .D(n10424), .Z(n5695) );
  AO4 U5865 ( .A(n10259), .B(n3523), .C(n3524), .D(n10423), .Z(n5696) );
  AO4 U5866 ( .A(n10259), .B(n3524), .C(n3525), .D(n10423), .Z(n5697) );
  AO4 U5867 ( .A(n10259), .B(n3525), .C(n3526), .D(n10423), .Z(n5698) );
  AO4 U5868 ( .A(n10259), .B(n3526), .C(n3527), .D(n10423), .Z(n5699) );
  AO4 U5869 ( .A(n10259), .B(n3527), .C(n3528), .D(n10423), .Z(n5700) );
  AO4 U5870 ( .A(n10259), .B(n3528), .C(n3529), .D(n10423), .Z(n5701) );
  AO4 U5871 ( .A(n10259), .B(n3529), .C(n3530), .D(n10423), .Z(n5702) );
  AO4 U5872 ( .A(n10259), .B(n3530), .C(n3531), .D(n10423), .Z(n5703) );
  AO4 U5873 ( .A(n10259), .B(n3531), .C(n3532), .D(n10423), .Z(n5704) );
  AO4 U5874 ( .A(n10259), .B(n3532), .C(n3533), .D(n10423), .Z(n5705) );
  AO4 U5875 ( .A(n10259), .B(n3533), .C(n10423), .D(n1420), .Z(n5706) );
  AO4 U5876 ( .A(n10423), .B(n3469), .C(n10259), .D(n1420), .Z(n5868) );
  EN U5877 ( .A(n10251), .B(n10582), .Z(n3535) );
  EN U5878 ( .A(n10244), .B(n10582), .Z(n3536) );
  EN U5879 ( .A(n10241), .B(n10582), .Z(n3537) );
  EN U5880 ( .A(n10238), .B(n10582), .Z(n3538) );
  EN U5881 ( .A(n10235), .B(n10582), .Z(n3539) );
  EN U5882 ( .A(n10232), .B(n10582), .Z(n3540) );
  EN U5883 ( .A(n10229), .B(n10582), .Z(n3541) );
  EN U5884 ( .A(n10226), .B(n10582), .Z(n3542) );
  EN U5885 ( .A(n10223), .B(n10582), .Z(n3543) );
  EN U5886 ( .A(n10220), .B(n10581), .Z(n3544) );
  EN U5887 ( .A(n10217), .B(n10581), .Z(n3545) );
  EN U5888 ( .A(n10214), .B(n10581), .Z(n3546) );
  EN U5889 ( .A(n10211), .B(n10581), .Z(n3547) );
  EN U5890 ( .A(n10208), .B(n10581), .Z(n3548) );
  EN U5891 ( .A(n10205), .B(n10581), .Z(n3549) );
  EN U5892 ( .A(n10202), .B(n10581), .Z(n3550) );
  EN U5893 ( .A(n10199), .B(n10581), .Z(n3551) );
  EN U5894 ( .A(n10196), .B(n10581), .Z(n3552) );
  EN U5895 ( .A(n10193), .B(n10581), .Z(n3553) );
  EN U5896 ( .A(n10190), .B(n10581), .Z(n3554) );
  EN U5897 ( .A(n10187), .B(n10581), .Z(n3555) );
  EN U5898 ( .A(n10184), .B(n10581), .Z(n3556) );
  EN U5899 ( .A(n10181), .B(n10581), .Z(n3557) );
  EN U5900 ( .A(n10178), .B(n10580), .Z(n3558) );
  EN U5901 ( .A(n10175), .B(n10580), .Z(n3559) );
  EN U5902 ( .A(n10172), .B(n10580), .Z(n3560) );
  EN U5903 ( .A(n10169), .B(n10580), .Z(n3561) );
  EN U5904 ( .A(n10166), .B(n10580), .Z(n3562) );
  EN U5905 ( .A(n10163), .B(n10580), .Z(n3563) );
  EN U5906 ( .A(n10160), .B(n10580), .Z(n3564) );
  EN U5907 ( .A(n10157), .B(n10580), .Z(n3565) );
  EN U5908 ( .A(n10154), .B(n10580), .Z(n3566) );
  EN U5909 ( .A(n10151), .B(n10580), .Z(n3567) );
  EN U5910 ( .A(n10148), .B(n10580), .Z(n3568) );
  EN U5911 ( .A(n10145), .B(n10580), .Z(n3569) );
  EN U5912 ( .A(n10142), .B(n10580), .Z(n3570) );
  EN U5913 ( .A(n10139), .B(n10580), .Z(n3571) );
  EN U5914 ( .A(n10136), .B(n10579), .Z(n3572) );
  EN U5915 ( .A(n10133), .B(n10579), .Z(n3573) );
  EN U5916 ( .A(n10130), .B(n10579), .Z(n3574) );
  EN U5917 ( .A(n10127), .B(n10579), .Z(n3575) );
  EN U5918 ( .A(n10124), .B(n10579), .Z(n3576) );
  EN U5919 ( .A(n10121), .B(n10579), .Z(n3577) );
  EN U5920 ( .A(n10118), .B(n10579), .Z(n3578) );
  EN U5921 ( .A(n10115), .B(n10579), .Z(n3579) );
  EN U5922 ( .A(n10112), .B(n10579), .Z(n3580) );
  EN U5923 ( .A(n10109), .B(n10579), .Z(n3581) );
  EN U5924 ( .A(n10106), .B(n10579), .Z(n3582) );
  EN U5925 ( .A(n10103), .B(n10579), .Z(n3583) );
  EN U5926 ( .A(n10100), .B(n10579), .Z(n3584) );
  EN U5927 ( .A(n10097), .B(n10579), .Z(n3585) );
  EN U5928 ( .A(n10094), .B(n10578), .Z(n3586) );
  EN U5929 ( .A(n10091), .B(n10578), .Z(n3587) );
  EN U5930 ( .A(n10088), .B(n10578), .Z(n3588) );
  EN U5931 ( .A(n10085), .B(n10578), .Z(n3589) );
  EN U5932 ( .A(n10082), .B(n10578), .Z(n3590) );
  EN U5933 ( .A(n10079), .B(n10578), .Z(n3591) );
  EN U5934 ( .A(n10076), .B(n10578), .Z(n3592) );
  EN U5935 ( .A(n10073), .B(n10578), .Z(n3593) );
  EN U5936 ( .A(n10070), .B(n10578), .Z(n3594) );
  EN U5937 ( .A(n10067), .B(n10578), .Z(n3595) );
  EN U5938 ( .A(n10064), .B(n10578), .Z(n3596) );
  EN U5939 ( .A(n10061), .B(n10578), .Z(n3597) );
  EN U5940 ( .A(n10058), .B(n10578), .Z(n3598) );
  AO4 U5941 ( .A(n10258), .B(n3535), .C(n3536), .D(n10422), .Z(n5709) );
  AO4 U5942 ( .A(n10258), .B(n3536), .C(n3537), .D(n10422), .Z(n5710) );
  AO4 U5943 ( .A(n10258), .B(n3537), .C(n3538), .D(n10422), .Z(n5711) );
  AO4 U5944 ( .A(n10258), .B(n3538), .C(n3539), .D(n10422), .Z(n5712) );
  AO4 U5945 ( .A(n10258), .B(n3539), .C(n3540), .D(n10422), .Z(n5713) );
  AO4 U5946 ( .A(n10258), .B(n3540), .C(n3541), .D(n10422), .Z(n5714) );
  AO4 U5947 ( .A(n10258), .B(n3541), .C(n3542), .D(n10422), .Z(n5715) );
  AO4 U5948 ( .A(n10258), .B(n3542), .C(n3543), .D(n10422), .Z(n5716) );
  AO4 U5949 ( .A(n10258), .B(n3543), .C(n3544), .D(n10422), .Z(n5717) );
  AO4 U5950 ( .A(n10258), .B(n3544), .C(n3545), .D(n10422), .Z(n5718) );
  AO4 U5951 ( .A(n10257), .B(n3545), .C(n3546), .D(n10422), .Z(n5719) );
  AO4 U5952 ( .A(n10257), .B(n3546), .C(n3547), .D(n10421), .Z(n5720) );
  AO4 U5953 ( .A(n10257), .B(n3547), .C(n3548), .D(n10421), .Z(n5721) );
  AO4 U5954 ( .A(n10257), .B(n3548), .C(n3549), .D(n10421), .Z(n5722) );
  AO4 U5955 ( .A(n10257), .B(n3549), .C(n3550), .D(n10421), .Z(n5723) );
  AO4 U5956 ( .A(n10257), .B(n3550), .C(n3551), .D(n10421), .Z(n5724) );
  AO4 U5957 ( .A(n10257), .B(n3551), .C(n3552), .D(n10421), .Z(n5725) );
  AO4 U5958 ( .A(n10257), .B(n3552), .C(n3553), .D(n10421), .Z(n5726) );
  AO4 U5959 ( .A(n10257), .B(n3553), .C(n3554), .D(n10421), .Z(n5727) );
  AO4 U5960 ( .A(n10257), .B(n3554), .C(n3555), .D(n10421), .Z(n5728) );
  AO4 U5961 ( .A(n10257), .B(n3555), .C(n3556), .D(n10421), .Z(n5729) );
  AO4 U5962 ( .A(n10257), .B(n3556), .C(n3557), .D(n10421), .Z(n5730) );
  AO4 U5963 ( .A(n10257), .B(n3557), .C(n3558), .D(n10421), .Z(n5731) );
  AO4 U5964 ( .A(n10257), .B(n3558), .C(n3559), .D(n10421), .Z(n5732) );
  AO4 U5965 ( .A(n10256), .B(n3559), .C(n3560), .D(n10421), .Z(n5733) );
  AO4 U5966 ( .A(n10256), .B(n3560), .C(n3561), .D(n10420), .Z(n5734) );
  AO4 U5967 ( .A(n10256), .B(n3561), .C(n3562), .D(n10420), .Z(n5735) );
  AO4 U5968 ( .A(n10256), .B(n3562), .C(n3563), .D(n10420), .Z(n5736) );
  AO4 U5969 ( .A(n10256), .B(n3563), .C(n3564), .D(n10420), .Z(n5737) );
  AO4 U5970 ( .A(n10256), .B(n3564), .C(n3565), .D(n10420), .Z(n5738) );
  AO4 U5971 ( .A(n10256), .B(n3565), .C(n3566), .D(n10420), .Z(n5739) );
  AO4 U5972 ( .A(n10256), .B(n3566), .C(n3567), .D(n10420), .Z(n5740) );
  AO4 U5973 ( .A(n10256), .B(n3567), .C(n3568), .D(n10420), .Z(n5741) );
  AO4 U5974 ( .A(n10256), .B(n3568), .C(n3569), .D(n10420), .Z(n5742) );
  AO4 U5975 ( .A(n10256), .B(n3569), .C(n3570), .D(n10420), .Z(n5743) );
  AO4 U5976 ( .A(n10256), .B(n3570), .C(n3571), .D(n10420), .Z(n5744) );
  AO4 U5977 ( .A(n10256), .B(n3571), .C(n3572), .D(n10420), .Z(n5745) );
  AO4 U5978 ( .A(n10256), .B(n3572), .C(n3573), .D(n10420), .Z(n5746) );
  AO4 U5979 ( .A(n10255), .B(n3573), .C(n3574), .D(n10420), .Z(n5747) );
  AO4 U5980 ( .A(n10255), .B(n3574), .C(n3575), .D(n10419), .Z(n5748) );
  AO4 U5981 ( .A(n10255), .B(n3575), .C(n3576), .D(n10419), .Z(n5749) );
  AO4 U5982 ( .A(n10255), .B(n3576), .C(n3577), .D(n10419), .Z(n5750) );
  AO4 U5983 ( .A(n10255), .B(n3577), .C(n3578), .D(n10419), .Z(n5751) );
  AO4 U5984 ( .A(n10255), .B(n3578), .C(n3579), .D(n10419), .Z(n5752) );
  AO4 U5985 ( .A(n10255), .B(n3579), .C(n3580), .D(n10419), .Z(n5753) );
  AO4 U5986 ( .A(n10255), .B(n3580), .C(n3581), .D(n10419), .Z(n5754) );
  AO4 U5987 ( .A(n10255), .B(n3581), .C(n3582), .D(n10419), .Z(n5755) );
  AO4 U5988 ( .A(n10255), .B(n3582), .C(n3583), .D(n10419), .Z(n5756) );
  AO4 U5989 ( .A(n10255), .B(n3583), .C(n3584), .D(n10419), .Z(n5757) );
  AO4 U5990 ( .A(n10255), .B(n3584), .C(n3585), .D(n10419), .Z(n5758) );
  AO4 U5991 ( .A(n10255), .B(n3585), .C(n3586), .D(n10419), .Z(n5759) );
  AO4 U5992 ( .A(n10255), .B(n3586), .C(n3587), .D(n10419), .Z(n5760) );
  AO4 U5993 ( .A(n10254), .B(n3587), .C(n3588), .D(n10419), .Z(n5761) );
  AO4 U5994 ( .A(n10254), .B(n3588), .C(n3589), .D(n10418), .Z(n5762) );
  AO4 U5995 ( .A(n10254), .B(n3589), .C(n3590), .D(n10418), .Z(n5763) );
  AO4 U5996 ( .A(n10254), .B(n3590), .C(n3591), .D(n10418), .Z(n5764) );
  AO4 U5997 ( .A(n10254), .B(n3591), .C(n3592), .D(n10418), .Z(n5765) );
  AO4 U5998 ( .A(n10254), .B(n3592), .C(n3593), .D(n10418), .Z(n5766) );
  AO4 U5999 ( .A(n10254), .B(n3593), .C(n3594), .D(n10418), .Z(n5767) );
  AO4 U6000 ( .A(n10254), .B(n3594), .C(n3595), .D(n10418), .Z(n5768) );
  AO4 U6001 ( .A(n10254), .B(n3595), .C(n3596), .D(n10418), .Z(n5769) );
  AO4 U6002 ( .A(n10254), .B(n3596), .C(n3597), .D(n10418), .Z(n5770) );
  AO4 U6003 ( .A(n10254), .B(n3597), .C(n3598), .D(n10418), .Z(n5771) );
  AO4 U6004 ( .A(n10254), .B(n3598), .C(n10418), .D(n1421), .Z(n5772) );
  AO4 U6005 ( .A(n10418), .B(n3534), .C(n10254), .D(n1421), .Z(n5869) );
  IVP U6006 ( .A(n10244), .Z(n3599) );
  IVP U6007 ( .A(n10241), .Z(n3600) );
  IVP U6008 ( .A(n10238), .Z(n3601) );
  IVP U6009 ( .A(n10235), .Z(n3602) );
  IVP U6010 ( .A(n10232), .Z(n3603) );
  IVP U6011 ( .A(n10229), .Z(n3604) );
  IVP U6012 ( .A(n10226), .Z(n3605) );
  IVP U6013 ( .A(n10223), .Z(n3606) );
  IVP U6014 ( .A(n10220), .Z(n3607) );
  IVP U6015 ( .A(n10217), .Z(n3608) );
  IVP U6016 ( .A(n10214), .Z(n3609) );
  IVP U6017 ( .A(n10211), .Z(n3610) );
  IVP U6018 ( .A(n10208), .Z(n3611) );
  IVP U6019 ( .A(n10205), .Z(n3612) );
  IVP U6020 ( .A(n10202), .Z(n3613) );
  IVP U6021 ( .A(n10199), .Z(n3614) );
  IVP U6022 ( .A(n10196), .Z(n3615) );
  IVP U6023 ( .A(n10193), .Z(n3616) );
  IVP U6024 ( .A(n10190), .Z(n3617) );
  IVP U6025 ( .A(n10187), .Z(n3618) );
  IVP U6026 ( .A(n10184), .Z(n3619) );
  IVP U6027 ( .A(n10181), .Z(n3620) );
  IVP U6028 ( .A(n10178), .Z(n3621) );
  IVP U6029 ( .A(n10175), .Z(n3622) );
  IVP U6030 ( .A(n10172), .Z(n3623) );
  IVP U6031 ( .A(n10169), .Z(n3624) );
  IVP U6032 ( .A(n10166), .Z(n3625) );
  IVP U6033 ( .A(n10163), .Z(n3626) );
  IVP U6034 ( .A(n10160), .Z(n3627) );
  IVP U6035 ( .A(n10157), .Z(n3628) );
  IVP U6036 ( .A(n10154), .Z(n3629) );
  IVP U6037 ( .A(n10151), .Z(n3630) );
  IVP U6038 ( .A(n10148), .Z(n3631) );
  IVP U6039 ( .A(n10145), .Z(n3632) );
  IVP U6040 ( .A(n10142), .Z(n3633) );
  IVP U6041 ( .A(n10139), .Z(n3634) );
  IVP U6042 ( .A(n10136), .Z(n3635) );
  IVP U6043 ( .A(n10133), .Z(n3636) );
  IVP U6044 ( .A(n10130), .Z(n3637) );
  IVP U6045 ( .A(n10127), .Z(n3638) );
  IVP U6046 ( .A(n10124), .Z(n3639) );
  IVP U6047 ( .A(n10121), .Z(n3640) );
  IVP U6048 ( .A(n10118), .Z(n3641) );
  IVP U6049 ( .A(n10115), .Z(n3642) );
  IVP U6050 ( .A(n10112), .Z(n3643) );
  IVP U6051 ( .A(n10109), .Z(n3644) );
  IVP U6052 ( .A(n10106), .Z(n3645) );
  IVP U6053 ( .A(n10103), .Z(n3646) );
  IVP U6054 ( .A(n10100), .Z(n3647) );
  IVP U6055 ( .A(n10097), .Z(n3648) );
  IVP U6056 ( .A(n10094), .Z(n3649) );
  IVP U6057 ( .A(n10091), .Z(n3650) );
  IVP U6058 ( .A(n10088), .Z(n3651) );
  IVP U6059 ( .A(n10085), .Z(n3652) );
  IVP U6060 ( .A(n10082), .Z(n3653) );
  IVP U6061 ( .A(n10079), .Z(n3654) );
  IVP U6062 ( .A(n10076), .Z(n3655) );
  IVP U6063 ( .A(n10073), .Z(n3656) );
  IVP U6064 ( .A(n10070), .Z(n3657) );
  IVP U6065 ( .A(n10067), .Z(n3658) );
  IVP U6066 ( .A(n10064), .Z(n3659) );
  IVP U6067 ( .A(n10061), .Z(n3660) );
  IVP U6068 ( .A(n10058), .Z(n3661) );
  NR2 U6069 ( .A(n3599), .B(n10417), .Z(n5775) );
  NR2 U6070 ( .A(n3600), .B(n10417), .Z(n5776) );
  NR2 U6071 ( .A(n3601), .B(n10417), .Z(n5777) );
  NR2 U6072 ( .A(n3602), .B(n10417), .Z(n5778) );
  NR2 U6073 ( .A(n3603), .B(n10417), .Z(n5779) );
  NR2 U6074 ( .A(n3604), .B(n10417), .Z(n5780) );
  NR2 U6075 ( .A(n3605), .B(n10417), .Z(n5781) );
  NR2 U6076 ( .A(n3606), .B(n10417), .Z(n5782) );
  NR2 U6077 ( .A(n3607), .B(n10417), .Z(n5783) );
  NR2 U6078 ( .A(n3608), .B(n10417), .Z(n5784) );
  NR2 U6079 ( .A(n3609), .B(n10417), .Z(n5785) );
  NR2 U6080 ( .A(n3610), .B(n10417), .Z(n5786) );
  NR2 U6081 ( .A(n3611), .B(n10417), .Z(n5787) );
  NR2 U6082 ( .A(n3612), .B(n10417), .Z(n5788) );
  NR2 U6083 ( .A(n3613), .B(n10417), .Z(n5789) );
  NR2 U6084 ( .A(n3614), .B(n10417), .Z(n5790) );
  NR2 U6085 ( .A(n3615), .B(n10416), .Z(n5791) );
  NR2 U6086 ( .A(n3616), .B(n10416), .Z(n5792) );
  NR2 U6087 ( .A(n3617), .B(n10416), .Z(n5793) );
  NR2 U6088 ( .A(n3618), .B(n10416), .Z(n5794) );
  NR2 U6089 ( .A(n3619), .B(n10416), .Z(n5795) );
  NR2 U6090 ( .A(n3620), .B(n10416), .Z(n5796) );
  NR2 U6091 ( .A(n3621), .B(n10416), .Z(n5797) );
  NR2 U6092 ( .A(n3622), .B(n10416), .Z(n5798) );
  NR2 U6093 ( .A(n3623), .B(n10416), .Z(n5799) );
  NR2 U6094 ( .A(n3624), .B(n10416), .Z(n5800) );
  NR2 U6095 ( .A(n3625), .B(n10416), .Z(n5801) );
  NR2 U6096 ( .A(n3626), .B(n10416), .Z(n5802) );
  NR2 U6097 ( .A(n3627), .B(n10416), .Z(n5803) );
  NR2 U6098 ( .A(n3628), .B(n10416), .Z(n5804) );
  NR2 U6099 ( .A(n3629), .B(n10416), .Z(n5805) );
  NR2 U6100 ( .A(n3630), .B(n10416), .Z(n5806) );
  NR2 U6101 ( .A(n3631), .B(n10415), .Z(n5807) );
  NR2 U6102 ( .A(n3632), .B(n10415), .Z(n5808) );
  NR2 U6103 ( .A(n3633), .B(n10415), .Z(n5809) );
  NR2 U6104 ( .A(n3634), .B(n10415), .Z(n5810) );
  NR2 U6105 ( .A(n3635), .B(n10415), .Z(n5811) );
  NR2 U6106 ( .A(n3636), .B(n10415), .Z(n5812) );
  NR2 U6107 ( .A(n3637), .B(n10415), .Z(n5813) );
  NR2 U6108 ( .A(n3638), .B(n10415), .Z(n5814) );
  NR2 U6109 ( .A(n3639), .B(n10415), .Z(n5815) );
  NR2 U6110 ( .A(n3640), .B(n10415), .Z(n5816) );
  NR2 U6111 ( .A(n3641), .B(n10415), .Z(n5817) );
  NR2 U6112 ( .A(n3642), .B(n10415), .Z(n5818) );
  NR2 U6113 ( .A(n3643), .B(n10415), .Z(n5819) );
  NR2 U6114 ( .A(n3644), .B(n10415), .Z(n5820) );
  NR2 U6115 ( .A(n3645), .B(n10415), .Z(n5821) );
  NR2 U6116 ( .A(n3646), .B(n10415), .Z(n5822) );
  NR2 U6117 ( .A(n3647), .B(n10414), .Z(n5823) );
  NR2 U6118 ( .A(n3648), .B(n10414), .Z(n5824) );
  NR2 U6119 ( .A(n3649), .B(n10414), .Z(n5825) );
  NR2 U6120 ( .A(n3650), .B(n10414), .Z(n5826) );
  NR2 U6121 ( .A(n3651), .B(n10414), .Z(n5827) );
  NR2 U6122 ( .A(n3652), .B(n10414), .Z(n5828) );
  NR2 U6123 ( .A(n3653), .B(n10414), .Z(n5829) );
  NR2 U6124 ( .A(n3654), .B(n10414), .Z(n5830) );
  NR2 U6125 ( .A(n3655), .B(n10414), .Z(n5831) );
  NR2 U6126 ( .A(n3656), .B(n10414), .Z(n5832) );
  NR2 U6127 ( .A(n3657), .B(n10414), .Z(n5833) );
  NR2 U6128 ( .A(n3658), .B(n10414), .Z(n5834) );
  NR2 U6129 ( .A(n3659), .B(n10414), .Z(n5835) );
  NR2 U6130 ( .A(n3660), .B(n10414), .Z(n5836) );
  NR2 U6131 ( .A(n3661), .B(n10414), .Z(n5837) );
  HA1 U6132 ( .A(n3729), .B(n3665), .S(n5870), .CO(n5871) );
  FA1A U6133 ( .CI(n3730), .A(n3666), .B(n10897), .S(n5872), .CO(n5873) );
  HA1 U6134 ( .A(n5840), .B(n3795), .S(n5874), .CO(n5875) );
  FA1A U6135 ( .CI(n5874), .A(n3731), .B(n3667), .S(n5876), .CO(n5877) );
  FA1A U6136 ( .CI(n3796), .A(n3668), .B(n10896), .S(n5878), .CO(n5879) );
  FA1A U6137 ( .CI(n5878), .A(n5875), .B(n3732), .S(n5880), .CO(n5881) );
  HA1 U6138 ( .A(n5841), .B(n3861), .S(n5882), .CO(n5883) );
  FA1A U6139 ( .CI(n3733), .A(n3797), .B(n3669), .S(n5884), .CO(n5885) );
  FA1A U6140 ( .CI(n5884), .A(n5879), .B(n5882), .S(n5886), .CO(n5887) );
  FA1A U6141 ( .CI(n3862), .A(n3798), .B(n10895), .S(n5888), .CO(n5889) );
  FA1A U6142 ( .CI(n5883), .A(n3734), .B(n3670), .S(n5890), .CO(n5891) );
  FA1A U6143 ( .CI(n5890), .A(n5885), .B(n5888), .S(n5892), .CO(n5893) );
  HA1 U6144 ( .A(n5842), .B(n3927), .S(n5894), .CO(n5895) );
  FA1A U6145 ( .CI(n3735), .A(n3863), .B(n3799), .S(n5896), .CO(n5897) );
  FA1A U6146 ( .CI(n5889), .A(n5894), .B(n3671), .S(n5898), .CO(n5899) );
  FA1A U6147 ( .CI(n5898), .A(n5896), .B(n5891), .S(n5900), .CO(n5901) );
  FA1A U6148 ( .CI(n3928), .A(n3864), .B(n10894), .S(n5902), .CO(n5903) );
  FA1A U6149 ( .CI(n5895), .A(n3736), .B(n3800), .S(n5904), .CO(n5905) );
  FA1A U6150 ( .CI(n5897), .A(n5902), .B(n3672), .S(n5906), .CO(n5907) );
  FA1A U6151 ( .CI(n5906), .A(n5899), .B(n5904), .S(n5908), .CO(n5909) );
  HA1 U6152 ( .A(n5843), .B(n3993), .S(n5910), .CO(n5911) );
  FA1A U6153 ( .CI(n3673), .A(n3929), .B(n3801), .S(n5912), .CO(n5913) );
  FA1A U6154 ( .CI(n5910), .A(n3865), .B(n3737), .S(n5914), .CO(n5915) );
  FA1A U6155 ( .CI(n5914), .A(n5912), .B(n5903), .S(n5916), .CO(n5917) );
  FA1A U6156 ( .CI(n5916), .A(n5907), .B(n5905), .S(n5918), .CO(n5919) );
  FA1A U6157 ( .CI(n3994), .A(n3930), .B(n10893), .S(n5920), .CO(n5921) );
  FA1A U6158 ( .CI(n5911), .A(n3674), .B(n3802), .S(n5922), .CO(n5923) );
  FA1A U6159 ( .CI(n5920), .A(n3866), .B(n3738), .S(n5924), .CO(n5925) );
  FA1A U6160 ( .CI(n5924), .A(n5922), .B(n5913), .S(n5926), .CO(n5927) );
  FA1A U6161 ( .CI(n5926), .A(n5917), .B(n5915), .S(n5928), .CO(n5929) );
  HA1 U6162 ( .A(n5844), .B(n4059), .S(n5930), .CO(n5931) );
  FA1A U6163 ( .CI(n3739), .A(n3675), .B(n3867), .S(n5932), .CO(n5933) );
  FA1A U6164 ( .CI(n3931), .A(n3995), .B(n3803), .S(n5934), .CO(n5935) );
  FA1A U6165 ( .CI(n5934), .A(n5921), .B(n5930), .S(n5936), .CO(n5937) );
  FA1A U6166 ( .CI(n5925), .A(n5932), .B(n5923), .S(n5938), .CO(n5939) );
  FA1A U6167 ( .CI(n5938), .A(n5927), .B(n5936), .S(n5940), .CO(n5941) );
  FA1A U6168 ( .CI(n4060), .A(n3996), .B(n10892), .S(n5942), .CO(n5943) );
  FA1A U6169 ( .CI(n5931), .A(n3932), .B(n3868), .S(n5944), .CO(n5945) );
  FA1A U6170 ( .CI(n3740), .A(n3804), .B(n3676), .S(n5946), .CO(n5947) );
  FA1A U6171 ( .CI(n5946), .A(n5935), .B(n5942), .S(n5948), .CO(n5949) );
  FA1A U6172 ( .CI(n5937), .A(n5944), .B(n5933), .S(n5950), .CO(n5951) );
  FA1A U6173 ( .CI(n5950), .A(n5939), .B(n5948), .S(n5952), .CO(n5953) );
  HA1 U6174 ( .A(n5845), .B(n4125), .S(n5954), .CO(n5955) );
  FA1A U6175 ( .CI(n3677), .A(n4061), .B(n3869), .S(n5956), .CO(n5957) );
  FA1A U6176 ( .CI(n3997), .A(n3741), .B(n3933), .S(n5958), .CO(n5959) );
  FA1A U6177 ( .CI(n5943), .A(n5954), .B(n3805), .S(n5960), .CO(n5961) );
  FA1A U6178 ( .CI(n5958), .A(n5956), .B(n5945), .S(n5962), .CO(n5963) );
  FA1A U6179 ( .CI(n5949), .A(n5960), .B(n5947), .S(n5964), .CO(n5965) );
  FA1A U6180 ( .CI(n5964), .A(n5951), .B(n5962), .S(n5966), .CO(n5967) );
  FA1A U6181 ( .CI(n4126), .A(n4062), .B(n10891), .S(n5968), .CO(n5969) );
  FA1A U6182 ( .CI(n5955), .A(n3678), .B(n3870), .S(n5970), .CO(n5971) );
  FA1A U6183 ( .CI(n3934), .A(n3998), .B(n3742), .S(n5972), .CO(n5973) );
  FA1A U6184 ( .CI(n5957), .A(n5968), .B(n3806), .S(n5974), .CO(n5975) );
  FA1A U6185 ( .CI(n5972), .A(n5970), .B(n5959), .S(n5976), .CO(n5977) );
  FA1A U6186 ( .CI(n5976), .A(n5974), .B(n5961), .S(n5978), .CO(n5979) );
  FA1A U6187 ( .CI(n5978), .A(n5965), .B(n5963), .S(n5980), .CO(n5981) );
  HA1 U6188 ( .A(n5846), .B(n4191), .S(n5982), .CO(n5983) );
  FA1A U6189 ( .CI(n3743), .A(n3679), .B(n3935), .S(n5984), .CO(n5985) );
  FA1A U6190 ( .CI(n3999), .A(n4127), .B(n4063), .S(n5986), .CO(n5987) );
  FA1A U6191 ( .CI(n5982), .A(n3871), .B(n3807), .S(n5988), .CO(n5989) );
  FA1A U6192 ( .CI(n5988), .A(n5986), .B(n5969), .S(n5990), .CO(n5991) );
  FA1A U6193 ( .CI(n5984), .A(n5973), .B(n5971), .S(n5992), .CO(n5993) );
  FA1A U6194 ( .CI(n5992), .A(n5990), .B(n5975), .S(n5994), .CO(n5995) );
  FA1A U6195 ( .CI(n5994), .A(n5979), .B(n5977), .S(n5996), .CO(n5997) );
  FA1A U6196 ( .CI(n4192), .A(n4128), .B(n10890), .S(n5998), .CO(n5999) );
  FA1A U6197 ( .CI(n5983), .A(n3680), .B(n3936), .S(n6000), .CO(n6001) );
  FA1A U6198 ( .CI(n4000), .A(n4064), .B(n3744), .S(n6002), .CO(n6003) );
  FA1A U6199 ( .CI(n5998), .A(n3872), .B(n3808), .S(n6004), .CO(n6005) );
  FA1A U6200 ( .CI(n6004), .A(n6000), .B(n5985), .S(n6006), .CO(n6007) );
  FA1A U6201 ( .CI(n5989), .A(n6002), .B(n5987), .S(n6008), .CO(n6009) );
  FA1A U6202 ( .CI(n6006), .A(n6008), .B(n5991), .S(n6010), .CO(n6011) );
  FA1A U6203 ( .CI(n6010), .A(n5995), .B(n5993), .S(n6012), .CO(n6013) );
  HA1 U6204 ( .A(n5847), .B(n4257), .S(n6014), .CO(n6015) );
  FA1A U6205 ( .CI(n4129), .A(n4193), .B(n3937), .S(n6016), .CO(n6017) );
  FA1A U6206 ( .CI(n4065), .A(n3681), .B(n3873), .S(n6018), .CO(n6019) );
  FA1A U6207 ( .CI(n3809), .A(n4001), .B(n3745), .S(n6020), .CO(n6021) );
  FA1A U6208 ( .CI(n6020), .A(n5999), .B(n6014), .S(n6022), .CO(n6023) );
  FA1A U6209 ( .CI(n6005), .A(n6016), .B(n6001), .S(n6024), .CO(n6025) );
  FA1A U6210 ( .CI(n6022), .A(n6018), .B(n6003), .S(n6026), .CO(n6027) );
  FA1A U6211 ( .CI(n6026), .A(n6024), .B(n6007), .S(n6028), .CO(n6029) );
  FA1A U6212 ( .CI(n6028), .A(n6011), .B(n6009), .S(n6030), .CO(n6031) );
  FA1A U6213 ( .CI(n4258), .A(n4194), .B(n10889), .S(n6032), .CO(n6033) );
  FA1A U6214 ( .CI(n6015), .A(n4130), .B(n3938), .S(n6034), .CO(n6035) );
  FA1A U6215 ( .CI(n4066), .A(n3682), .B(n3874), .S(n6036), .CO(n6037) );
  FA1A U6216 ( .CI(n3810), .A(n4002), .B(n3746), .S(n6038), .CO(n6039) );
  FA1A U6217 ( .CI(n6038), .A(n6021), .B(n6032), .S(n6040), .CO(n6041) );
  FA1A U6218 ( .CI(n6036), .A(n6034), .B(n6017), .S(n6042), .CO(n6043) );
  FA1A U6219 ( .CI(n6040), .A(n6023), .B(n6019), .S(n6044), .CO(n6045) );
  FA1A U6220 ( .CI(n6027), .A(n6042), .B(n6025), .S(n6046), .CO(n6047) );
  FA1A U6221 ( .CI(n6046), .A(n6029), .B(n6044), .S(n6048), .CO(n6049) );
  HA1 U6222 ( .A(n5848), .B(n4323), .S(n6050), .CO(n6051) );
  FA1A U6223 ( .CI(n3747), .A(n3683), .B(n4003), .S(n6052), .CO(n6053) );
  FA1A U6224 ( .CI(n4195), .A(n4259), .B(n4131), .S(n6054), .CO(n6055) );
  FA1A U6225 ( .CI(n3939), .A(n4067), .B(n3811), .S(n6056), .CO(n6057) );
  FA1A U6226 ( .CI(n6033), .A(n6050), .B(n3875), .S(n6058), .CO(n6059) );
  FA1A U6227 ( .CI(n6054), .A(n6056), .B(n6035), .S(n6060), .CO(n6061) );
  FA1A U6228 ( .CI(n6052), .A(n6039), .B(n6037), .S(n6062), .CO(n6063) );
  FA1A U6229 ( .CI(n6062), .A(n6041), .B(n6058), .S(n6064), .CO(n6065) );
  FA1A U6230 ( .CI(n6064), .A(n6060), .B(n6043), .S(n6066), .CO(n6067) );
  FA1A U6231 ( .CI(n6066), .A(n6047), .B(n6045), .S(n6068), .CO(n6069) );
  FA1A U6232 ( .CI(n4324), .A(n4260), .B(n10888), .S(n6070), .CO(n6071) );
  FA1A U6233 ( .CI(n6051), .A(n3684), .B(n4004), .S(n6072), .CO(n6073) );
  FA1A U6234 ( .CI(n3748), .A(n4196), .B(n3940), .S(n6074), .CO(n6075) );
  FA1A U6235 ( .CI(n4068), .A(n4132), .B(n3812), .S(n6076), .CO(n6077) );
  FA1A U6236 ( .CI(n6053), .A(n6070), .B(n3876), .S(n6078), .CO(n6079) );
  FA1A U6237 ( .CI(n6074), .A(n6072), .B(n6055), .S(n6080), .CO(n6081) );
  FA1A U6238 ( .CI(n6059), .A(n6076), .B(n6057), .S(n6082), .CO(n6083) );
  FA1A U6239 ( .CI(n6082), .A(n6061), .B(n6078), .S(n6084), .CO(n6085) );
  FA1A U6240 ( .CI(n6084), .A(n6080), .B(n6063), .S(n6086), .CO(n6087) );
  FA1A U6241 ( .CI(n6086), .A(n6067), .B(n6065), .S(n6088), .CO(n6089) );
  HA1 U6242 ( .A(n5849), .B(n4389), .S(n6090), .CO(n6091) );
  FA1A U6243 ( .CI(n4261), .A(n4325), .B(n4005), .S(n6092), .CO(n6093) );
  FA1A U6244 ( .CI(n3749), .A(n3685), .B(n4069), .S(n6094), .CO(n6095) );
  FA1A U6245 ( .CI(n4133), .A(n4197), .B(n3813), .S(n6096), .CO(n6097) );
  FA1A U6246 ( .CI(n6090), .A(n3941), .B(n3877), .S(n6098), .CO(n6099) );
  FA1A U6247 ( .CI(n6098), .A(n6096), .B(n6071), .S(n6100), .CO(n6101) );
  FA1A U6248 ( .CI(n6092), .A(n6094), .B(n6073), .S(n6102), .CO(n6103) );
  FA1A U6249 ( .CI(n6079), .A(n6077), .B(n6075), .S(n6104), .CO(n6105) );
  FA1A U6250 ( .CI(n6104), .A(n6102), .B(n6100), .S(n6106), .CO(n6107) );
  FA1A U6251 ( .CI(n6085), .A(n6083), .B(n6081), .S(n6108), .CO(n6109) );
  FA1A U6252 ( .CI(n6108), .A(n6087), .B(n6106), .S(n6110), .CO(n6111) );
  FA1A U6253 ( .CI(n4390), .A(n4326), .B(n10887), .S(n6112), .CO(n6113) );
  FA1A U6254 ( .CI(n6091), .A(n4262), .B(n4006), .S(n6114), .CO(n6115) );
  FA1A U6255 ( .CI(n3750), .A(n3686), .B(n3942), .S(n6116), .CO(n6117) );
  FA1A U6256 ( .CI(n4134), .A(n4198), .B(n3814), .S(n6118), .CO(n6119) );
  FA1A U6257 ( .CI(n6112), .A(n4070), .B(n3878), .S(n6120), .CO(n6121) );
  FA1A U6258 ( .CI(n6120), .A(n6118), .B(n6093), .S(n6122), .CO(n6123) );
  FA1A U6259 ( .CI(n6099), .A(n6114), .B(n6095), .S(n6124), .CO(n6125) );
  FA1A U6260 ( .CI(n6101), .A(n6116), .B(n6097), .S(n6126), .CO(n6127) );
  FA1A U6261 ( .CI(n6105), .A(n6122), .B(n6103), .S(n6128), .CO(n6129) );
  FA1A U6262 ( .CI(n6107), .A(n6126), .B(n6124), .S(n6130), .CO(n6131) );
  FA1A U6263 ( .CI(n6130), .A(n6109), .B(n6128), .S(n6132), .CO(n6133) );
  HA1 U6264 ( .A(n5850), .B(n4455), .S(n6134), .CO(n6135) );
  FA1A U6265 ( .CI(n3751), .A(n3687), .B(n4007), .S(n6136), .CO(n6137) );
  FA1A U6266 ( .CI(n4327), .A(n4391), .B(n4199), .S(n6138), .CO(n6139) );
  FA1A U6267 ( .CI(n4135), .A(n4263), .B(n3815), .S(n6140), .CO(n6141) );
  FA1A U6268 ( .CI(n3943), .A(n4071), .B(n3879), .S(n6142), .CO(n6143) );
  FA1A U6269 ( .CI(n6142), .A(n6113), .B(n6134), .S(n6144), .CO(n6145) );
  FA1A U6270 ( .CI(n6121), .A(n6140), .B(n6115), .S(n6146), .CO(n6147) );
  FA1A U6271 ( .CI(n6138), .A(n6136), .B(n6117), .S(n6148), .CO(n6149) );
  FA1A U6272 ( .CI(n6123), .A(n6144), .B(n6119), .S(n6150), .CO(n6151) );
  FA1A U6273 ( .CI(n6148), .A(n6146), .B(n6125), .S(n6152), .CO(n6153) );
  FA1A U6274 ( .CI(n6129), .A(n6150), .B(n6127), .S(n6154), .CO(n6155) );
  FA1A U6275 ( .CI(n6154), .A(n6131), .B(n6152), .S(n6156), .CO(n6157) );
  FA1A U6276 ( .CI(n4456), .A(n4392), .B(n10886), .S(n6158), .CO(n6159) );
  FA1A U6277 ( .CI(n6135), .A(n3688), .B(n4072), .S(n6160), .CO(n6161) );
  FA1A U6278 ( .CI(n3816), .A(n3752), .B(n4136), .S(n6162), .CO(n6163) );
  FA1A U6279 ( .CI(n4264), .A(n4328), .B(n3880), .S(n6164), .CO(n6165) );
  FA1A U6280 ( .CI(n4008), .A(n4200), .B(n3944), .S(n6166), .CO(n6167) );
  FA1A U6281 ( .CI(n6166), .A(n6143), .B(n6158), .S(n6168), .CO(n6169) );
  FA1A U6282 ( .CI(n6162), .A(n6164), .B(n6137), .S(n6170), .CO(n6171) );
  FA1A U6283 ( .CI(n6160), .A(n6141), .B(n6139), .S(n6172), .CO(n6173) );
  FA1A U6284 ( .CI(n6170), .A(n6172), .B(n6145), .S(n6174), .CO(n6175) );
  FA1A U6285 ( .CI(n6147), .A(n6149), .B(n6168), .S(n6176), .CO(n6177) );
  FA1A U6286 ( .CI(n6153), .A(n6174), .B(n6151), .S(n6178), .CO(n6179) );
  FA1A U6287 ( .CI(n6178), .A(n6155), .B(n6176), .S(n6180), .CO(n6181) );
  HA1 U6288 ( .A(n5851), .B(n4521), .S(n6182), .CO(n6183) );
  FA1A U6289 ( .CI(n4393), .A(n4457), .B(n4073), .S(n6184), .CO(n6185) );
  FA1A U6290 ( .CI(n3689), .A(n4329), .B(n4009), .S(n6186), .CO(n6187) );
  FA1A U6291 ( .CI(n4265), .A(n3753), .B(n4137), .S(n6188), .CO(n6189) );
  FA1A U6292 ( .CI(n3945), .A(n4201), .B(n3817), .S(n6190), .CO(n6191) );
  FA1A U6293 ( .CI(n6159), .A(n6182), .B(n3881), .S(n6192), .CO(n6193) );
  FA1A U6294 ( .CI(n6188), .A(n6190), .B(n6165), .S(n6194), .CO(n6195) );
  FA1A U6295 ( .CI(n6186), .A(n6184), .B(n6161), .S(n6196), .CO(n6197) );
  FA1A U6296 ( .CI(n6192), .A(n6167), .B(n6163), .S(n6198), .CO(n6199) );
  FA1A U6297 ( .CI(n6198), .A(n6196), .B(n6169), .S(n6200), .CO(n6201) );
  FA1A U6298 ( .CI(n6194), .A(n6173), .B(n6171), .S(n6202), .CO(n6203) );
  FA1A U6299 ( .CI(n6202), .A(n6200), .B(n6177), .S(n6204), .CO(n6205) );
  FA1A U6300 ( .CI(n6204), .A(n6179), .B(n6175), .S(n6206), .CO(n6207) );
  FA1A U6301 ( .CI(n4522), .A(n4458), .B(n10885), .S(n6208), .CO(n6209) );
  FA1A U6302 ( .CI(n6183), .A(n4394), .B(n4074), .S(n6210), .CO(n6211) );
  FA1A U6303 ( .CI(n4266), .A(n4330), .B(n4010), .S(n6212), .CO(n6213) );
  FA1A U6304 ( .CI(n4138), .A(n4202), .B(n3690), .S(n6214), .CO(n6215) );
  FA1A U6305 ( .CI(n3882), .A(n3946), .B(n3754), .S(n6216), .CO(n6217) );
  FA1A U6306 ( .CI(n6185), .A(n6208), .B(n3818), .S(n6218), .CO(n6219) );
  FA1A U6307 ( .CI(n6214), .A(n6216), .B(n6191), .S(n6220), .CO(n6221) );
  FA1A U6308 ( .CI(n6212), .A(n6210), .B(n6187), .S(n6222), .CO(n6223) );
  FA1A U6309 ( .CI(n6218), .A(n6193), .B(n6189), .S(n6224), .CO(n6225) );
  FA1A U6310 ( .CI(n6199), .A(n6220), .B(n6195), .S(n6226), .CO(n6227) );
  FA1A U6311 ( .CI(n6224), .A(n6222), .B(n6197), .S(n6228), .CO(n6229) );
  FA1A U6312 ( .CI(n6228), .A(n6226), .B(n6201), .S(n6230), .CO(n6231) );
  FA1A U6313 ( .CI(n6230), .A(n6205), .B(n6203), .S(n6232), .CO(n6233) );
  HA1 U6314 ( .A(n5852), .B(n4587), .S(n6234), .CO(n6235) );
  FA1A U6315 ( .CI(n3755), .A(n3691), .B(n4075), .S(n6236), .CO(n6237) );
  FA1A U6316 ( .CI(n3883), .A(n3819), .B(n4267), .S(n6238), .CO(n6239) );
  FA1A U6317 ( .CI(n4459), .A(n4523), .B(n4395), .S(n6240), .CO(n6241) );
  FA1A U6318 ( .CI(n4203), .A(n4331), .B(n3947), .S(n6242), .CO(n6243) );
  FA1A U6319 ( .CI(n6234), .A(n4011), .B(n4139), .S(n6244), .CO(n6245) );
  FA1A U6320 ( .CI(n6244), .A(n6242), .B(n6209), .S(n6246), .CO(n6247) );
  FA1A U6321 ( .CI(n6238), .A(n6240), .B(n6211), .S(n6248), .CO(n6249) );
  FA1A U6322 ( .CI(n6236), .A(n6217), .B(n6213), .S(n6250), .CO(n6251) );
  FA1A U6323 ( .CI(n6246), .A(n6219), .B(n6215), .S(n6252), .CO(n6253) );
  FA1A U6324 ( .CI(n6250), .A(n6248), .B(n6221), .S(n6254), .CO(n6255) );
  FA1A U6325 ( .CI(n6252), .A(n6225), .B(n6223), .S(n6256), .CO(n6257) );
  FA1A U6326 ( .CI(n6229), .A(n6254), .B(n6227), .S(n6258), .CO(n6259) );
  FA1A U6327 ( .CI(n6258), .A(n6231), .B(n6256), .S(n6260), .CO(n6261) );
  FA1A U6328 ( .CI(n4588), .A(n4524), .B(n10884), .S(n6262), .CO(n6263) );
  FA1A U6329 ( .CI(n6235), .A(n3692), .B(n4140), .S(n6264), .CO(n6265) );
  FA1A U6330 ( .CI(n4460), .A(n3756), .B(n4076), .S(n6266), .CO(n6267) );
  FA1A U6331 ( .CI(n4268), .A(n4396), .B(n4332), .S(n6268), .CO(n6269) );
  FA1A U6332 ( .CI(n4012), .A(n4204), .B(n3820), .S(n6270), .CO(n6271) );
  FA1A U6333 ( .CI(n6262), .A(n3884), .B(n3948), .S(n6272), .CO(n6273) );
  FA1A U6334 ( .CI(n6272), .A(n6270), .B(n6241), .S(n6274), .CO(n6275) );
  FA1A U6335 ( .CI(n6245), .A(n6268), .B(n6237), .S(n6276), .CO(n6277) );
  FA1A U6336 ( .CI(n6264), .A(n6266), .B(n6239), .S(n6278), .CO(n6279) );
  FA1A U6337 ( .CI(n6249), .A(n6247), .B(n6243), .S(n6280), .CO(n6281) );
  FA1A U6338 ( .CI(n6276), .A(n6274), .B(n6251), .S(n6282), .CO(n6283) );
  FA1A U6339 ( .CI(n6280), .A(n6253), .B(n6278), .S(n6284), .CO(n6285) );
  FA1A U6340 ( .CI(n6257), .A(n6282), .B(n6255), .S(n6286), .CO(n6287) );
  FA1A U6341 ( .CI(n6286), .A(n6259), .B(n6284), .S(n6288), .CO(n6289) );
  HA1 U6342 ( .A(n5853), .B(n4653), .S(n6290), .CO(n6291) );
  FA1A U6343 ( .CI(n4525), .A(n4589), .B(n4141), .S(n6292), .CO(n6293) );
  FA1A U6344 ( .CI(n3757), .A(n3693), .B(n4077), .S(n6294), .CO(n6295) );
  FA1A U6345 ( .CI(n3885), .A(n3821), .B(n4269), .S(n6296), .CO(n6297) );
  FA1A U6346 ( .CI(n4397), .A(n4461), .B(n3949), .S(n6298), .CO(n6299) );
  FA1A U6347 ( .CI(n4205), .A(n4013), .B(n4333), .S(n6300), .CO(n6301) );
  FA1A U6348 ( .CI(n6300), .A(n6263), .B(n6290), .S(n6302), .CO(n6303) );
  FA1A U6349 ( .CI(n6273), .A(n6298), .B(n6269), .S(n6304), .CO(n6305) );
  FA1A U6350 ( .CI(n6294), .A(n6292), .B(n6267), .S(n6306), .CO(n6307) );
  FA1A U6351 ( .CI(n6296), .A(n6271), .B(n6265), .S(n6308), .CO(n6309) );
  FA1A U6352 ( .CI(n6308), .A(n6275), .B(n6302), .S(n6310), .CO(n6311) );
  FA1A U6353 ( .CI(n6306), .A(n6304), .B(n6277), .S(n6312), .CO(n6313) );
  FA1A U6354 ( .CI(n6281), .A(n6310), .B(n6279), .S(n6314), .CO(n6315) );
  FA1A U6355 ( .CI(n6285), .A(n6312), .B(n6283), .S(n6316), .CO(n6317) );
  FA1A U6356 ( .CI(n6316), .A(n6287), .B(n6314), .S(n6318), .CO(n6319) );
  FA1A U6357 ( .CI(n4654), .A(n4590), .B(n10883), .S(n6320), .CO(n6321) );
  FA1A U6358 ( .CI(n6291), .A(n3694), .B(n4142), .S(n6322), .CO(n6323) );
  FA1A U6359 ( .CI(n3822), .A(n3758), .B(n4206), .S(n6324), .CO(n6325) );
  FA1A U6360 ( .CI(n3886), .A(n4526), .B(n4334), .S(n6326), .CO(n6327) );
  FA1A U6361 ( .CI(n4398), .A(n4462), .B(n3950), .S(n6328), .CO(n6329) );
  FA1A U6362 ( .CI(n4078), .A(n4014), .B(n4270), .S(n6330), .CO(n6331) );
  FA1A U6363 ( .CI(n6330), .A(n6301), .B(n6320), .S(n6332), .CO(n6333) );
  FA1A U6364 ( .CI(n6324), .A(n6328), .B(n6297), .S(n6334), .CO(n6335) );
  FA1A U6365 ( .CI(n6322), .A(n6326), .B(n6293), .S(n6336), .CO(n6337) );
  FA1A U6366 ( .CI(n6303), .A(n6299), .B(n6295), .S(n6338), .CO(n6339) );
  FA1A U6367 ( .CI(n6334), .A(n6336), .B(n6332), .S(n6340), .CO(n6341) );
  FA1A U6368 ( .CI(n6338), .A(n6309), .B(n6305), .S(n6342), .CO(n6343) );
  FA1A U6369 ( .CI(n6311), .A(n6340), .B(n6307), .S(n6344), .CO(n6345) );
  FA1A U6370 ( .CI(n6344), .A(n6342), .B(n6313), .S(n6346), .CO(n6347) );
  FA1A U6371 ( .CI(n6346), .A(n6317), .B(n6315), .S(n6348), .CO(n6349) );
  HA1 U6372 ( .A(n5854), .B(n4719), .S(n6350), .CO(n6351) );
  FA1A U6373 ( .CI(n3759), .A(n3695), .B(n4143), .S(n6352), .CO(n6353) );
  FA1A U6374 ( .CI(n3887), .A(n3823), .B(n4335), .S(n6354), .CO(n6355) );
  FA1A U6375 ( .CI(n3951), .A(n4655), .B(n4399), .S(n6356), .CO(n6357) );
  FA1A U6376 ( .CI(n4527), .A(n4591), .B(n4015), .S(n6358), .CO(n6359) );
  FA1A U6377 ( .CI(n4271), .A(n4207), .B(n4079), .S(n6360), .CO(n6361) );
  FA1A U6378 ( .CI(n6321), .A(n6350), .B(n4463), .S(n6362), .CO(n6363) );
  FA1A U6379 ( .CI(n6358), .A(n6360), .B(n6329), .S(n6364), .CO(n6365) );
  FA1A U6380 ( .CI(n6352), .A(n6356), .B(n6327), .S(n6366), .CO(n6367) );
  FA1A U6381 ( .CI(n6354), .A(n6331), .B(n6323), .S(n6368), .CO(n6369) );
  FA1A U6382 ( .CI(n6333), .A(n6362), .B(n6325), .S(n6370), .CO(n6371) );
  FA1A U6383 ( .CI(n6339), .A(n6364), .B(n6335), .S(n6372), .CO(n6373) );
  FA1A U6384 ( .CI(n6368), .A(n6366), .B(n6337), .S(n6374), .CO(n6375) );
  FA1A U6385 ( .CI(n6374), .A(n6341), .B(n6370), .S(n6376), .CO(n6377) );
  FA1A U6386 ( .CI(n6376), .A(n6372), .B(n6343), .S(n6378), .CO(n6379) );
  FA1A U6387 ( .CI(n6378), .A(n6347), .B(n6345), .S(n6380), .CO(n6381) );
  FA1A U6388 ( .CI(n4720), .A(n4656), .B(n10882), .S(n6382), .CO(n6383) );
  FA1A U6389 ( .CI(n6351), .A(n3696), .B(n4208), .S(n6384), .CO(n6385) );
  FA1A U6390 ( .CI(n3760), .A(n4592), .B(n4272), .S(n6386), .CO(n6387) );
  FA1A U6391 ( .CI(n3824), .A(n4528), .B(n4144), .S(n6388), .CO(n6389) );
  FA1A U6392 ( .CI(n4400), .A(n4464), .B(n3888), .S(n6390), .CO(n6391) );
  FA1A U6393 ( .CI(n4080), .A(n4016), .B(n3952), .S(n6392), .CO(n6393) );
  FA1A U6394 ( .CI(n6353), .A(n6382), .B(n4336), .S(n6394), .CO(n6395) );
  FA1A U6395 ( .CI(n6390), .A(n6392), .B(n6361), .S(n6396), .CO(n6397) );
  FA1A U6396 ( .CI(n6386), .A(n6384), .B(n6357), .S(n6398), .CO(n6399) );
  FA1A U6397 ( .CI(n6388), .A(n6359), .B(n6355), .S(n6400), .CO(n6401) );
  FA1A U6398 ( .CI(n6400), .A(n6394), .B(n6363), .S(n6402), .CO(n6403) );
  FA1A U6399 ( .CI(n6396), .A(n6398), .B(n6365), .S(n6404), .CO(n6405) );
  FA1A U6400 ( .CI(n6371), .A(n6369), .B(n6367), .S(n6406), .CO(n6407) );
  FA1A U6401 ( .CI(n6406), .A(n6373), .B(n6402), .S(n6408), .CO(n6409) );
  FA1A U6402 ( .CI(n6408), .A(n6404), .B(n6375), .S(n6410), .CO(n6411) );
  FA1A U6403 ( .CI(n6410), .A(n6379), .B(n6377), .S(n6412), .CO(n6413) );
  HA1 U6404 ( .A(n5855), .B(n4785), .S(n6414), .CO(n6415) );
  FA1A U6405 ( .CI(n4721), .A(n3697), .B(n4209), .S(n6416), .CO(n6417) );
  FA1A U6406 ( .CI(n3761), .A(n4657), .B(n4337), .S(n6418), .CO(n6419) );
  FA1A U6407 ( .CI(n4593), .A(n3825), .B(n4273), .S(n6420), .CO(n6421) );
  FA1A U6408 ( .CI(n4465), .A(n4529), .B(n3889), .S(n6422), .CO(n6423) );
  FA1A U6409 ( .CI(n4145), .A(n4401), .B(n3953), .S(n6424), .CO(n6425) );
  FA1A U6410 ( .CI(n6414), .A(n4081), .B(n4017), .S(n6426), .CO(n6427) );
  FA1A U6411 ( .CI(n6426), .A(n6424), .B(n6383), .S(n6428), .CO(n6429) );
  FA1A U6412 ( .CI(n6418), .A(n6422), .B(n6391), .S(n6430), .CO(n6431) );
  FA1A U6413 ( .CI(n6420), .A(n6416), .B(n6385), .S(n6432), .CO(n6433) );
  FA1A U6414 ( .CI(n6389), .A(n6393), .B(n6387), .S(n6434), .CO(n6435) );
  FA1A U6415 ( .CI(n6434), .A(n6428), .B(n6395), .S(n6436), .CO(n6437) );
  FA1A U6416 ( .CI(n6430), .A(n6432), .B(n6397), .S(n6438), .CO(n6439) );
  FA1A U6417 ( .CI(n6403), .A(n6401), .B(n6399), .S(n6440), .CO(n6441) );
  FA1A U6418 ( .CI(n6440), .A(n6405), .B(n6436), .S(n6442), .CO(n6443) );
  FA1A U6419 ( .CI(n6442), .A(n6407), .B(n6438), .S(n6444), .CO(n6445) );
  FA1A U6420 ( .CI(n6444), .A(n6411), .B(n6409), .S(n6446), .CO(n6447) );
  FA1A U6421 ( .CI(n4786), .A(n4722), .B(n10881), .S(n6448), .CO(n6449) );
  FA1A U6422 ( .CI(n6415), .A(n4658), .B(n4210), .S(n6450), .CO(n6451) );
  FA1A U6423 ( .CI(n3762), .A(n3698), .B(n4146), .S(n6452), .CO(n6453) );
  FA1A U6424 ( .CI(n4530), .A(n4594), .B(n4274), .S(n6454), .CO(n6455) );
  FA1A U6425 ( .CI(n4402), .A(n4466), .B(n3826), .S(n6456), .CO(n6457) );
  FA1A U6426 ( .CI(n4082), .A(n4338), .B(n3890), .S(n6458), .CO(n6459) );
  FA1A U6427 ( .CI(n6448), .A(n4018), .B(n3954), .S(n6460), .CO(n6461) );
  FA1A U6428 ( .CI(n6460), .A(n6458), .B(n6423), .S(n6462), .CO(n6463) );
  FA1A U6429 ( .CI(n6427), .A(n6456), .B(n6421), .S(n6464), .CO(n6465) );
  FA1A U6430 ( .CI(n6452), .A(n6450), .B(n6419), .S(n6466), .CO(n6467) );
  FA1A U6431 ( .CI(n6454), .A(n6425), .B(n6417), .S(n6468), .CO(n6469) );
  FA1A U6432 ( .CI(n6466), .A(n6468), .B(n6429), .S(n6470), .CO(n6471) );
  FA1A U6433 ( .CI(n6462), .A(n6464), .B(n6431), .S(n6472), .CO(n6473) );
  FA1A U6434 ( .CI(n6437), .A(n6435), .B(n6433), .S(n6474), .CO(n6475) );
  FA1A U6435 ( .CI(n6441), .A(n6472), .B(n6470), .S(n6476), .CO(n6477) );
  FA1A U6436 ( .CI(n6443), .A(n6474), .B(n6439), .S(n6478), .CO(n6479) );
  FA1A U6437 ( .CI(n6478), .A(n6445), .B(n6476), .S(n6480), .CO(n6481) );
  HA1 U6438 ( .A(n5856), .B(n4851), .S(n6482), .CO(n6483) );
  FA1A U6439 ( .CI(n4787), .A(n3699), .B(n4211), .S(n6484), .CO(n6485) );
  FA1A U6440 ( .CI(n4659), .A(n4723), .B(n4339), .S(n6486), .CO(n6487) );
  FA1A U6441 ( .CI(n3827), .A(n3763), .B(n4147), .S(n6488), .CO(n6489) );
  FA1A U6442 ( .CI(n4531), .A(n4595), .B(n3891), .S(n6490), .CO(n6491) );
  FA1A U6443 ( .CI(n4403), .A(n4467), .B(n3955), .S(n6492), .CO(n6493) );
  FA1A U6444 ( .CI(n4083), .A(n4275), .B(n4019), .S(n6494), .CO(n6495) );
  FA1A U6445 ( .CI(n6494), .A(n6449), .B(n6482), .S(n6496), .CO(n6497) );
  FA1A U6446 ( .CI(n6461), .A(n6492), .B(n6457), .S(n6498), .CO(n6499) );
  FA1A U6447 ( .CI(n6488), .A(n6490), .B(n6455), .S(n6500), .CO(n6501) );
  FA1A U6448 ( .CI(n6486), .A(n6484), .B(n6451), .S(n6502), .CO(n6503) );
  FA1A U6449 ( .CI(n6496), .A(n6459), .B(n6453), .S(n6504), .CO(n6505) );
  FA1A U6450 ( .CI(n6504), .A(n6502), .B(n6463), .S(n6506), .CO(n6507) );
  FA1A U6451 ( .CI(n6498), .A(n6500), .B(n6465), .S(n6508), .CO(n6509) );
  FA1A U6452 ( .CI(n6471), .A(n6469), .B(n6467), .S(n6510), .CO(n6511) );
  FA1A U6453 ( .CI(n6475), .A(n6506), .B(n6473), .S(n6512), .CO(n6513) );
  FA1A U6454 ( .CI(n6477), .A(n6510), .B(n6508), .S(n6514), .CO(n6515) );
  FA1A U6455 ( .CI(n6514), .A(n6479), .B(n6512), .S(n6516), .CO(n6517) );
  FA1A U6456 ( .CI(n4852), .A(n4788), .B(n10880), .S(n6518), .CO(n6519) );
  FA1A U6457 ( .CI(n6483), .A(n4724), .B(n4276), .S(n6520), .CO(n6521) );
  FA1A U6458 ( .CI(n4660), .A(n3700), .B(n4212), .S(n6522), .CO(n6523) );
  FA1A U6459 ( .CI(n4532), .A(n4596), .B(n4148), .S(n6524), .CO(n6525) );
  FA1A U6460 ( .CI(n4404), .A(n4468), .B(n3764), .S(n6526), .CO(n6527) );
  FA1A U6461 ( .CI(n4084), .A(n4340), .B(n3828), .S(n6528), .CO(n6529) );
  FA1A U6462 ( .CI(n3956), .A(n4020), .B(n3892), .S(n6530), .CO(n6531) );
  FA1A U6463 ( .CI(n6530), .A(n6495), .B(n6518), .S(n6532), .CO(n6533) );
  FA1A U6464 ( .CI(n6526), .A(n6528), .B(n6491), .S(n6534), .CO(n6535) );
  FA1A U6465 ( .CI(n6520), .A(n6524), .B(n6489), .S(n6536), .CO(n6537) );
  FA1A U6466 ( .CI(n6522), .A(n6493), .B(n6485), .S(n6538), .CO(n6539) );
  FA1A U6467 ( .CI(n6532), .A(n6497), .B(n6487), .S(n6540), .CO(n6541) );
  FA1A U6468 ( .CI(n6505), .A(n6538), .B(n6499), .S(n6542), .CO(n6543) );
  FA1A U6469 ( .CI(n6536), .A(n6534), .B(n6501), .S(n6544), .CO(n6545) );
  FA1A U6470 ( .CI(n6507), .A(n6540), .B(n6503), .S(n6546), .CO(n6547) );
  FA1A U6471 ( .CI(n6544), .A(n6542), .B(n6509), .S(n6548), .CO(n6549) );
  FA1A U6472 ( .CI(n6513), .A(n6546), .B(n6511), .S(n6550), .CO(n6551) );
  FA1A U6473 ( .CI(n6550), .A(n6515), .B(n6548), .S(n6552), .CO(n6553) );
  HA1 U6474 ( .A(n5857), .B(n4917), .S(n6554), .CO(n6555) );
  FA1A U6475 ( .CI(n3765), .A(n3701), .B(n4277), .S(n6556), .CO(n6557) );
  FA1A U6476 ( .CI(n4789), .A(n4853), .B(n4469), .S(n6558), .CO(n6559) );
  FA1A U6477 ( .CI(n3829), .A(n4725), .B(n4341), .S(n6560), .CO(n6561) );
  FA1A U6478 ( .CI(n4597), .A(n4661), .B(n4405), .S(n6562), .CO(n6563) );
  FA1A U6479 ( .CI(n4213), .A(n4533), .B(n3893), .S(n6564), .CO(n6565) );
  FA1A U6480 ( .CI(n4085), .A(n4149), .B(n3957), .S(n6566), .CO(n6567) );
  FA1A U6481 ( .CI(n6519), .A(n6554), .B(n4021), .S(n6568), .CO(n6569) );
  FA1A U6482 ( .CI(n6564), .A(n6566), .B(n6529), .S(n6570), .CO(n6571) );
  FA1A U6483 ( .CI(n6560), .A(n6562), .B(n6527), .S(n6572), .CO(n6573) );
  FA1A U6484 ( .CI(n6558), .A(n6556), .B(n6521), .S(n6574), .CO(n6575) );
  FA1A U6485 ( .CI(n6525), .A(n6531), .B(n6523), .S(n6576), .CO(n6577) );
  FA1A U6486 ( .CI(n6576), .A(n6533), .B(n6568), .S(n6578), .CO(n6579) );
  FA1A U6487 ( .CI(n6572), .A(n6574), .B(n6535), .S(n6580), .CO(n6581) );
  FA1A U6488 ( .CI(n6570), .A(n6539), .B(n6537), .S(n6582), .CO(n6583) );
  FA1A U6489 ( .CI(n6582), .A(n6541), .B(n6578), .S(n6584), .CO(n6585) );
  FA1A U6490 ( .CI(n6580), .A(n6545), .B(n6543), .S(n6586), .CO(n6587) );
  FA1A U6491 ( .CI(n6586), .A(n6584), .B(n6547), .S(n6588), .CO(n6589) );
  FA1A U6492 ( .CI(n6588), .A(n6551), .B(n6549), .S(n6590), .CO(n6591) );
  FA1A U6493 ( .CI(n4918), .A(n4854), .B(n10879), .S(n6592), .CO(n6593) );
  FA1A U6494 ( .CI(n6555), .A(n3702), .B(n4342), .S(n6594), .CO(n6595) );
  FA1A U6495 ( .CI(n3830), .A(n3766), .B(n4278), .S(n6596), .CO(n6597) );
  FA1A U6496 ( .CI(n3958), .A(n3894), .B(n4470), .S(n6598), .CO(n6599) );
  FA1A U6497 ( .CI(n4662), .A(n4726), .B(n4790), .S(n6600), .CO(n6601) );
  FA1A U6498 ( .CI(n4534), .A(n4598), .B(n4022), .S(n6602), .CO(n6603) );
  FA1A U6499 ( .CI(n4214), .A(n4406), .B(n4086), .S(n6604), .CO(n6605) );
  FA1A U6500 ( .CI(n6557), .A(n6592), .B(n4150), .S(n6606), .CO(n6607) );
  FA1A U6501 ( .CI(n6602), .A(n6604), .B(n6567), .S(n6608), .CO(n6609) );
  FA1A U6502 ( .CI(n6598), .A(n6600), .B(n6563), .S(n6610), .CO(n6611) );
  FA1A U6503 ( .CI(n6594), .A(n6596), .B(n6559), .S(n6612), .CO(n6613) );
  FA1A U6504 ( .CI(n6569), .A(n6565), .B(n6561), .S(n6614), .CO(n6615) );
  FA1A U6505 ( .CI(n6614), .A(n6571), .B(n6606), .S(n6616), .CO(n6617) );
  FA1A U6506 ( .CI(n6610), .A(n6612), .B(n6573), .S(n6618), .CO(n6619) );
  FA1A U6507 ( .CI(n6608), .A(n6577), .B(n6575), .S(n6620), .CO(n6621) );
  FA1A U6508 ( .CI(n6620), .A(n6583), .B(n6616), .S(n6622), .CO(n6623) );
  FA1A U6509 ( .CI(n6618), .A(n6581), .B(n6579), .S(n6624), .CO(n6625) );
  FA1A U6510 ( .CI(n6587), .A(n6624), .B(n6585), .S(n6626), .CO(n6627) );
  FA1A U6511 ( .CI(n6626), .A(n6589), .B(n6622), .S(n6628), .CO(n6629) );
  HA1 U6512 ( .A(n5858), .B(n4983), .S(n6630), .CO(n6631) );
  FA1A U6513 ( .CI(n4919), .A(n3703), .B(n4279), .S(n6632), .CO(n6633) );
  FA1A U6514 ( .CI(n3767), .A(n4855), .B(n4407), .S(n6634), .CO(n6635) );
  FA1A U6515 ( .CI(n4791), .A(n3831), .B(n4471), .S(n6636), .CO(n6637) );
  FA1A U6516 ( .CI(n3959), .A(n3895), .B(n4343), .S(n6638), .CO(n6639) );
  FA1A U6517 ( .CI(n4663), .A(n4727), .B(n4023), .S(n6640), .CO(n6641) );
  FA1A U6518 ( .CI(n4535), .A(n4599), .B(n4087), .S(n6642), .CO(n6643) );
  FA1A U6519 ( .CI(n6630), .A(n4215), .B(n4151), .S(n6644), .CO(n6645) );
  FA1A U6520 ( .CI(n6644), .A(n6642), .B(n6593), .S(n6646), .CO(n6647) );
  FA1A U6521 ( .CI(n6638), .A(n6640), .B(n6595), .S(n6648), .CO(n6649) );
  FA1A U6522 ( .CI(n6632), .A(n6636), .B(n6601), .S(n6650), .CO(n6651) );
  FA1A U6523 ( .CI(n6634), .A(n6605), .B(n6597), .S(n6652), .CO(n6653) );
  FA1A U6524 ( .CI(n6607), .A(n6603), .B(n6599), .S(n6654), .CO(n6655) );
  FA1A U6525 ( .CI(n6654), .A(n6652), .B(n6646), .S(n6656), .CO(n6657) );
  FA1A U6526 ( .CI(n6615), .A(n6650), .B(n6609), .S(n6658), .CO(n6659) );
  FA1A U6527 ( .CI(n6648), .A(n6613), .B(n6611), .S(n6660), .CO(n6661) );
  FA1A U6528 ( .CI(n6658), .A(n6660), .B(n6617), .S(n6662), .CO(n6663) );
  FA1A U6529 ( .CI(n6619), .A(n6621), .B(n6656), .S(n6664), .CO(n6665) );
  FA1A U6530 ( .CI(n6664), .A(n6662), .B(n6623), .S(n6666), .CO(n6667) );
  FA1A U6531 ( .CI(n6666), .A(n6627), .B(n6625), .S(n6668), .CO(n6669) );
  FA1A U6532 ( .CI(n4984), .A(n4920), .B(n10878), .S(n6670), .CO(n6671) );
  FA1A U6533 ( .CI(n6631), .A(n4856), .B(n4344), .S(n6672), .CO(n6673) );
  FA1A U6534 ( .CI(n3768), .A(n3704), .B(n4280), .S(n6674), .CO(n6675) );
  FA1A U6535 ( .CI(n4728), .A(n4792), .B(n4408), .S(n6676), .CO(n6677) );
  FA1A U6536 ( .CI(n3896), .A(n3832), .B(n4600), .S(n6678), .CO(n6679) );
  FA1A U6537 ( .CI(n4536), .A(n4664), .B(n3960), .S(n6680), .CO(n6681) );
  FA1A U6538 ( .CI(n4216), .A(n4472), .B(n4024), .S(n6682), .CO(n6683) );
  FA1A U6539 ( .CI(n6670), .A(n4152), .B(n4088), .S(n6684), .CO(n6685) );
  FA1A U6540 ( .CI(n6684), .A(n6682), .B(n6641), .S(n6686), .CO(n6687) );
  FA1A U6541 ( .CI(n6645), .A(n6680), .B(n6633), .S(n6688), .CO(n6689) );
  FA1A U6542 ( .CI(n6676), .A(n6678), .B(n6639), .S(n6690), .CO(n6691) );
  FA1A U6543 ( .CI(n6672), .A(n6674), .B(n6637), .S(n6692), .CO(n6693) );
  FA1A U6544 ( .CI(n6647), .A(n6643), .B(n6635), .S(n6694), .CO(n6695) );
  FA1A U6545 ( .CI(n6655), .A(n6692), .B(n6653), .S(n6696), .CO(n6697) );
  FA1A U6546 ( .CI(n6686), .A(n6688), .B(n6649), .S(n6698), .CO(n6699) );
  FA1A U6547 ( .CI(n6694), .A(n6690), .B(n6651), .S(n6700), .CO(n6701) );
  FA1A U6548 ( .CI(n6700), .A(n6698), .B(n6657), .S(n6702), .CO(n6703) );
  FA1A U6549 ( .CI(n6696), .A(n6661), .B(n6659), .S(n6704), .CO(n6705) );
  FA1A U6550 ( .CI(n6704), .A(n6702), .B(n6663), .S(n6706), .CO(n6707) );
  FA1A U6551 ( .CI(n6706), .A(n6667), .B(n6665), .S(n6708), .CO(n6709) );
  HA1 U6552 ( .A(n5859), .B(n5049), .S(n6710), .CO(n6711) );
  FA1A U6553 ( .CI(n4985), .A(n3705), .B(n4345), .S(n6712), .CO(n6713) );
  FA1A U6554 ( .CI(n3769), .A(n4921), .B(n4473), .S(n6714), .CO(n6715) );
  FA1A U6555 ( .CI(n3897), .A(n3833), .B(n4409), .S(n6716), .CO(n6717) );
  FA1A U6556 ( .CI(n3961), .A(n4857), .B(n4601), .S(n6718), .CO(n6719) );
  FA1A U6557 ( .CI(n4729), .A(n4793), .B(n4025), .S(n6720), .CO(n6721) );
  FA1A U6558 ( .CI(n4537), .A(n4665), .B(n4089), .S(n6722), .CO(n6723) );
  FA1A U6559 ( .CI(n4153), .A(n4217), .B(n4281), .S(n6724), .CO(n6725) );
  FA1A U6560 ( .CI(n6724), .A(n6671), .B(n6710), .S(n6726), .CO(n6727) );
  FA1A U6561 ( .CI(n6685), .A(n6722), .B(n6681), .S(n6728), .CO(n6729) );
  FA1A U6562 ( .CI(n6718), .A(n6720), .B(n6679), .S(n6730), .CO(n6731) );
  FA1A U6563 ( .CI(n6714), .A(n6712), .B(n6673), .S(n6732), .CO(n6733) );
  FA1A U6564 ( .CI(n6716), .A(n6683), .B(n6677), .S(n6734), .CO(n6735) );
  FA1A U6565 ( .CI(n6687), .A(n6726), .B(n6675), .S(n6736), .CO(n6737) );
  FA1A U6566 ( .CI(n6732), .A(n6734), .B(n6693), .S(n6738), .CO(n6739) );
  FA1A U6567 ( .CI(n6730), .A(n6728), .B(n6689), .S(n6740), .CO(n6741) );
  FA1A U6568 ( .CI(n6736), .A(n6695), .B(n6691), .S(n6742), .CO(n6743) );
  FA1A U6569 ( .CI(n6742), .A(n6701), .B(n6697), .S(n6744), .CO(n6745) );
  FA1A U6570 ( .CI(n6740), .A(n6738), .B(n6699), .S(n6746), .CO(n6747) );
  FA1A U6571 ( .CI(n6744), .A(n6746), .B(n6703), .S(n6748), .CO(n6749) );
  FA1A U6572 ( .CI(n6748), .A(n6707), .B(n6705), .S(n6750), .CO(n6751) );
  FA1A U6573 ( .CI(n5050), .A(n4986), .B(n10877), .S(n6752), .CO(n6753) );
  FA1A U6574 ( .CI(n6711), .A(n3706), .B(n4346), .S(n6754), .CO(n6755) );
  FA1A U6575 ( .CI(n3770), .A(n4922), .B(n4474), .S(n6756), .CO(n6757) );
  FA1A U6576 ( .CI(n4858), .A(n3834), .B(n4410), .S(n6758), .CO(n6759) );
  FA1A U6577 ( .CI(n3962), .A(n3898), .B(n4282), .S(n6760), .CO(n6761) );
  FA1A U6578 ( .CI(n4730), .A(n4794), .B(n4026), .S(n6762), .CO(n6763) );
  FA1A U6579 ( .CI(n4602), .A(n4666), .B(n4090), .S(n6764), .CO(n6765) );
  FA1A U6580 ( .CI(n4154), .A(n4218), .B(n4538), .S(n6766), .CO(n6767) );
  FA1A U6581 ( .CI(n6766), .A(n6725), .B(n6752), .S(n6768), .CO(n6769) );
  FA1A U6582 ( .CI(n6756), .A(n6764), .B(n6721), .S(n6770), .CO(n6771) );
  FA1A U6583 ( .CI(n6760), .A(n6762), .B(n6713), .S(n6772), .CO(n6773) );
  FA1A U6584 ( .CI(n6754), .A(n6758), .B(n6715), .S(n6774), .CO(n6775) );
  FA1A U6585 ( .CI(n6719), .A(n6723), .B(n6717), .S(n6776), .CO(n6777) );
  FA1A U6586 ( .CI(n6774), .A(n6776), .B(n6727), .S(n6778), .CO(n6779) );
  FA1A U6587 ( .CI(n6770), .A(n6772), .B(n6768), .S(n6780), .CO(n6781) );
  FA1A U6588 ( .CI(n6733), .A(n6735), .B(n6729), .S(n6782), .CO(n6783) );
  FA1A U6589 ( .CI(n6778), .A(n6737), .B(n6731), .S(n6784), .CO(n6785) );
  FA1A U6590 ( .CI(n6782), .A(n6739), .B(n6780), .S(n6786), .CO(n6787) );
  FA1A U6591 ( .CI(n6784), .A(n6743), .B(n6741), .S(n6788), .CO(n6789) );
  FA1A U6592 ( .CI(n6788), .A(n6747), .B(n6786), .S(n6790), .CO(n6791) );
  FA1A U6593 ( .CI(n6749), .A(n6790), .B(n6745), .S(n6792), .CO(n6793) );
  HA1 U6594 ( .A(n5860), .B(n5115), .S(n6794), .CO(n6795) );
  FA1A U6595 ( .CI(n5051), .A(n3707), .B(n4347), .S(n6796), .CO(n6797) );
  FA1A U6596 ( .CI(n4987), .A(n3771), .B(n4475), .S(n6798), .CO(n6799) );
  FA1A U6597 ( .CI(n4923), .A(n3835), .B(n4539), .S(n6800), .CO(n6801) );
  FA1A U6598 ( .CI(n4795), .A(n4859), .B(n4411), .S(n6802), .CO(n6803) );
  FA1A U6599 ( .CI(n4667), .A(n4731), .B(n3899), .S(n6804), .CO(n6805) );
  FA1A U6600 ( .CI(n4283), .A(n4603), .B(n3963), .S(n6806), .CO(n6807) );
  FA1A U6601 ( .CI(n4155), .A(n4091), .B(n4027), .S(n6808), .CO(n6809) );
  FA1A U6602 ( .CI(n6753), .A(n6794), .B(n4219), .S(n6810), .CO(n6811) );
  FA1A U6603 ( .CI(n6806), .A(n6808), .B(n6765), .S(n6812), .CO(n6813) );
  FA1A U6604 ( .CI(n6796), .A(n6804), .B(n6763), .S(n6814), .CO(n6815) );
  FA1A U6605 ( .CI(n6800), .A(n6798), .B(n6755), .S(n6816), .CO(n6817) );
  FA1A U6606 ( .CI(n6802), .A(n6767), .B(n6761), .S(n6818), .CO(n6819) );
  FA1A U6607 ( .CI(n6810), .A(n6757), .B(n6759), .S(n6820), .CO(n6821) );
  FA1A U6608 ( .CI(n6820), .A(n6818), .B(n6769), .S(n6822), .CO(n6823) );
  FA1A U6609 ( .CI(n6814), .A(n6816), .B(n6771), .S(n6824), .CO(n6825) );
  FA1A U6610 ( .CI(n6812), .A(n6777), .B(n6773), .S(n6826), .CO(n6827) );
  FA1A U6611 ( .CI(n6781), .A(n6779), .B(n6775), .S(n6828), .CO(n6829) );
  FA1A U6612 ( .CI(n6826), .A(n6824), .B(n6822), .S(n6830), .CO(n6831) );
  FA1A U6613 ( .CI(n6828), .A(n6785), .B(n6783), .S(n6832), .CO(n6833) );
  FA1A U6614 ( .CI(n6789), .A(n6830), .B(n6787), .S(n6834), .CO(n6835) );
  FA1A U6615 ( .CI(n6834), .A(n6791), .B(n6832), .S(n6836), .CO(n6837) );
  FA1A U6616 ( .CI(n5116), .A(n5052), .B(n10876), .S(n6838), .CO(n6839) );
  FA1A U6617 ( .CI(n6795), .A(n4988), .B(n4412), .S(n6840), .CO(n6841) );
  FA1A U6618 ( .CI(n3708), .A(n4924), .B(n4348), .S(n6842), .CO(n6843) );
  FA1A U6619 ( .CI(n3836), .A(n3772), .B(n4284), .S(n6844), .CO(n6845) );
  FA1A U6620 ( .CI(n3900), .A(n4860), .B(n4540), .S(n6846), .CO(n6847) );
  FA1A U6621 ( .CI(n4732), .A(n4796), .B(n3964), .S(n6848), .CO(n6849) );
  FA1A U6622 ( .CI(n4604), .A(n4668), .B(n4028), .S(n6850), .CO(n6851) );
  FA1A U6623 ( .CI(n4476), .A(n4156), .B(n4092), .S(n6852), .CO(n6853) );
  FA1A U6624 ( .CI(n6797), .A(n6838), .B(n4220), .S(n6854), .CO(n6855) );
  FA1A U6625 ( .CI(n6850), .A(n6852), .B(n6809), .S(n6856), .CO(n6857) );
  FA1A U6626 ( .CI(n6840), .A(n6848), .B(n6805), .S(n6858), .CO(n6859) );
  FA1A U6627 ( .CI(n6846), .A(n6844), .B(n6799), .S(n6860), .CO(n6861) );
  FA1A U6628 ( .CI(n6842), .A(n6803), .B(n6807), .S(n6862), .CO(n6863) );
  FA1A U6629 ( .CI(n6854), .A(n6811), .B(n6801), .S(n6864), .CO(n6865) );
  FA1A U6630 ( .CI(n6821), .A(n6862), .B(n6817), .S(n6866), .CO(n6867) );
  FA1A U6631 ( .CI(n6858), .A(n6856), .B(n6815), .S(n6868), .CO(n6869) );
  FA1A U6632 ( .CI(n6860), .A(n6819), .B(n6813), .S(n6870), .CO(n6871) );
  FA1A U6633 ( .CI(n6870), .A(n6823), .B(n6864), .S(n6872), .CO(n6873) );
  FA1A U6634 ( .CI(n6868), .A(n6866), .B(n6825), .S(n6874), .CO(n6875) );
  FA1A U6635 ( .CI(n6829), .A(n6872), .B(n6827), .S(n6876), .CO(n6877) );
  FA1A U6636 ( .CI(n6833), .A(n6874), .B(n6831), .S(n6878), .CO(n6879) );
  FA1A U6637 ( .CI(n6878), .A(n6835), .B(n6876), .S(n6880), .CO(n6881) );
  HA1 U6638 ( .A(n5861), .B(n5181), .S(n6882), .CO(n6883) );
  FA1A U6639 ( .CI(n3773), .A(n3709), .B(n4349), .S(n6884), .CO(n6885) );
  FA1A U6640 ( .CI(n3837), .A(n5117), .B(n4541), .S(n6886), .CO(n6887) );
  FA1A U6641 ( .CI(n3965), .A(n3901), .B(n4669), .S(n6888), .CO(n6889) );
  FA1A U6642 ( .CI(n5053), .A(n4029), .B(n4733), .S(n6890), .CO(n6891) );
  FA1A U6643 ( .CI(n4925), .A(n4989), .B(n4093), .S(n6892), .CO(n6893) );
  FA1A U6644 ( .CI(n4797), .A(n4861), .B(n4157), .S(n6894), .CO(n6895) );
  FA1A U6645 ( .CI(n4477), .A(n4605), .B(n4221), .S(n6896), .CO(n6897) );
  FA1A U6646 ( .CI(n6882), .A(n4413), .B(n4285), .S(n6898), .CO(n6899) );
  FA1A U6647 ( .CI(n6898), .A(n6896), .B(n6839), .S(n6900), .CO(n6901) );
  FA1A U6648 ( .CI(n6886), .A(n6894), .B(n6851), .S(n6902), .CO(n6903) );
  FA1A U6649 ( .CI(n6888), .A(n6884), .B(n6841), .S(n6904), .CO(n6905) );
  FA1A U6650 ( .CI(n6892), .A(n6890), .B(n6843), .S(n6906), .CO(n6907) );
  FA1A U6651 ( .CI(n6849), .A(n6853), .B(n6845), .S(n6908), .CO(n6909) );
  FA1A U6652 ( .CI(n6900), .A(n6855), .B(n6847), .S(n6910), .CO(n6911) );
  FA1A U6653 ( .CI(n6904), .A(n6908), .B(n6861), .S(n6912), .CO(n6913) );
  FA1A U6654 ( .CI(n6902), .A(n6906), .B(n6857), .S(n6914), .CO(n6915) );
  FA1A U6655 ( .CI(n6865), .A(n6863), .B(n6859), .S(n6916), .CO(n6917) );
  FA1A U6656 ( .CI(n6916), .A(n6867), .B(n6910), .S(n6918), .CO(n6919) );
  FA1A U6657 ( .CI(n6914), .A(n6912), .B(n6869), .S(n6920), .CO(n6921) );
  FA1A U6658 ( .CI(n6873), .A(n6918), .B(n6871), .S(n6922), .CO(n6923) );
  FA1A U6659 ( .CI(n6922), .A(n6920), .B(n6875), .S(n6924), .CO(n6925) );
  FA1A U6660 ( .CI(n6924), .A(n6879), .B(n6877), .S(n6926), .CO(n6927) );
  FA1A U6661 ( .CI(n5182), .A(n5118), .B(n10875), .S(n6928), .CO(n6929) );
  FA1A U6662 ( .CI(n6883), .A(n3710), .B(n4414), .S(n6930), .CO(n6931) );
  FA1A U6663 ( .CI(n3838), .A(n3774), .B(n4478), .S(n6932), .CO(n6933) );
  FA1A U6664 ( .CI(n5054), .A(n3902), .B(n4606), .S(n6934), .CO(n6935) );
  FA1A U6665 ( .CI(n3966), .A(n4990), .B(n4542), .S(n6936), .CO(n6937) );
  FA1A U6666 ( .CI(n4862), .A(n4926), .B(n4030), .S(n6938), .CO(n6939) );
  FA1A U6667 ( .CI(n4734), .A(n4798), .B(n4094), .S(n6940), .CO(n6941) );
  FA1A U6668 ( .CI(n4350), .A(n4670), .B(n4158), .S(n6942), .CO(n6943) );
  FA1A U6669 ( .CI(n6928), .A(n4286), .B(n4222), .S(n6944), .CO(n6945) );
  FA1A U6670 ( .CI(n6944), .A(n6942), .B(n6895), .S(n6946), .CO(n6947) );
  FA1A U6671 ( .CI(n6899), .A(n6940), .B(n6893), .S(n6948), .CO(n6949) );
  FA1A U6672 ( .CI(n6930), .A(n6938), .B(n6891), .S(n6950), .CO(n6951) );
  FA1A U6673 ( .CI(n6936), .A(n6932), .B(n6885), .S(n6952), .CO(n6953) );
  FA1A U6674 ( .CI(n6934), .A(n6889), .B(n6897), .S(n6954), .CO(n6955) );
  FA1A U6675 ( .CI(n6903), .A(n6901), .B(n6887), .S(n6956), .CO(n6957) );
  FA1A U6676 ( .CI(n6948), .A(n6946), .B(n6909), .S(n6958), .CO(n6959) );
  FA1A U6677 ( .CI(n6952), .A(n6950), .B(n6905), .S(n6960), .CO(n6961) );
  FA1A U6678 ( .CI(n6911), .A(n6954), .B(n6907), .S(n6962), .CO(n6963) );
  FA1A U6679 ( .CI(n6917), .A(n6913), .B(n6956), .S(n6964), .CO(n6965) );
  FA1A U6680 ( .CI(n6962), .A(n6958), .B(n6915), .S(n6966), .CO(n6967) );
  FA1A U6681 ( .CI(n6919), .A(n6964), .B(n6960), .S(n6968), .CO(n6969) );
  FA1A U6682 ( .CI(n6968), .A(n6966), .B(n6921), .S(n6970), .CO(n6971) );
  FA1A U6683 ( .CI(n6970), .A(n6925), .B(n6923), .S(n6972), .CO(n6973) );
  HA1 U6684 ( .A(n5862), .B(n5247), .S(n6974), .CO(n6975) );
  FA1A U6685 ( .CI(n3775), .A(n3711), .B(n4415), .S(n6976), .CO(n6977) );
  FA1A U6686 ( .CI(n3903), .A(n3839), .B(n4607), .S(n6978), .CO(n6979) );
  FA1A U6687 ( .CI(n4031), .A(n3967), .B(n4735), .S(n6980), .CO(n6981) );
  FA1A U6688 ( .CI(n5119), .A(n5183), .B(n4799), .S(n6982), .CO(n6983) );
  FA1A U6689 ( .CI(n4927), .A(n4991), .B(n5055), .S(n6984), .CO(n6985) );
  FA1A U6690 ( .CI(n4671), .A(n4863), .B(n4095), .S(n6986), .CO(n6987) );
  FA1A U6691 ( .CI(n4479), .A(n4543), .B(n4159), .S(n6988), .CO(n6989) );
  FA1A U6692 ( .CI(n4287), .A(n4351), .B(n4223), .S(n6990), .CO(n6991) );
  FA1A U6693 ( .CI(n6990), .A(n6929), .B(n6974), .S(n6992), .CO(n6993) );
  FA1A U6694 ( .CI(n6945), .A(n6988), .B(n6941), .S(n6994), .CO(n6995) );
  FA1A U6695 ( .CI(n6984), .A(n6986), .B(n6939), .S(n6996), .CO(n6997) );
  FA1A U6696 ( .CI(n6976), .A(n6982), .B(n6937), .S(n6998), .CO(n6999) );
  FA1A U6697 ( .CI(n6980), .A(n6978), .B(n6931), .S(n7000), .CO(n7001) );
  FA1A U6698 ( .CI(n6935), .A(n6933), .B(n6943), .S(n7002), .CO(n7003) );
  FA1A U6699 ( .CI(n7002), .A(n6947), .B(n6992), .S(n7004), .CO(n7005) );
  FA1A U6700 ( .CI(n6994), .A(n7000), .B(n6953), .S(n7006), .CO(n7007) );
  FA1A U6701 ( .CI(n6998), .A(n6996), .B(n6949), .S(n7008), .CO(n7009) );
  FA1A U6702 ( .CI(n7004), .A(n6955), .B(n6951), .S(n7010), .CO(n7011) );
  FA1A U6703 ( .CI(n6963), .A(n7008), .B(n6957), .S(n7012), .CO(n7013) );
  FA1A U6704 ( .CI(n7010), .A(n7006), .B(n6959), .S(n7014), .CO(n7015) );
  FA1A U6705 ( .CI(n6965), .A(n7012), .B(n6961), .S(n7016), .CO(n7017) );
  FA1A U6706 ( .CI(n7016), .A(n7014), .B(n6967), .S(n7018), .CO(n7019) );
  FA1A U6707 ( .CI(n7018), .A(n6971), .B(n6969), .S(n7020), .CO(n7021) );
  FA1A U6708 ( .CI(n5248), .A(n5184), .B(n10874), .S(n7022), .CO(n7023) );
  FA1A U6709 ( .CI(n6975), .A(n3712), .B(n4480), .S(n7024), .CO(n7025) );
  FA1A U6710 ( .CI(n3776), .A(n5120), .B(n4544), .S(n7026), .CO(n7027) );
  FA1A U6711 ( .CI(n4992), .A(n5056), .B(n4608), .S(n7028), .CO(n7029) );
  FA1A U6712 ( .CI(n4928), .A(n3840), .B(n4352), .S(n7030), .CO(n7031) );
  FA1A U6713 ( .CI(n4736), .A(n4800), .B(n4864), .S(n7032), .CO(n7033) );
  FA1A U6714 ( .CI(n4416), .A(n4672), .B(n3904), .S(n7034), .CO(n7035) );
  FA1A U6715 ( .CI(n4224), .A(n4288), .B(n3968), .S(n7036), .CO(n7037) );
  FA1A U6716 ( .CI(n4096), .A(n4160), .B(n4032), .S(n7038), .CO(n7039) );
  FA1A U6717 ( .CI(n7038), .A(n6991), .B(n7022), .S(n7040), .CO(n7041) );
  FA1A U6718 ( .CI(n7034), .A(n7036), .B(n6987), .S(n7042), .CO(n7043) );
  FA1A U6719 ( .CI(n7024), .A(n7032), .B(n6985), .S(n7044), .CO(n7045) );
  FA1A U6720 ( .CI(n7028), .A(n7026), .B(n6977), .S(n7046), .CO(n7047) );
  FA1A U6721 ( .CI(n7030), .A(n6989), .B(n6979), .S(n7048), .CO(n7049) );
  FA1A U6722 ( .CI(n6993), .A(n6981), .B(n6983), .S(n7050), .CO(n7051) );
  FA1A U6723 ( .CI(n7042), .A(n7048), .B(n7040), .S(n7052), .CO(n7053) );
  FA1A U6724 ( .CI(n7050), .A(n7044), .B(n6995), .S(n7054), .CO(n7055) );
  FA1A U6725 ( .CI(n7046), .A(n7003), .B(n6997), .S(n7056), .CO(n7057) );
  FA1A U6726 ( .CI(n7052), .A(n7001), .B(n6999), .S(n7058), .CO(n7059) );
  FA1A U6727 ( .CI(n7054), .A(n7056), .B(n7005), .S(n7060), .CO(n7061) );
  FA1A U6728 ( .CI(n7058), .A(n7009), .B(n7007), .S(n7062), .CO(n7063) );
  FA1A U6729 ( .CI(n7013), .A(n7060), .B(n7011), .S(n7064), .CO(n7065) );
  FA1A U6730 ( .CI(n7064), .A(n7062), .B(n7015), .S(n7066), .CO(n7067) );
  FA1A U6731 ( .CI(n7066), .A(n7019), .B(n7017), .S(n7068), .CO(n7069) );
  HA1 U6732 ( .A(n5863), .B(n5313), .S(n7070), .CO(n7071) );
  FA1A U6733 ( .CI(n3713), .A(n5249), .B(n4417), .S(n7072), .CO(n7073) );
  FA1A U6734 ( .CI(n5185), .A(n3777), .B(n4609), .S(n7074), .CO(n7075) );
  FA1A U6735 ( .CI(n5057), .A(n5121), .B(n4545), .S(n7076), .CO(n7077) );
  FA1A U6736 ( .CI(n4929), .A(n4993), .B(n4481), .S(n7078), .CO(n7079) );
  FA1A U6737 ( .CI(n3841), .A(n4865), .B(n4353), .S(n7080), .CO(n7081) );
  FA1A U6738 ( .CI(n4737), .A(n4801), .B(n3905), .S(n7082), .CO(n7083) );
  FA1A U6739 ( .CI(n4289), .A(n4673), .B(n3969), .S(n7084), .CO(n7085) );
  FA1A U6740 ( .CI(n4161), .A(n4225), .B(n4033), .S(n7086), .CO(n7087) );
  FA1A U6741 ( .CI(n7023), .A(n7070), .B(n4097), .S(n7088), .CO(n7089) );
  FA1A U6742 ( .CI(n7084), .A(n7086), .B(n7037), .S(n7090), .CO(n7091) );
  FA1A U6743 ( .CI(n7080), .A(n7082), .B(n7035), .S(n7092), .CO(n7093) );
  FA1A U6744 ( .CI(n7072), .A(n7078), .B(n7031), .S(n7094), .CO(n7095) );
  FA1A U6745 ( .CI(n7076), .A(n7074), .B(n7025), .S(n7096), .CO(n7097) );
  FA1A U6746 ( .CI(n7033), .A(n7029), .B(n7027), .S(n7098), .CO(n7099) );
  FA1A U6747 ( .CI(n7041), .A(n7088), .B(n7039), .S(n7100), .CO(n7101) );
  FA1A U6748 ( .CI(n7051), .A(n7098), .B(n7049), .S(n7102), .CO(n7103) );
  FA1A U6749 ( .CI(n7090), .A(n7092), .B(n7047), .S(n7104), .CO(n7105) );
  FA1A U6750 ( .CI(n7096), .A(n7094), .B(n7043), .S(n7106), .CO(n7107) );
  FA1A U6751 ( .CI(n7053), .A(n7100), .B(n7045), .S(n7108), .CO(n7109) );
  FA1A U6752 ( .CI(n7059), .A(n7102), .B(n7055), .S(n7110), .CO(n7111) );
  FA1A U6753 ( .CI(n7106), .A(n7104), .B(n7057), .S(n7112), .CO(n7113) );
  FA1A U6754 ( .CI(n7063), .A(n7061), .B(n7108), .S(n7114), .CO(n7115) );
  FA1A U6755 ( .CI(n7114), .A(n7110), .B(n7112), .S(n7116), .CO(n7117) );
  FA1A U6756 ( .CI(n7116), .A(n7067), .B(n7065), .S(n7118), .CO(n7119) );
  FA1A U6757 ( .CI(n5314), .A(n5250), .B(n10873), .S(n7120), .CO(n7121) );
  FA1A U6758 ( .CI(n7071), .A(n3714), .B(n4546), .S(n7122), .CO(n7123) );
  FA1A U6759 ( .CI(n3778), .A(n5186), .B(n4482), .S(n7124), .CO(n7125) );
  FA1A U6760 ( .CI(n3842), .A(n5122), .B(n4610), .S(n7126), .CO(n7127) );
  FA1A U6761 ( .CI(n4994), .A(n5058), .B(n4674), .S(n7128), .CO(n7129) );
  FA1A U6762 ( .CI(n3970), .A(n3906), .B(n4866), .S(n7130), .CO(n7131) );
  FA1A U6763 ( .CI(n4802), .A(n4930), .B(n4034), .S(n7132), .CO(n7133) );
  FA1A U6764 ( .CI(n4418), .A(n4738), .B(n4098), .S(n7134), .CO(n7135) );
  FA1A U6765 ( .CI(n4290), .A(n4354), .B(n4162), .S(n7136), .CO(n7137) );
  FA1A U6766 ( .CI(n7073), .A(n7120), .B(n4226), .S(n7138), .CO(n7139) );
  FA1A U6767 ( .CI(n7134), .A(n7136), .B(n7085), .S(n7140), .CO(n7141) );
  FA1A U6768 ( .CI(n7130), .A(n7132), .B(n7083), .S(n7142), .CO(n7143) );
  FA1A U6769 ( .CI(n7122), .A(n7128), .B(n7081), .S(n7144), .CO(n7145) );
  FA1A U6770 ( .CI(n7124), .A(n7126), .B(n7075), .S(n7146), .CO(n7147) );
  FA1A U6771 ( .CI(n7087), .A(n7079), .B(n7077), .S(n7148), .CO(n7149) );
  FA1A U6772 ( .CI(n7148), .A(n7138), .B(n7089), .S(n7150), .CO(n7151) );
  FA1A U6773 ( .CI(n7142), .A(n7146), .B(n7097), .S(n7152), .CO(n7153) );
  FA1A U6774 ( .CI(n7144), .A(n7140), .B(n7091), .S(n7154), .CO(n7155) );
  FA1A U6775 ( .CI(n7095), .A(n7099), .B(n7093), .S(n7156), .CO(n7157) );
  FA1A U6776 ( .CI(n7156), .A(n7150), .B(n7101), .S(n7158), .CO(n7159) );
  FA1A U6777 ( .CI(n7152), .A(n7154), .B(n7103), .S(n7160), .CO(n7161) );
  FA1A U6778 ( .CI(n7109), .A(n7107), .B(n7105), .S(n7162), .CO(n7163) );
  FA1A U6779 ( .CI(n7162), .A(n7111), .B(n7158), .S(n7164), .CO(n7165) );
  FA1A U6780 ( .CI(n7164), .A(n7160), .B(n7113), .S(n7166), .CO(n7167) );
  FA1A U6781 ( .CI(n7166), .A(n7117), .B(n7115), .S(n7168), .CO(n7169) );
  HA1 U6782 ( .A(n5864), .B(n5379), .S(n7170), .CO(n7171) );
  FA1A U6783 ( .CI(n5315), .A(n3715), .B(n4483), .S(n7172), .CO(n7173) );
  FA1A U6784 ( .CI(n3843), .A(n3779), .B(n4611), .S(n7174), .CO(n7175) );
  FA1A U6785 ( .CI(n3971), .A(n3907), .B(n4739), .S(n7176), .CO(n7177) );
  FA1A U6786 ( .CI(n5251), .A(n4035), .B(n4867), .S(n7178), .CO(n7179) );
  FA1A U6787 ( .CI(n4099), .A(n5187), .B(n4803), .S(n7180), .CO(n7181) );
  FA1A U6788 ( .CI(n5059), .A(n5123), .B(n4163), .S(n7182), .CO(n7183) );
  FA1A U6789 ( .CI(n4931), .A(n4995), .B(n4227), .S(n7184), .CO(n7185) );
  FA1A U6790 ( .CI(n4547), .A(n4675), .B(n4291), .S(n7186), .CO(n7187) );
  FA1A U6791 ( .CI(n7170), .A(n4355), .B(n4419), .S(n7188), .CO(n7189) );
  FA1A U6792 ( .CI(n7188), .A(n7186), .B(n7121), .S(n7190), .CO(n7191) );
  FA1A U6793 ( .CI(n7182), .A(n7184), .B(n7123), .S(n7192), .CO(n7193) );
  FA1A U6794 ( .CI(n7172), .A(n7180), .B(n7133), .S(n7194), .CO(n7195) );
  FA1A U6795 ( .CI(n7174), .A(n7176), .B(n7125), .S(n7196), .CO(n7197) );
  FA1A U6796 ( .CI(n7178), .A(n7137), .B(n7127), .S(n7198), .CO(n7199) );
  FA1A U6797 ( .CI(n7135), .A(n7131), .B(n7129), .S(n7200), .CO(n7201) );
  FA1A U6798 ( .CI(n7200), .A(n7190), .B(n7139), .S(n7202), .CO(n7203) );
  FA1A U6799 ( .CI(n7194), .A(n7198), .B(n7147), .S(n7204), .CO(n7205) );
  FA1A U6800 ( .CI(n7196), .A(n7192), .B(n7141), .S(n7206), .CO(n7207) );
  FA1A U6801 ( .CI(n7145), .A(n7149), .B(n7143), .S(n7208), .CO(n7209) );
  FA1A U6802 ( .CI(n7208), .A(n7202), .B(n7151), .S(n7210), .CO(n7211) );
  FA1A U6803 ( .CI(n7204), .A(n7206), .B(n7153), .S(n7212), .CO(n7213) );
  FA1A U6804 ( .CI(n7159), .A(n7157), .B(n7155), .S(n7214), .CO(n7215) );
  FA1A U6805 ( .CI(n7214), .A(n7161), .B(n7210), .S(n7216), .CO(n7217) );
  FA1A U6806 ( .CI(n7216), .A(n7163), .B(n7212), .S(n7218), .CO(n7219) );
  FA1A U6807 ( .CI(n7218), .A(n7167), .B(n7165), .S(n7220), .CO(n7221) );
  FA1A U6808 ( .CI(n5380), .A(n5316), .B(n10872), .S(n7222), .CO(n7223) );
  FA1A U6809 ( .CI(n7171), .A(n5252), .B(n4548), .S(n7224), .CO(n7225) );
  FA1A U6810 ( .CI(n3780), .A(n3716), .B(n4484), .S(n7226), .CO(n7227) );
  FA1A U6811 ( .CI(n5188), .A(n3844), .B(n4612), .S(n7228), .CO(n7229) );
  FA1A U6812 ( .CI(n3908), .A(n5124), .B(n4676), .S(n7230), .CO(n7231) );
  FA1A U6813 ( .CI(n3972), .A(n5060), .B(n4996), .S(n7232), .CO(n7233) );
  FA1A U6814 ( .CI(n4868), .A(n4932), .B(n4036), .S(n7234), .CO(n7235) );
  FA1A U6815 ( .CI(n4740), .A(n4804), .B(n4100), .S(n7236), .CO(n7237) );
  FA1A U6816 ( .CI(n4356), .A(n4420), .B(n4164), .S(n7238), .CO(n7239) );
  FA1A U6817 ( .CI(n7222), .A(n4228), .B(n4292), .S(n7240), .CO(n7241) );
  FA1A U6818 ( .CI(n7240), .A(n7238), .B(n7185), .S(n7242), .CO(n7243) );
  FA1A U6819 ( .CI(n7189), .A(n7236), .B(n7173), .S(n7244), .CO(n7245) );
  FA1A U6820 ( .CI(n7232), .A(n7234), .B(n7183), .S(n7246), .CO(n7247) );
  FA1A U6821 ( .CI(n7224), .A(n7230), .B(n7181), .S(n7248), .CO(n7249) );
  FA1A U6822 ( .CI(n7226), .A(n7228), .B(n7175), .S(n7250), .CO(n7251) );
  FA1A U6823 ( .CI(n7179), .A(n7187), .B(n7177), .S(n7252), .CO(n7253) );
  FA1A U6824 ( .CI(n7250), .A(n7252), .B(n7191), .S(n7254), .CO(n7255) );
  FA1A U6825 ( .CI(n7244), .A(n7248), .B(n7199), .S(n7256), .CO(n7257) );
  FA1A U6826 ( .CI(n7246), .A(n7242), .B(n7193), .S(n7258), .CO(n7259) );
  FA1A U6827 ( .CI(n7197), .A(n7201), .B(n7195), .S(n7260), .CO(n7261) );
  FA1A U6828 ( .CI(n7258), .A(n7260), .B(n7203), .S(n7262), .CO(n7263) );
  FA1A U6829 ( .CI(n7256), .A(n7205), .B(n7254), .S(n7264), .CO(n7265) );
  FA1A U6830 ( .CI(n7211), .A(n7209), .B(n7207), .S(n7266), .CO(n7267) );
  FA1A U6831 ( .CI(n7266), .A(n7213), .B(n7262), .S(n7268), .CO(n7269) );
  FA1A U6832 ( .CI(n7268), .A(n7215), .B(n7264), .S(n7270), .CO(n7271) );
  FA1A U6833 ( .CI(n7270), .A(n7219), .B(n7217), .S(n7272), .CO(n7273) );
  HA1 U6834 ( .A(n5865), .B(n5445), .S(n7274), .CO(n7275) );
  FA1A U6835 ( .CI(n5317), .A(n5381), .B(n4485), .S(n7276), .CO(n7277) );
  FA1A U6836 ( .CI(n3717), .A(n5253), .B(n4613), .S(n7278), .CO(n7279) );
  FA1A U6837 ( .CI(n3781), .A(n5189), .B(n4549), .S(n7280), .CO(n7281) );
  FA1A U6838 ( .CI(n5061), .A(n5125), .B(n4677), .S(n7282), .CO(n7283) );
  FA1A U6839 ( .CI(n3909), .A(n3845), .B(n4421), .S(n7284), .CO(n7285) );
  FA1A U6840 ( .CI(n4933), .A(n4997), .B(n3973), .S(n7286), .CO(n7287) );
  FA1A U6841 ( .CI(n4805), .A(n4869), .B(n4037), .S(n7288), .CO(n7289) );
  FA1A U6842 ( .CI(n4357), .A(n4741), .B(n4101), .S(n7290), .CO(n7291) );
  FA1A U6843 ( .CI(n4293), .A(n4229), .B(n4165), .S(n7292), .CO(n7293) );
  FA1A U6844 ( .CI(n7292), .A(n7223), .B(n7274), .S(n7294), .CO(n7295) );
  FA1A U6845 ( .CI(n7241), .A(n7290), .B(n7237), .S(n7296), .CO(n7297) );
  FA1A U6846 ( .CI(n7286), .A(n7288), .B(n7235), .S(n7298), .CO(n7299) );
  FA1A U6847 ( .CI(n7282), .A(n7284), .B(n7233), .S(n7300), .CO(n7301) );
  FA1A U6848 ( .CI(n7280), .A(n7276), .B(n7225), .S(n7302), .CO(n7303) );
  FA1A U6849 ( .CI(n7278), .A(n7239), .B(n7227), .S(n7304), .CO(n7305) );
  FA1A U6850 ( .CI(n7294), .A(n7231), .B(n7229), .S(n7306), .CO(n7307) );
  FA1A U6851 ( .CI(n7306), .A(n7304), .B(n7251), .S(n7308), .CO(n7309) );
  FA1A U6852 ( .CI(n7300), .A(n7302), .B(n7249), .S(n7310), .CO(n7311) );
  FA1A U6853 ( .CI(n7298), .A(n7296), .B(n7243), .S(n7312), .CO(n7313) );
  FA1A U6854 ( .CI(n7247), .A(n7253), .B(n7245), .S(n7314), .CO(n7315) );
  FA1A U6855 ( .CI(n7312), .A(n7314), .B(n7255), .S(n7316), .CO(n7317) );
  FA1A U6856 ( .CI(n7308), .A(n7310), .B(n7257), .S(n7318), .CO(n7319) );
  FA1A U6857 ( .CI(n7263), .A(n7261), .B(n7259), .S(n7320), .CO(n7321) );
  FA1A U6858 ( .CI(n7267), .A(n7318), .B(n7265), .S(n7322), .CO(n7323) );
  FA1A U6859 ( .CI(n7269), .A(n7320), .B(n7316), .S(n7324), .CO(n7325) );
  FA1A U6860 ( .CI(n7324), .A(n7271), .B(n7322), .S(n7326), .CO(n7327) );
  FA1A U6861 ( .CI(n5446), .A(n5382), .B(n10871), .S(n7328), .CO(n7329) );
  FA1A U6862 ( .CI(n7275), .A(n5318), .B(n4614), .S(n7330), .CO(n7331) );
  FA1A U6863 ( .CI(n3782), .A(n3718), .B(n4486), .S(n7332), .CO(n7333) );
  FA1A U6864 ( .CI(n3846), .A(n5254), .B(n4678), .S(n7334), .CO(n7335) );
  FA1A U6865 ( .CI(n5190), .A(n3910), .B(n4742), .S(n7336), .CO(n7337) );
  FA1A U6866 ( .CI(n3974), .A(n5126), .B(n4550), .S(n7338), .CO(n7339) );
  FA1A U6867 ( .CI(n4998), .A(n5062), .B(n4038), .S(n7340), .CO(n7341) );
  FA1A U6868 ( .CI(n4870), .A(n4934), .B(n4102), .S(n7342), .CO(n7343) );
  FA1A U6869 ( .CI(n4422), .A(n4806), .B(n4166), .S(n7344), .CO(n7345) );
  FA1A U6870 ( .CI(n4358), .A(n4294), .B(n4230), .S(n7346), .CO(n7347) );
  FA1A U6871 ( .CI(n7346), .A(n7293), .B(n7328), .S(n7348), .CO(n7349) );
  FA1A U6872 ( .CI(n7330), .A(n7344), .B(n7289), .S(n7350), .CO(n7351) );
  FA1A U6873 ( .CI(n7340), .A(n7342), .B(n7277), .S(n7352), .CO(n7353) );
  FA1A U6874 ( .CI(n7334), .A(n7338), .B(n7285), .S(n7354), .CO(n7355) );
  FA1A U6875 ( .CI(n7332), .A(n7336), .B(n7279), .S(n7356), .CO(n7357) );
  FA1A U6876 ( .CI(n7287), .A(n7291), .B(n7281), .S(n7358), .CO(n7359) );
  FA1A U6877 ( .CI(n7348), .A(n7295), .B(n7283), .S(n7360), .CO(n7361) );
  FA1A U6878 ( .CI(n7307), .A(n7358), .B(n7303), .S(n7362), .CO(n7363) );
  FA1A U6879 ( .CI(n7354), .A(n7356), .B(n7301), .S(n7364), .CO(n7365) );
  FA1A U6880 ( .CI(n7352), .A(n7350), .B(n7297), .S(n7366), .CO(n7367) );
  FA1A U6881 ( .CI(n7360), .A(n7305), .B(n7299), .S(n7368), .CO(n7369) );
  FA1A U6882 ( .CI(n7368), .A(n7366), .B(n7309), .S(n7370), .CO(n7371) );
  FA1A U6883 ( .CI(n7362), .A(n7364), .B(n7311), .S(n7372), .CO(n7373) );
  FA1A U6884 ( .CI(n7317), .A(n7315), .B(n7313), .S(n7374), .CO(n7375) );
  FA1A U6885 ( .CI(n7372), .A(n7370), .B(n7319), .S(n7376), .CO(n7377) );
  FA1A U6886 ( .CI(n7323), .A(n7374), .B(n7321), .S(n7378), .CO(n7379) );
  FA1A U6887 ( .CI(n7378), .A(n7325), .B(n7376), .S(n7380), .CO(n7381) );
  HA1 U6888 ( .A(n5866), .B(n5511), .S(n7382), .CO(n7383) );
  FA1A U6889 ( .CI(n3783), .A(n3719), .B(n4551), .S(n7384), .CO(n7385) );
  FA1A U6890 ( .CI(n5383), .A(n5447), .B(n4743), .S(n7386), .CO(n7387) );
  FA1A U6891 ( .CI(n5255), .A(n5319), .B(n4679), .S(n7388), .CO(n7389) );
  FA1A U6892 ( .CI(n5127), .A(n5191), .B(n4487), .S(n7390), .CO(n7391) );
  FA1A U6893 ( .CI(n3847), .A(n5063), .B(n4423), .S(n7392), .CO(n7393) );
  FA1A U6894 ( .CI(n4935), .A(n4999), .B(n3911), .S(n7394), .CO(n7395) );
  FA1A U6895 ( .CI(n4807), .A(n4871), .B(n3975), .S(n7396), .CO(n7397) );
  FA1A U6896 ( .CI(n4359), .A(n4615), .B(n4039), .S(n7398), .CO(n7399) );
  FA1A U6897 ( .CI(n4295), .A(n4167), .B(n4103), .S(n7400), .CO(n7401) );
  FA1A U6898 ( .CI(n7329), .A(n7382), .B(n4231), .S(n7402), .CO(n7403) );
  FA1A U6899 ( .CI(n7398), .A(n7400), .B(n7345), .S(n7404), .CO(n7405) );
  FA1A U6900 ( .CI(n7394), .A(n7396), .B(n7341), .S(n7406), .CO(n7407) );
  FA1A U6901 ( .CI(n7390), .A(n7392), .B(n7331), .S(n7408), .CO(n7409) );
  FA1A U6902 ( .CI(n7388), .A(n7384), .B(n7333), .S(n7410), .CO(n7411) );
  FA1A U6903 ( .CI(n7386), .A(n7347), .B(n7335), .S(n7412), .CO(n7413) );
  FA1A U6904 ( .CI(n7339), .A(n7343), .B(n7337), .S(n7414), .CO(n7415) );
  FA1A U6905 ( .CI(n7414), .A(n7349), .B(n7402), .S(n7416), .CO(n7417) );
  FA1A U6906 ( .CI(n7410), .A(n7412), .B(n7357), .S(n7418), .CO(n7419) );
  FA1A U6907 ( .CI(n7404), .A(n7408), .B(n7355), .S(n7420), .CO(n7421) );
  FA1A U6908 ( .CI(n7406), .A(n7359), .B(n7351), .S(n7422), .CO(n7423) );
  FA1A U6909 ( .CI(n7361), .A(n7416), .B(n7353), .S(n7424), .CO(n7425) );
  FA1A U6910 ( .CI(n7369), .A(n7422), .B(n7363), .S(n7426), .CO(n7427) );
  FA1A U6911 ( .CI(n7420), .A(n7418), .B(n7365), .S(n7428), .CO(n7429) );
  FA1A U6912 ( .CI(n7371), .A(n7424), .B(n7367), .S(n7430), .CO(n7431) );
  FA1A U6913 ( .CI(n7428), .A(n7426), .B(n7373), .S(n7432), .CO(n7433) );
  FA1A U6914 ( .CI(n7377), .A(n7430), .B(n7375), .S(n7434), .CO(n7435) );
  FA1A U6915 ( .CI(n7434), .A(n7379), .B(n7432), .S(n7436), .CO(n7437) );
  FA1A U6916 ( .CI(n5512), .A(n5448), .B(n10870), .S(n7438), .CO(n7439) );
  FA1A U6917 ( .CI(n7383), .A(n3720), .B(n4616), .S(n7440), .CO(n7441) );
  FA1A U6918 ( .CI(n3784), .A(n5384), .B(n4680), .S(n7442), .CO(n7443) );
  FA1A U6919 ( .CI(n3912), .A(n3848), .B(n4744), .S(n7444), .CO(n7445) );
  FA1A U6920 ( .CI(n5256), .A(n5320), .B(n4808), .S(n7446), .CO(n7447) );
  FA1A U6921 ( .CI(n5192), .A(n3976), .B(n4552), .S(n7448), .CO(n7449) );
  FA1A U6922 ( .CI(n5064), .A(n5128), .B(n4040), .S(n7450), .CO(n7451) );
  FA1A U6923 ( .CI(n4936), .A(n5000), .B(n4104), .S(n7452), .CO(n7453) );
  FA1A U6924 ( .CI(n4488), .A(n4872), .B(n4168), .S(n7454), .CO(n7455) );
  FA1A U6925 ( .CI(n4296), .A(n4424), .B(n4232), .S(n7456), .CO(n7457) );
  FA1A U6926 ( .CI(n7385), .A(n7438), .B(n4360), .S(n7458), .CO(n7459) );
  FA1A U6927 ( .CI(n7454), .A(n7456), .B(n7399), .S(n7460), .CO(n7461) );
  FA1A U6928 ( .CI(n7450), .A(n7452), .B(n7397), .S(n7462), .CO(n7463) );
  FA1A U6929 ( .CI(n7446), .A(n7448), .B(n7387), .S(n7464), .CO(n7465) );
  FA1A U6930 ( .CI(n7440), .A(n7442), .B(n7389), .S(n7466), .CO(n7467) );
  FA1A U6931 ( .CI(n7444), .A(n7401), .B(n7391), .S(n7468), .CO(n7469) );
  FA1A U6932 ( .CI(n7403), .A(n7395), .B(n7393), .S(n7470), .CO(n7471) );
  FA1A U6933 ( .CI(n7470), .A(n7413), .B(n7458), .S(n7472), .CO(n7473) );
  FA1A U6934 ( .CI(n7466), .A(n7468), .B(n7411), .S(n7474), .CO(n7475) );
  FA1A U6935 ( .CI(n7460), .A(n7464), .B(n7409), .S(n7476), .CO(n7477) );
  FA1A U6936 ( .CI(n7462), .A(n7415), .B(n7405), .S(n7478), .CO(n7479) );
  FA1A U6937 ( .CI(n7417), .A(n7472), .B(n7407), .S(n7480), .CO(n7481) );
  FA1A U6938 ( .CI(n7476), .A(n7478), .B(n7419), .S(n7482), .CO(n7483) );
  FA1A U6939 ( .CI(n7474), .A(n7423), .B(n7421), .S(n7484), .CO(n7485) );
  FA1A U6940 ( .CI(n7484), .A(n7425), .B(n7480), .S(n7486), .CO(n7487) );
  FA1A U6941 ( .CI(n7482), .A(n7429), .B(n7427), .S(n7488), .CO(n7489) );
  FA1A U6942 ( .CI(n7488), .A(n7486), .B(n7431), .S(n7490), .CO(n7491) );
  FA1A U6943 ( .CI(n7490), .A(n7435), .B(n7433), .S(n7492), .CO(n7493) );
  HA1 U6944 ( .A(n5867), .B(n5577), .S(n7494), .CO(n7495) );
  FA1A U6945 ( .CI(n3721), .A(n5513), .B(n4553), .S(n7496), .CO(n7497) );
  FA1A U6946 ( .CI(n3785), .A(n5449), .B(n4745), .S(n7498), .CO(n7499) );
  FA1A U6947 ( .CI(n5385), .A(n3849), .B(n4809), .S(n7500), .CO(n7501) );
  FA1A U6948 ( .CI(n3977), .A(n3913), .B(n4681), .S(n7502), .CO(n7503) );
  FA1A U6949 ( .CI(n4041), .A(n5321), .B(n4937), .S(n7504), .CO(n7505) );
  FA1A U6950 ( .CI(n5129), .A(n5193), .B(n5257), .S(n7506), .CO(n7507) );
  FA1A U6951 ( .CI(n5001), .A(n5065), .B(n4105), .S(n7508), .CO(n7509) );
  FA1A U6952 ( .CI(n4617), .A(n4873), .B(n4169), .S(n7510), .CO(n7511) );
  FA1A U6953 ( .CI(n4425), .A(n4489), .B(n4233), .S(n7512), .CO(n7513) );
  FA1A U6954 ( .CI(n7494), .A(n4361), .B(n4297), .S(n7514), .CO(n7515) );
  FA1A U6955 ( .CI(n7514), .A(n7512), .B(n7439), .S(n7516), .CO(n7517) );
  FA1A U6956 ( .CI(n7498), .A(n7510), .B(n7453), .S(n7518), .CO(n7519) );
  FA1A U6957 ( .CI(n7506), .A(n7508), .B(n7441), .S(n7520), .CO(n7521) );
  FA1A U6958 ( .CI(n7500), .A(n7504), .B(n7443), .S(n7522), .CO(n7523) );
  FA1A U6959 ( .CI(n7496), .A(n7502), .B(n7445), .S(n7524), .CO(n7525) );
  FA1A U6960 ( .CI(n7455), .A(n7457), .B(n7447), .S(n7526), .CO(n7527) );
  FA1A U6961 ( .CI(n7459), .A(n7451), .B(n7449), .S(n7528), .CO(n7529) );
  FA1A U6962 ( .CI(n7528), .A(n7526), .B(n7516), .S(n7530), .CO(n7531) );
  FA1A U6963 ( .CI(n7471), .A(n7524), .B(n7467), .S(n7532), .CO(n7533) );
  FA1A U6964 ( .CI(n7518), .A(n7522), .B(n7465), .S(n7534), .CO(n7535) );
  FA1A U6965 ( .CI(n7520), .A(n7469), .B(n7461), .S(n7536), .CO(n7537) );
  FA1A U6966 ( .CI(n7530), .A(n7473), .B(n7463), .S(n7538), .CO(n7539) );
  FA1A U6967 ( .CI(n7534), .A(n7536), .B(n7475), .S(n7540), .CO(n7541) );
  FA1A U6968 ( .CI(n7532), .A(n7479), .B(n7477), .S(n7542), .CO(n7543) );
  FA1A U6969 ( .CI(n7542), .A(n7538), .B(n7481), .S(n7544), .CO(n7545) );
  FA1A U6970 ( .CI(n7540), .A(n7485), .B(n7483), .S(n7546), .CO(n7547) );
  FA1A U6971 ( .CI(n7546), .A(n7544), .B(n7487), .S(n7548), .CO(n7549) );
  FA1A U6972 ( .CI(n7548), .A(n7491), .B(n7489), .S(n7550), .CO(n7551) );
  FA1A U6973 ( .CI(n5578), .A(n5514), .B(n10869), .S(n7552), .CO(n7553) );
  FA1A U6974 ( .CI(n7495), .A(n3722), .B(n4682), .S(n7554), .CO(n7555) );
  FA1A U6975 ( .CI(n3786), .A(n5450), .B(n4746), .S(n7556), .CO(n7557) );
  FA1A U6976 ( .CI(n3914), .A(n3850), .B(n4618), .S(n7558), .CO(n7559) );
  FA1A U6977 ( .CI(n4042), .A(n3978), .B(n4810), .S(n7560), .CO(n7561) );
  FA1A U6978 ( .CI(n5386), .A(n4106), .B(n4938), .S(n7562), .CO(n7563) );
  FA1A U6979 ( .CI(n5194), .A(n5258), .B(n5322), .S(n7564), .CO(n7565) );
  FA1A U6980 ( .CI(n5066), .A(n5130), .B(n4170), .S(n7566), .CO(n7567) );
  FA1A U6981 ( .CI(n4874), .A(n5002), .B(n4234), .S(n7568), .CO(n7569) );
  FA1A U6982 ( .CI(n4490), .A(n4554), .B(n4298), .S(n7570), .CO(n7571) );
  FA1A U6983 ( .CI(n7552), .A(n4426), .B(n4362), .S(n7572), .CO(n7573) );
  FA1A U6984 ( .CI(n7572), .A(n7570), .B(n7511), .S(n7574), .CO(n7575) );
  FA1A U6985 ( .CI(n7515), .A(n7568), .B(n7509), .S(n7576), .CO(n7577) );
  FA1A U6986 ( .CI(n7564), .A(n7566), .B(n7507), .S(n7578), .CO(n7579) );
  FA1A U6987 ( .CI(n7560), .A(n7562), .B(n7497), .S(n7580), .CO(n7581) );
  FA1A U6988 ( .CI(n7558), .A(n7556), .B(n7505), .S(n7582), .CO(n7583) );
  FA1A U6989 ( .CI(n7554), .A(n7513), .B(n7499), .S(n7584), .CO(n7585) );
  FA1A U6990 ( .CI(n7517), .A(n7503), .B(n7501), .S(n7586), .CO(n7587) );
  FA1A U6991 ( .CI(n7529), .A(n7584), .B(n7527), .S(n7588), .CO(n7589) );
  FA1A U6992 ( .CI(n7580), .A(n7582), .B(n7525), .S(n7590), .CO(n7591) );
  FA1A U6993 ( .CI(n7578), .A(n7574), .B(n7519), .S(n7592), .CO(n7593) );
  FA1A U6994 ( .CI(n7576), .A(n7521), .B(n7523), .S(n7594), .CO(n7595) );
  FA1A U6995 ( .CI(n7533), .A(n7531), .B(n7586), .S(n7596), .CO(n7597) );
  FA1A U6996 ( .CI(n7592), .A(n7588), .B(n7535), .S(n7598), .CO(n7599) );
  FA1A U6997 ( .CI(n7594), .A(n7590), .B(n7537), .S(n7600), .CO(n7601) );
  FA1A U6998 ( .CI(n7600), .A(n7539), .B(n7596), .S(n7602), .CO(n7603) );
  FA1A U6999 ( .CI(n7598), .A(n7543), .B(n7541), .S(n7604), .CO(n7605) );
  FA1A U7000 ( .CI(n7604), .A(n7602), .B(n7545), .S(n7606), .CO(n7607) );
  FA1A U7001 ( .CI(n7606), .A(n7549), .B(n7547), .S(n7608), .CO(n7609) );
  HA1 U7002 ( .A(n5868), .B(n5643), .S(n7610), .CO(n7611) );
  FA1A U7003 ( .CI(n5579), .A(n3723), .B(n4619), .S(n7612), .CO(n7613) );
  FA1A U7004 ( .CI(n5515), .A(n3787), .B(n4747), .S(n7614), .CO(n7615) );
  FA1A U7005 ( .CI(n5451), .A(n3851), .B(n4811), .S(n7616), .CO(n7617) );
  FA1A U7006 ( .CI(n3915), .A(n5387), .B(n4683), .S(n7618), .CO(n7619) );
  FA1A U7007 ( .CI(n5323), .A(n3979), .B(n4875), .S(n7620), .CO(n7621) );
  FA1A U7008 ( .CI(n4107), .A(n4043), .B(n5259), .S(n7622), .CO(n7623) );
  FA1A U7009 ( .CI(n5131), .A(n5195), .B(n4171), .S(n7624), .CO(n7625) );
  FA1A U7010 ( .CI(n5003), .A(n5067), .B(n4235), .S(n7626), .CO(n7627) );
  FA1A U7011 ( .CI(n4555), .A(n4939), .B(n4299), .S(n7628), .CO(n7629) );
  FA1A U7012 ( .CI(n4427), .A(n4491), .B(n4363), .S(n7630), .CO(n7631) );
  FA1A U7013 ( .CI(n7630), .A(n7553), .B(n7610), .S(n7632), .CO(n7633) );
  FA1A U7014 ( .CI(n7573), .A(n7628), .B(n7569), .S(n7634), .CO(n7635) );
  FA1A U7015 ( .CI(n7624), .A(n7626), .B(n7567), .S(n7636), .CO(n7637) );
  FA1A U7016 ( .CI(n7612), .A(n7622), .B(n7565), .S(n7638), .CO(n7639) );
  FA1A U7017 ( .CI(n7616), .A(n7614), .B(n7555), .S(n7640), .CO(n7641) );
  FA1A U7018 ( .CI(n7618), .A(n7620), .B(n7563), .S(n7642), .CO(n7643) );
  FA1A U7019 ( .CI(n7561), .A(n7571), .B(n7557), .S(n7644), .CO(n7645) );
  FA1A U7020 ( .CI(n7575), .A(n7632), .B(n7559), .S(n7646), .CO(n7647) );
  FA1A U7021 ( .CI(n7642), .A(n7644), .B(n7585), .S(n7648), .CO(n7649) );
  FA1A U7022 ( .CI(n7638), .A(n7640), .B(n7581), .S(n7650), .CO(n7651) );
  FA1A U7023 ( .CI(n7634), .A(n7636), .B(n7577), .S(n7652), .CO(n7653) );
  FA1A U7024 ( .CI(n7587), .A(n7583), .B(n7579), .S(n7654), .CO(n7655) );
  FA1A U7025 ( .CI(n7654), .A(n7589), .B(n7646), .S(n7656), .CO(n7657) );
  FA1A U7026 ( .CI(n7650), .A(n7652), .B(n7591), .S(n7658), .CO(n7659) );
  FA1A U7027 ( .CI(n7648), .A(n7595), .B(n7593), .S(n7660), .CO(n7661) );
  FA1A U7028 ( .CI(n7660), .A(n7601), .B(n7656), .S(n7662), .CO(n7663) );
  FA1A U7029 ( .CI(n7658), .A(n7599), .B(n7597), .S(n7664), .CO(n7665) );
  FA1A U7030 ( .CI(n7605), .A(n7664), .B(n7603), .S(n7666), .CO(n7667) );
  FA1A U7031 ( .CI(n7666), .A(n7607), .B(n7662), .S(n7668), .CO(n7669) );
  FA1A U7032 ( .CI(n5644), .A(n5580), .B(n10868), .S(n7670), .CO(n7671) );
  FA1A U7033 ( .CI(n7611), .A(n3724), .B(n4684), .S(n7672), .CO(n7673) );
  FA1A U7034 ( .CI(n5452), .A(n5516), .B(n4748), .S(n7674), .CO(n7675) );
  FA1A U7035 ( .CI(n5388), .A(n3788), .B(n4620), .S(n7676), .CO(n7677) );
  FA1A U7036 ( .CI(n3916), .A(n3852), .B(n4556), .S(n7678), .CO(n7679) );
  FA1A U7037 ( .CI(n3980), .A(n5324), .B(n4876), .S(n7680), .CO(n7681) );
  FA1A U7038 ( .CI(n4108), .A(n4044), .B(n5260), .S(n7682), .CO(n7683) );
  FA1A U7039 ( .CI(n5132), .A(n5196), .B(n4172), .S(n7684), .CO(n7685) );
  FA1A U7040 ( .CI(n5004), .A(n5068), .B(n4236), .S(n7686), .CO(n7687) );
  FA1A U7041 ( .CI(n4812), .A(n4940), .B(n4300), .S(n7688), .CO(n7689) );
  FA1A U7042 ( .CI(n4428), .A(n4492), .B(n4364), .S(n7690), .CO(n7691) );
  FA1A U7043 ( .CI(n7690), .A(n7631), .B(n7670), .S(n7692), .CO(n7693) );
  FA1A U7044 ( .CI(n7686), .A(n7688), .B(n7627), .S(n7694), .CO(n7695) );
  FA1A U7045 ( .CI(n7682), .A(n7684), .B(n7623), .S(n7696), .CO(n7697) );
  FA1A U7046 ( .CI(n7674), .A(n7672), .B(n7613), .S(n7698), .CO(n7699) );
  FA1A U7047 ( .CI(n7678), .A(n7676), .B(n7615), .S(n7700), .CO(n7701) );
  FA1A U7048 ( .CI(n7680), .A(n7629), .B(n7617), .S(n7702), .CO(n7703) );
  FA1A U7049 ( .CI(n7621), .A(n7625), .B(n7619), .S(n7704), .CO(n7705) );
  FA1A U7050 ( .CI(n7702), .A(n7704), .B(n7633), .S(n7706), .CO(n7707) );
  FA1A U7051 ( .CI(n7694), .A(n7700), .B(n7692), .S(n7708), .CO(n7709) );
  FA1A U7052 ( .CI(n7698), .A(n7696), .B(n7635), .S(n7710), .CO(n7711) );
  FA1A U7053 ( .CI(n7643), .A(n7645), .B(n7637), .S(n7712), .CO(n7713) );
  FA1A U7054 ( .CI(n7647), .A(n7641), .B(n7639), .S(n7714), .CO(n7715) );
  FA1A U7055 ( .CI(n7714), .A(n7655), .B(n7706), .S(n7716), .CO(n7717) );
  FA1A U7056 ( .CI(n7710), .A(n7712), .B(n7708), .S(n7718), .CO(n7719) );
  FA1A U7057 ( .CI(n7651), .A(n7653), .B(n7649), .S(n7720), .CO(n7721) );
  FA1A U7058 ( .CI(n7720), .A(n7661), .B(n7716), .S(n7722), .CO(n7723) );
  FA1A U7059 ( .CI(n7659), .A(n7657), .B(n7718), .S(n7724), .CO(n7725) );
  FA1A U7060 ( .CI(n7663), .A(n7665), .B(n7722), .S(n7726), .CO(n7727) );
  FA1A U7061 ( .CI(n7726), .A(n7667), .B(n7724), .S(n7728), .CO(n7729) );
  HA1 U7062 ( .A(n5869), .B(n5709), .S(n7730), .CO(n7731) );
  FA1A U7063 ( .CI(n3725), .A(n5645), .B(n4621), .S(n7732), .CO(n7733) );
  FA1A U7064 ( .CI(n3789), .A(n5581), .B(n4813), .S(n7734), .CO(n7735) );
  FA1A U7065 ( .CI(n5517), .A(n3853), .B(n4877), .S(n7736), .CO(n7737) );
  FA1A U7066 ( .CI(n5389), .A(n5453), .B(n4749), .S(n7738), .CO(n7739) );
  FA1A U7067 ( .CI(n3981), .A(n3917), .B(n4685), .S(n7740), .CO(n7741) );
  FA1A U7068 ( .CI(n4109), .A(n4045), .B(n5005), .S(n7742), .CO(n7743) );
  FA1A U7069 ( .CI(n5261), .A(n5325), .B(n4173), .S(n7744), .CO(n7745) );
  FA1A U7070 ( .CI(n5133), .A(n5197), .B(n4237), .S(n7746), .CO(n7747) );
  FA1A U7071 ( .CI(n4941), .A(n5069), .B(n4301), .S(n7748), .CO(n7749) );
  FA1A U7072 ( .CI(n4493), .A(n4557), .B(n4365), .S(n7750), .CO(n7751) );
  FA1A U7073 ( .CI(n7671), .A(n7730), .B(n4429), .S(n7752), .CO(n7753) );
  FA1A U7074 ( .CI(n7748), .A(n7750), .B(n7689), .S(n7754), .CO(n7755) );
  FA1A U7075 ( .CI(n7744), .A(n7746), .B(n7685), .S(n7756), .CO(n7757) );
  FA1A U7076 ( .CI(n7732), .A(n7742), .B(n7683), .S(n7758), .CO(n7759) );
  FA1A U7077 ( .CI(n7740), .A(n7736), .B(n7673), .S(n7760), .CO(n7761) );
  FA1A U7078 ( .CI(n7738), .A(n7734), .B(n7675), .S(n7762), .CO(n7763) );
  FA1A U7079 ( .CI(n7687), .A(n7691), .B(n7677), .S(n7764), .CO(n7765) );
  FA1A U7080 ( .CI(n7752), .A(n7681), .B(n7679), .S(n7766), .CO(n7767) );
  FA1A U7081 ( .CI(n7766), .A(n7764), .B(n7693), .S(n7768), .CO(n7769) );
  FA1A U7082 ( .CI(n7760), .A(n7762), .B(n7695), .S(n7770), .CO(n7771) );
  FA1A U7083 ( .CI(n7754), .A(n7758), .B(n7701), .S(n7772), .CO(n7773) );
  FA1A U7084 ( .CI(n7756), .A(n7705), .B(n7697), .S(n7774), .CO(n7775) );
  FA1A U7085 ( .CI(n7707), .A(n7703), .B(n7699), .S(n7776), .CO(n7777) );
  FA1A U7086 ( .CI(n7715), .A(n7774), .B(n7709), .S(n7778), .CO(n7779) );
  FA1A U7087 ( .CI(n7772), .A(n7770), .B(n7768), .S(n7780), .CO(n7781) );
  FA1A U7088 ( .CI(n7776), .A(n7713), .B(n7711), .S(n7782), .CO(n7783) );
  FA1A U7089 ( .CI(n7782), .A(n7721), .B(n7719), .S(n7784), .CO(n7785) );
  FA1A U7090 ( .CI(n7780), .A(n7778), .B(n7717), .S(n7786), .CO(n7787) );
  FA1A U7091 ( .CI(n7786), .A(n7784), .B(n7725), .S(n7788), .CO(n7789) );
  FA1A U7092 ( .CI(n7788), .A(n7727), .B(n7723), .S(n7790), .CO(n7791) );
  FA1A U7093 ( .CI(n3726), .A(n5646), .B(n10867), .S(n7792), .CO(n7793) );
  FA1A U7094 ( .CI(n7731), .A(n3790), .B(n4814), .S(n7794), .CO(n7795) );
  FA1A U7095 ( .CI(n3918), .A(n3854), .B(n4878), .S(n7796), .CO(n7797) );
  FA1A U7096 ( .CI(n4046), .A(n3982), .B(n4942), .S(n7798), .CO(n7799) );
  FA1A U7097 ( .CI(n5710), .A(n4110), .B(n5070), .S(n7800), .CO(n7801) );
  FA1A U7098 ( .CI(n4238), .A(n4174), .B(n5006), .S(n7802), .CO(n7803) );
  FA1A U7099 ( .CI(n4366), .A(n4302), .B(n5518), .S(n7804), .CO(n7805) );
  FA1A U7100 ( .CI(n5454), .A(n5582), .B(n4430), .S(n7806), .CO(n7807) );
  FA1A U7101 ( .CI(n5326), .A(n5390), .B(n4494), .S(n7808), .CO(n7809) );
  FA1A U7102 ( .CI(n5198), .A(n5262), .B(n4558), .S(n7810), .CO(n7811) );
  FA1A U7103 ( .CI(n4750), .A(n5134), .B(n4622), .S(n7812), .CO(n7813) );
  FA1A U7104 ( .CI(n7733), .A(n7792), .B(n4686), .S(n7814), .CO(n7815) );
  FA1A U7105 ( .CI(n7810), .A(n7812), .B(n7749), .S(n7816), .CO(n7817) );
  FA1A U7106 ( .CI(n7806), .A(n7808), .B(n7747), .S(n7818), .CO(n7819) );
  FA1A U7107 ( .CI(n7794), .A(n7804), .B(n7745), .S(n7820), .CO(n7821) );
  FA1A U7108 ( .CI(n7802), .A(n7796), .B(n7735), .S(n7822), .CO(n7823) );
  FA1A U7109 ( .CI(n7800), .A(n7798), .B(n7737), .S(n7824), .CO(n7825) );
  FA1A U7110 ( .CI(n7743), .A(n7751), .B(n7739), .S(n7826), .CO(n7827) );
  FA1A U7111 ( .CI(n7814), .A(n7753), .B(n7741), .S(n7828), .CO(n7829) );
  FA1A U7112 ( .CI(n7767), .A(n7826), .B(n7763), .S(n7830), .CO(n7831) );
  FA1A U7113 ( .CI(n7822), .A(n7824), .B(n7761), .S(n7832), .CO(n7833) );
  FA1A U7114 ( .CI(n7818), .A(n7816), .B(n7755), .S(n7834), .CO(n7835) );
  FA1A U7115 ( .CI(n7820), .A(n7765), .B(n7759), .S(n7836), .CO(n7837) );
  FA1A U7116 ( .CI(n7769), .A(n7828), .B(n7757), .S(n7838), .CO(n7839) );
  FA1A U7117 ( .CI(n7834), .A(n7836), .B(n7775), .S(n7840), .CO(n7841) );
  FA1A U7118 ( .CI(n7832), .A(n7830), .B(n7771), .S(n7842), .CO(n7843) );
  FA1A U7119 ( .CI(n7838), .A(n7777), .B(n7773), .S(n7844), .CO(n7845) );
  FA1A U7120 ( .CI(n7844), .A(n7783), .B(n7779), .S(n7846), .CO(n7847) );
  FA1A U7121 ( .CI(n7842), .A(n7840), .B(n7781), .S(n7848), .CO(n7849) );
  FA1A U7122 ( .CI(n7846), .A(n7848), .B(n7785), .S(n7850), .CO(n7851) );
  FA1A U7123 ( .CI(n7850), .A(n7789), .B(n7787), .S(n7852), .CO(n7853) );
  IVP U7124 ( .A(n5775), .Z(n7854) );
  FA1A U7125 ( .CI(n3791), .A(n3727), .B(n7854), .S(n7855), .CO(n7856) );
  FA1A U7126 ( .CI(n5711), .A(n3855), .B(n4879), .S(n7857), .CO(n7858) );
  FA1A U7127 ( .CI(n3983), .A(n3919), .B(n4943), .S(n7859), .CO(n7860) );
  FA1A U7128 ( .CI(n4047), .A(n5647), .B(n5007), .S(n7861), .CO(n7862) );
  FA1A U7129 ( .CI(n5519), .A(n5583), .B(n5071), .S(n7863), .CO(n7864) );
  FA1A U7130 ( .CI(n4175), .A(n4111), .B(n4751), .S(n7865), .CO(n7866) );
  FA1A U7131 ( .CI(n4303), .A(n4239), .B(n5455), .S(n7867), .CO(n7868) );
  FA1A U7132 ( .CI(n5327), .A(n5391), .B(n4367), .S(n7869), .CO(n7870) );
  FA1A U7133 ( .CI(n5199), .A(n5263), .B(n4431), .S(n7871), .CO(n7872) );
  FA1A U7134 ( .CI(n4815), .A(n5135), .B(n4495), .S(n7873), .CO(n7874) );
  FA1A U7135 ( .CI(n4623), .A(n4687), .B(n4559), .S(n7875), .CO(n7876) );
  FA1A U7136 ( .CI(n7875), .A(n7793), .B(n7855), .S(n7877), .CO(n7878) );
  FA1A U7137 ( .CI(n7871), .A(n7873), .B(n7795), .S(n7879), .CO(n7880) );
  FA1A U7138 ( .CI(n7865), .A(n7869), .B(n7809), .S(n7881), .CO(n7882) );
  FA1A U7139 ( .CI(n7859), .A(n7857), .B(n7797), .S(n7883), .CO(n7884) );
  FA1A U7140 ( .CI(n7863), .A(n7867), .B(n7799), .S(n7885), .CO(n7886) );
  FA1A U7141 ( .CI(n7861), .A(n7813), .B(n7801), .S(n7887), .CO(n7888) );
  FA1A U7142 ( .CI(n7807), .A(n7811), .B(n7803), .S(n7889), .CO(n7890) );
  FA1A U7143 ( .CI(n7815), .A(n7877), .B(n7805), .S(n7891), .CO(n7892) );
  FA1A U7144 ( .CI(n7881), .A(n7889), .B(n7825), .S(n7893), .CO(n7894) );
  FA1A U7145 ( .CI(n7885), .A(n7887), .B(n7817), .S(n7895), .CO(n7896) );
  FA1A U7146 ( .CI(n7879), .A(n7883), .B(n7819), .S(n7897), .CO(n7898) );
  FA1A U7147 ( .CI(n7823), .A(n7827), .B(n7821), .S(n7899), .CO(n7900) );
  FA1A U7148 ( .CI(n7899), .A(n7891), .B(n7829), .S(n7901), .CO(n7902) );
  FA1A U7149 ( .CI(n7895), .A(n7897), .B(n7831), .S(n7903), .CO(n7904) );
  FA1A U7150 ( .CI(n7893), .A(n7837), .B(n7833), .S(n7905), .CO(n7906) );
  FA1A U7151 ( .CI(n7901), .A(n7839), .B(n7835), .S(n7907), .CO(n7908) );
  FA1A U7152 ( .CI(n7845), .A(n7903), .B(n7841), .S(n7909), .CO(n7910) );
  FA1A U7153 ( .CI(n7907), .A(n7905), .B(n7843), .S(n7911), .CO(n7912) );
  FA1A U7154 ( .CI(n7911), .A(n7909), .B(n7849), .S(n7913), .CO(n7914) );
  FA1A U7155 ( .CI(n7913), .A(n7851), .B(n7847), .S(n7915), .CO(n7916) );
  FA1A U7157 ( .CI(n3792), .A(n7854), .B(n5776), .S(n7918), .CO(n7919) );
  FA1A U7158 ( .CI(n5712), .A(n3856), .B(n4880), .S(n7920), .CO(n7921) );
  FA1A U7159 ( .CI(n3984), .A(n3920), .B(n4944), .S(n7922), .CO(n7923) );
  FA1A U7160 ( .CI(n4048), .A(n5648), .B(n5008), .S(n7924), .CO(n7925) );
  FA1A U7161 ( .CI(n5520), .A(n5584), .B(n5072), .S(n7926), .CO(n7927) );
  FA1A U7162 ( .CI(n4176), .A(n4112), .B(n4752), .S(n7928), .CO(n7929) );
  FA1A U7163 ( .CI(n4304), .A(n4240), .B(n5456), .S(n7930), .CO(n7931) );
  FA1A U7164 ( .CI(n5328), .A(n5392), .B(n4368), .S(n7932), .CO(n7933) );
  FA1A U7165 ( .CI(n5200), .A(n5264), .B(n4432), .S(n7934), .CO(n7935) );
  FA1A U7166 ( .CI(n4816), .A(n5136), .B(n4496), .S(n7936), .CO(n7937) );
  FA1A U7167 ( .CI(n4624), .A(n4688), .B(n4560), .S(n7938), .CO(n7939) );
  FA1A U7168 ( .CI(n7876), .A(n7856), .B(n7918), .S(n7940), .CO(n7941) );
  FA1A U7169 ( .CI(n7936), .A(n7938), .B(n7872), .S(n7942), .CO(n7943) );
  FA1A U7170 ( .CI(n7932), .A(n7934), .B(n7870), .S(n7944), .CO(n7945) );
  FA1A U7171 ( .CI(n7920), .A(n7930), .B(n7868), .S(n7946), .CO(n7947) );
  FA1A U7172 ( .CI(n7928), .A(n7922), .B(n7858), .S(n7948), .CO(n7949) );
  FA1A U7173 ( .CI(n7926), .A(n7924), .B(n7860), .S(n7950), .CO(n7951) );
  FA1A U7174 ( .CI(n7866), .A(n7874), .B(n7862), .S(n7952), .CO(n7953) );
  FA1A U7175 ( .CI(n7878), .A(n7940), .B(n7864), .S(n7954), .CO(n7955) );
  FA1A U7176 ( .CI(n7942), .A(n7952), .B(n7888), .S(n7956), .CO(n7957) );
  FA1A U7177 ( .CI(n7948), .A(n7950), .B(n7880), .S(n7958), .CO(n7959) );
  FA1A U7178 ( .CI(n7946), .A(n7944), .B(n7882), .S(n7960), .CO(n7961) );
  FA1A U7179 ( .CI(n7886), .A(n7890), .B(n7884), .S(n7962), .CO(n7963) );
  FA1A U7180 ( .CI(n7962), .A(n7892), .B(n7954), .S(n7964), .CO(n7965) );
  FA1A U7181 ( .CI(n7958), .A(n7960), .B(n7894), .S(n7966), .CO(n7967) );
  FA1A U7182 ( .CI(n7956), .A(n7900), .B(n7896), .S(n7968), .CO(n7969) );
  FA1A U7183 ( .CI(n7964), .A(n7902), .B(n7898), .S(n7970), .CO(n7971) );
  FA1A U7184 ( .CI(n7968), .A(n7966), .B(n7904), .S(n7972), .CO(n7973) );
  FA1A U7185 ( .CI(n7970), .A(n7908), .B(n7906), .S(n7974), .CO(n7975) );
  FA1A U7186 ( .CI(n7974), .A(n7972), .B(n7910), .S(n7976), .CO(n7977) );
  FA1A U7187 ( .CI(n7976), .A(n7914), .B(n7912), .S(n7978), .CO(n7979) );
  FA1A U7188 ( .CI(n3793), .A(n5777), .B(n5775), .S(n7980), .CO(n7981) );
  FA1A U7189 ( .CI(n7980), .A(n3857), .B(n4881), .S(n7982), .CO(n7983) );
  FA1A U7190 ( .CI(n5649), .A(n5713), .B(n3921), .S(n7984), .CO(n7985) );
  FA1A U7191 ( .CI(n4049), .A(n3985), .B(n4817), .S(n7986), .CO(n7987) );
  FA1A U7192 ( .CI(n5585), .A(n4113), .B(n5009), .S(n7988), .CO(n7989) );
  FA1A U7193 ( .CI(n5521), .A(n4177), .B(n4945), .S(n7990), .CO(n7991) );
  FA1A U7194 ( .CI(n4305), .A(n5457), .B(n4241), .S(n7992), .CO(n7993) );
  FA1A U7195 ( .CI(n4369), .A(n5393), .B(n4753), .S(n7994), .CO(n7995) );
  FA1A U7196 ( .CI(n5265), .A(n5329), .B(n4433), .S(n7996), .CO(n7997) );
  FA1A U7197 ( .CI(n5137), .A(n5201), .B(n4497), .S(n7998), .CO(n7999) );
  FA1A U7198 ( .CI(n4689), .A(n5073), .B(n4561), .S(n8000), .CO(n8001) );
  FA1A U7199 ( .CI(n7921), .A(n7919), .B(n4625), .S(n8002), .CO(n8003) );
  FA1A U7200 ( .CI(n7998), .A(n8000), .B(n7937), .S(n8004), .CO(n8005) );
  FA1A U7201 ( .CI(n7994), .A(n7996), .B(n7935), .S(n8006), .CO(n8007) );
  FA1A U7202 ( .CI(n7982), .A(n7992), .B(n7933), .S(n8008), .CO(n8009) );
  FA1A U7203 ( .CI(n7990), .A(n7984), .B(n7923), .S(n8010), .CO(n8011) );
  FA1A U7204 ( .CI(n7988), .A(n7986), .B(n7925), .S(n8012), .CO(n8013) );
  FA1A U7205 ( .CI(n7931), .A(n7939), .B(n7927), .S(n8014), .CO(n8015) );
  FA1A U7206 ( .CI(n7941), .A(n8002), .B(n7929), .S(n8016), .CO(n8017) );
  FA1A U7207 ( .CI(n8016), .A(n8014), .B(n7951), .S(n8018), .CO(n8019) );
  FA1A U7208 ( .CI(n8010), .A(n8012), .B(n7943), .S(n8020), .CO(n8021) );
  FA1A U7209 ( .CI(n8006), .A(n8008), .B(n7949), .S(n8022), .CO(n8023) );
  FA1A U7210 ( .CI(n8004), .A(n7953), .B(n7945), .S(n8024), .CO(n8025) );
  FA1A U7211 ( .CI(n7957), .A(n7955), .B(n7947), .S(n8026), .CO(n8027) );
  FA1A U7212 ( .CI(n8022), .A(n8024), .B(n7963), .S(n8028), .CO(n8029) );
  FA1A U7213 ( .CI(n8020), .A(n8018), .B(n7959), .S(n8030), .CO(n8031) );
  FA1A U7214 ( .CI(n7965), .A(n8026), .B(n7961), .S(n8032), .CO(n8033) );
  FA1A U7215 ( .CI(n8030), .A(n8028), .B(n7967), .S(n8034), .CO(n8035) );
  FA1A U7216 ( .CI(n7971), .A(n8032), .B(n7969), .S(n8036), .CO(n8037) );
  FA1A U7217 ( .CI(n7975), .A(n8034), .B(n7973), .S(n8038), .CO(n8039) );
  FA1A U7218 ( .CI(n8038), .A(n7977), .B(n8036), .S(n8040), .CO(n8041) );
  IVP U7219 ( .A(n5778), .Z(n8042) );
  FA1A U7220 ( .CI(n4882), .A(n3858), .B(n8042), .S(n8043), .CO(n8044) );
  FA1A U7221 ( .CI(n7981), .A(n5714), .B(n4946), .S(n8045), .CO(n8046) );
  FA1A U7222 ( .CI(n3922), .A(n5650), .B(n4818), .S(n8047), .CO(n8048) );
  FA1A U7223 ( .CI(n3986), .A(n5586), .B(n4754), .S(n8049), .CO(n8050) );
  FA1A U7224 ( .CI(n4114), .A(n4050), .B(n5010), .S(n8051), .CO(n8052) );
  FA1A U7225 ( .CI(n5522), .A(n4178), .B(n5138), .S(n8053), .CO(n8054) );
  FA1A U7226 ( .CI(n5458), .A(n4242), .B(n4626), .S(n8055), .CO(n8056) );
  FA1A U7227 ( .CI(n5330), .A(n5394), .B(n4306), .S(n8057), .CO(n8058) );
  FA1A U7228 ( .CI(n5202), .A(n5266), .B(n4370), .S(n8059), .CO(n8060) );
  FA1A U7229 ( .CI(n4690), .A(n5074), .B(n4434), .S(n8061), .CO(n8062) );
  FA1A U7230 ( .CI(n8043), .A(n4562), .B(n4498), .S(n8063), .CO(n8064) );
  FA1A U7231 ( .CI(n8063), .A(n8061), .B(n7983), .S(n8065), .CO(n8066) );
  FA1A U7232 ( .CI(n8057), .A(n8059), .B(n7997), .S(n8067), .CO(n8068) );
  FA1A U7233 ( .CI(n8053), .A(n8055), .B(n7985), .S(n8069), .CO(n8070) );
  FA1A U7234 ( .CI(n8049), .A(n8045), .B(n7987), .S(n8071), .CO(n8072) );
  FA1A U7235 ( .CI(n8051), .A(n8047), .B(n7989), .S(n8073), .CO(n8074) );
  FA1A U7236 ( .CI(n7999), .A(n8001), .B(n7991), .S(n8075), .CO(n8076) );
  FA1A U7237 ( .CI(n8003), .A(n7995), .B(n7993), .S(n8077), .CO(n8078) );
  FA1A U7238 ( .CI(n8077), .A(n8075), .B(n8013), .S(n8079), .CO(n8080) );
  FA1A U7239 ( .CI(n8071), .A(n8073), .B(n8005), .S(n8081), .CO(n8082) );
  FA1A U7240 ( .CI(n8067), .A(n8069), .B(n8011), .S(n8083), .CO(n8084) );
  FA1A U7241 ( .CI(n8065), .A(n8015), .B(n8007), .S(n8085), .CO(n8086) );
  FA1A U7242 ( .CI(n8019), .A(n8017), .B(n8009), .S(n8087), .CO(n8088) );
  FA1A U7243 ( .CI(n8083), .A(n8085), .B(n8025), .S(n8089), .CO(n8090) );
  FA1A U7244 ( .CI(n8081), .A(n8079), .B(n8021), .S(n8091), .CO(n8092) );
  FA1A U7245 ( .CI(n8027), .A(n8087), .B(n8023), .S(n8093), .CO(n8094) );
  FA1A U7246 ( .CI(n8093), .A(n8089), .B(n8029), .S(n8095), .CO(n8096) );
  FA1A U7247 ( .CI(n8033), .A(n8091), .B(n8031), .S(n8097), .CO(n8098) );
  FA1A U7248 ( .CI(n8097), .A(n8095), .B(n8035), .S(n8099), .CO(n8100) );
  FA1A U7249 ( .CI(n8099), .A(n8039), .B(n8037), .S(n8101), .CO(n8102) );
  FA1A U7250 ( .CI(n3859), .A(n5779), .B(n5778), .S(n8103), .CO(n8104) );
  FA1A U7251 ( .CI(n8103), .A(n5715), .B(n4883), .S(n8105), .CO(n8106) );
  FA1A U7252 ( .CI(n5587), .A(n5651), .B(n3923), .S(n8107), .CO(n8108) );
  FA1A U7253 ( .CI(n4051), .A(n3987), .B(n4819), .S(n8109), .CO(n8110) );
  FA1A U7254 ( .CI(n5459), .A(n5523), .B(n4947), .S(n8111), .CO(n8112) );
  FA1A U7255 ( .CI(n5331), .A(n5395), .B(n4115), .S(n8113), .CO(n8114) );
  FA1A U7256 ( .CI(n4243), .A(n4179), .B(n5203), .S(n8115), .CO(n8116) );
  FA1A U7257 ( .CI(n5139), .A(n5267), .B(n4627), .S(n8117), .CO(n8118) );
  FA1A U7258 ( .CI(n5011), .A(n5075), .B(n4307), .S(n8119), .CO(n8120) );
  FA1A U7259 ( .CI(n4691), .A(n4755), .B(n4371), .S(n8121), .CO(n8122) );
  FA1A U7260 ( .CI(n4499), .A(n4563), .B(n4435), .S(n8123), .CO(n8124) );
  FA1A U7261 ( .CI(n8121), .A(n8123), .B(n8044), .S(n8125), .CO(n8126) );
  FA1A U7262 ( .CI(n8064), .A(n8119), .B(n8058), .S(n8127), .CO(n8128) );
  FA1A U7263 ( .CI(n8115), .A(n8117), .B(n8056), .S(n8129), .CO(n8130) );
  FA1A U7264 ( .CI(n8107), .A(n8105), .B(n8046), .S(n8131), .CO(n8132) );
  FA1A U7265 ( .CI(n8113), .A(n8109), .B(n8048), .S(n8133), .CO(n8134) );
  FA1A U7266 ( .CI(n8111), .A(n8062), .B(n8050), .S(n8135), .CO(n8136) );
  FA1A U7267 ( .CI(n8054), .A(n8060), .B(n8052), .S(n8137), .CO(n8138) );
  FA1A U7268 ( .CI(n8078), .A(n8137), .B(n8125), .S(n8139), .CO(n8140) );
  FA1A U7269 ( .CI(n8133), .A(n8135), .B(n8066), .S(n8141), .CO(n8142) );
  FA1A U7270 ( .CI(n8127), .A(n8131), .B(n8072), .S(n8143), .CO(n8144) );
  FA1A U7271 ( .CI(n8129), .A(n8076), .B(n8068), .S(n8145), .CO(n8146) );
  FA1A U7272 ( .CI(n8139), .A(n8074), .B(n8070), .S(n8147), .CO(n8148) );
  FA1A U7273 ( .CI(n8143), .A(n8145), .B(n8080), .S(n8149), .CO(n8150) );
  FA1A U7274 ( .CI(n8141), .A(n8086), .B(n8082), .S(n8151), .CO(n8152) );
  FA1A U7275 ( .CI(n8088), .A(n8147), .B(n8084), .S(n8153), .CO(n8154) );
  FA1A U7276 ( .CI(n8153), .A(n8149), .B(n8090), .S(n8155), .CO(n8156) );
  FA1A U7277 ( .CI(n8094), .A(n8151), .B(n8092), .S(n8157), .CO(n8158) );
  FA1A U7278 ( .CI(n8098), .A(n8157), .B(n8096), .S(n8159), .CO(n8160) );
  FA1A U7279 ( .CI(n8159), .A(n8100), .B(n8155), .S(n8161), .CO(n8162) );
  IVP U7280 ( .A(n5780), .Z(n8163) );
  FA1A U7281 ( .CI(n4948), .A(n3924), .B(n8163), .S(n8164), .CO(n8165) );
  FA1A U7282 ( .CI(n8104), .A(n5716), .B(n5012), .S(n8166), .CO(n8167) );
  FA1A U7283 ( .CI(n4052), .A(n3988), .B(n4820), .S(n8168), .CO(n8169) );
  FA1A U7284 ( .CI(n4116), .A(n5652), .B(n5076), .S(n8170), .CO(n8171) );
  FA1A U7285 ( .CI(n5524), .A(n5588), .B(n4884), .S(n8172), .CO(n8173) );
  FA1A U7286 ( .CI(n4244), .A(n4180), .B(n4756), .S(n8174), .CO(n8175) );
  FA1A U7287 ( .CI(n5396), .A(n5460), .B(n4628), .S(n8176), .CO(n8177) );
  FA1A U7288 ( .CI(n5268), .A(n5332), .B(n4308), .S(n8178), .CO(n8179) );
  FA1A U7289 ( .CI(n5140), .A(n5204), .B(n4372), .S(n8180), .CO(n8181) );
  FA1A U7290 ( .CI(n4564), .A(n4692), .B(n4436), .S(n8182), .CO(n8183) );
  FA1A U7291 ( .CI(n8106), .A(n8164), .B(n4500), .S(n8184), .CO(n8185) );
  FA1A U7292 ( .CI(n8180), .A(n8182), .B(n8122), .S(n8186), .CO(n8187) );
  FA1A U7293 ( .CI(n8176), .A(n8178), .B(n8118), .S(n8188), .CO(n8189) );
  FA1A U7294 ( .CI(n8168), .A(n8166), .B(n8108), .S(n8190), .CO(n8191) );
  FA1A U7295 ( .CI(n8172), .A(n8170), .B(n8110), .S(n8192), .CO(n8193) );
  FA1A U7296 ( .CI(n8174), .A(n8124), .B(n8112), .S(n8194), .CO(n8195) );
  FA1A U7297 ( .CI(n8116), .A(n8120), .B(n8114), .S(n8196), .CO(n8197) );
  FA1A U7298 ( .CI(n8196), .A(n8126), .B(n8184), .S(n8198), .CO(n8199) );
  FA1A U7299 ( .CI(n8192), .A(n8194), .B(n8128), .S(n8200), .CO(n8201) );
  FA1A U7300 ( .CI(n8186), .A(n8190), .B(n8134), .S(n8202), .CO(n8203) );
  FA1A U7301 ( .CI(n8188), .A(n8138), .B(n8130), .S(n8204), .CO(n8205) );
  FA1A U7302 ( .CI(n8198), .A(n8136), .B(n8132), .S(n8206), .CO(n8207) );
  FA1A U7303 ( .CI(n8206), .A(n8204), .B(n8140), .S(n8208), .CO(n8209) );
  FA1A U7304 ( .CI(n8200), .A(n8202), .B(n8142), .S(n8210), .CO(n8211) );
  FA1A U7305 ( .CI(n8148), .A(n8146), .B(n8144), .S(n8212), .CO(n8213) );
  FA1A U7306 ( .CI(n8212), .A(n8210), .B(n8208), .S(n8214), .CO(n8215) );
  FA1A U7307 ( .CI(n8154), .A(n8152), .B(n8150), .S(n8216), .CO(n8217) );
  FA1A U7308 ( .CI(n8158), .A(n8216), .B(n8214), .S(n8218), .CO(n8219) );
  FA1A U7309 ( .CI(n8160), .A(n8218), .B(n8156), .S(n8220), .CO(n8221) );
  FA1A U7310 ( .CI(n3925), .A(n5781), .B(n5780), .S(n8222), .CO(n8223) );
  FA1A U7311 ( .CI(n8222), .A(n3989), .B(n4949), .S(n8224), .CO(n8225) );
  FA1A U7312 ( .CI(n5653), .A(n5717), .B(n4053), .S(n8226), .CO(n8227) );
  FA1A U7313 ( .CI(n4181), .A(n4117), .B(n4885), .S(n8228), .CO(n8229) );
  FA1A U7314 ( .CI(n4309), .A(n4245), .B(n5013), .S(n8230), .CO(n8231) );
  FA1A U7315 ( .CI(n5525), .A(n5589), .B(n4373), .S(n8232), .CO(n8233) );
  FA1A U7316 ( .CI(n5397), .A(n4437), .B(n5461), .S(n8234), .CO(n8235) );
  FA1A U7317 ( .CI(n5269), .A(n5333), .B(n4501), .S(n8236), .CO(n8237) );
  FA1A U7318 ( .CI(n5141), .A(n5205), .B(n4565), .S(n8238), .CO(n8239) );
  FA1A U7319 ( .CI(n4821), .A(n5077), .B(n4629), .S(n8240), .CO(n8241) );
  FA1A U7320 ( .CI(n8165), .A(n4757), .B(n4693), .S(n8242), .CO(n8243) );
  FA1A U7321 ( .CI(n8238), .A(n8240), .B(n8181), .S(n8244), .CO(n8245) );
  FA1A U7322 ( .CI(n8234), .A(n8236), .B(n8177), .S(n8246), .CO(n8247) );
  FA1A U7323 ( .CI(n8226), .A(n8224), .B(n8167), .S(n8248), .CO(n8249) );
  FA1A U7324 ( .CI(n8230), .A(n8228), .B(n8169), .S(n8250), .CO(n8251) );
  FA1A U7325 ( .CI(n8232), .A(n8183), .B(n8171), .S(n8252), .CO(n8253) );
  FA1A U7326 ( .CI(n8175), .A(n8179), .B(n8173), .S(n8254), .CO(n8255) );
  FA1A U7327 ( .CI(n8187), .A(n8185), .B(n8242), .S(n8256), .CO(n8257) );
  FA1A U7328 ( .CI(n8252), .A(n8254), .B(n8197), .S(n8258), .CO(n8259) );
  FA1A U7329 ( .CI(n8248), .A(n8250), .B(n8193), .S(n8260), .CO(n8261) );
  FA1A U7330 ( .CI(n8244), .A(n8246), .B(n8189), .S(n8262), .CO(n8263) );
  FA1A U7331 ( .CI(n8256), .A(n8195), .B(n8191), .S(n8264), .CO(n8265) );
  FA1A U7332 ( .CI(n8264), .A(n8262), .B(n8199), .S(n8266), .CO(n8267) );
  FA1A U7333 ( .CI(n8207), .A(n8260), .B(n8201), .S(n8268), .CO(n8269) );
  FA1A U7334 ( .CI(n8258), .A(n8205), .B(n8203), .S(n8270), .CO(n8271) );
  FA1A U7335 ( .CI(n8213), .A(n8270), .B(n8266), .S(n8272), .CO(n8273) );
  FA1A U7336 ( .CI(n8268), .A(n8211), .B(n8209), .S(n8274), .CO(n8275) );
  FA1A U7337 ( .CI(n8217), .A(n8274), .B(n8272), .S(n8276), .CO(n8277) );
  FA1A U7338 ( .CI(n8219), .A(n8276), .B(n8215), .S(n8278), .CO(n8279) );
  IVP U7339 ( .A(n5782), .Z(n8280) );
  FA1A U7340 ( .CI(n4054), .A(n3990), .B(n8280), .S(n8281), .CO(n8282) );
  FA1A U7341 ( .CI(n8223), .A(n5718), .B(n5014), .S(n8283), .CO(n8284) );
  FA1A U7342 ( .CI(n4182), .A(n4118), .B(n4950), .S(n8285), .CO(n8286) );
  FA1A U7343 ( .CI(n4310), .A(n4246), .B(n5078), .S(n8287), .CO(n8288) );
  FA1A U7344 ( .CI(n4374), .A(n5654), .B(n5206), .S(n8289), .CO(n8290) );
  FA1A U7345 ( .CI(n4438), .A(n5590), .B(n5526), .S(n8291), .CO(n8292) );
  FA1A U7346 ( .CI(n5398), .A(n5462), .B(n4502), .S(n8293), .CO(n8294) );
  FA1A U7347 ( .CI(n5270), .A(n5334), .B(n4566), .S(n8295), .CO(n8296) );
  FA1A U7348 ( .CI(n4886), .A(n5142), .B(n4630), .S(n8297), .CO(n8298) );
  FA1A U7349 ( .CI(n4822), .A(n4758), .B(n4694), .S(n8299), .CO(n8300) );
  FA1A U7350 ( .CI(n8299), .A(n8241), .B(n8281), .S(n8301), .CO(n8302) );
  FA1A U7351 ( .CI(n8283), .A(n8297), .B(n8237), .S(n8303), .CO(n8304) );
  FA1A U7352 ( .CI(n8285), .A(n8295), .B(n8225), .S(n8305), .CO(n8306) );
  FA1A U7353 ( .CI(n8291), .A(n8293), .B(n8227), .S(n8307), .CO(n8308) );
  FA1A U7354 ( .CI(n8289), .A(n8287), .B(n8229), .S(n8309), .CO(n8310) );
  FA1A U7355 ( .CI(n8235), .A(n8239), .B(n8231), .S(n8311), .CO(n8312) );
  FA1A U7356 ( .CI(n8301), .A(n8243), .B(n8233), .S(n8313), .CO(n8314) );
  FA1A U7357 ( .CI(n8313), .A(n8311), .B(n8245), .S(n8315), .CO(n8316) );
  FA1A U7358 ( .CI(n8307), .A(n8309), .B(n8253), .S(n8317), .CO(n8318) );
  FA1A U7359 ( .CI(n8305), .A(n8303), .B(n8247), .S(n8319), .CO(n8320) );
  FA1A U7360 ( .CI(n8251), .A(n8255), .B(n8249), .S(n8321), .CO(n8322) );
  FA1A U7361 ( .CI(n8321), .A(n8259), .B(n8257), .S(n8323), .CO(n8324) );
  FA1A U7362 ( .CI(n8265), .A(n8315), .B(n8261), .S(n8325), .CO(n8326) );
  FA1A U7363 ( .CI(n8319), .A(n8317), .B(n8263), .S(n8327), .CO(n8328) );
  FA1A U7364 ( .CI(n8327), .A(n8271), .B(n8323), .S(n8329), .CO(n8330) );
  FA1A U7365 ( .CI(n8325), .A(n8269), .B(n8267), .S(n8331), .CO(n8332) );
  FA1A U7366 ( .CI(n8331), .A(n8275), .B(n8329), .S(n8333), .CO(n8334) );
  FA1A U7367 ( .CI(n8277), .A(n8333), .B(n8273), .S(n8335), .CO(n8336) );
  FA1A U7368 ( .CI(n3991), .A(n5783), .B(n5782), .S(n8337), .CO(n8338) );
  FA1A U7369 ( .CI(n8337), .A(n4055), .B(n4951), .S(n8339), .CO(n8340) );
  FA1A U7370 ( .CI(n5655), .A(n5719), .B(n4119), .S(n8341), .CO(n8342) );
  FA1A U7371 ( .CI(n4247), .A(n4183), .B(n5015), .S(n8343), .CO(n8344) );
  FA1A U7372 ( .CI(n5527), .A(n5591), .B(n5079), .S(n8345), .CO(n8346) );
  FA1A U7373 ( .CI(n5399), .A(n5463), .B(n4311), .S(n8347), .CO(n8348) );
  FA1A U7374 ( .CI(n4375), .A(n5271), .B(n5335), .S(n8349), .CO(n8350) );
  FA1A U7375 ( .CI(n5143), .A(n5207), .B(n4439), .S(n8351), .CO(n8352) );
  FA1A U7376 ( .CI(n4823), .A(n4887), .B(n4503), .S(n8353), .CO(n8354) );
  FA1A U7377 ( .CI(n4695), .A(n4759), .B(n4567), .S(n8355), .CO(n8356) );
  FA1A U7378 ( .CI(n8284), .A(n8282), .B(n4631), .S(n8357), .CO(n8358) );
  FA1A U7379 ( .CI(n8353), .A(n8355), .B(n8298), .S(n8359), .CO(n8360) );
  FA1A U7380 ( .CI(n8349), .A(n8351), .B(n8296), .S(n8361), .CO(n8362) );
  FA1A U7381 ( .CI(n8345), .A(n8347), .B(n8286), .S(n8363), .CO(n8364) );
  FA1A U7382 ( .CI(n8343), .A(n8339), .B(n8288), .S(n8365), .CO(n8366) );
  FA1A U7383 ( .CI(n8341), .A(n8300), .B(n8290), .S(n8367), .CO(n8368) );
  FA1A U7384 ( .CI(n8357), .A(n8294), .B(n8292), .S(n8369), .CO(n8370) );
  FA1A U7385 ( .CI(n8369), .A(n8367), .B(n8302), .S(n8371), .CO(n8372) );
  FA1A U7386 ( .CI(n8314), .A(n8365), .B(n8310), .S(n8373), .CO(n8374) );
  FA1A U7387 ( .CI(n8359), .A(n8363), .B(n8308), .S(n8375), .CO(n8376) );
  FA1A U7388 ( .CI(n8361), .A(n8312), .B(n8304), .S(n8377), .CO(n8378) );
  FA1A U7389 ( .CI(n8316), .A(n8371), .B(n8306), .S(n8379), .CO(n8380) );
  FA1A U7390 ( .CI(n8375), .A(n8377), .B(n8318), .S(n8381), .CO(n8382) );
  FA1A U7391 ( .CI(n8373), .A(n8322), .B(n8320), .S(n8383), .CO(n8384) );
  FA1A U7392 ( .CI(n8383), .A(n8324), .B(n8379), .S(n8385), .CO(n8386) );
  FA1A U7393 ( .CI(n8381), .A(n8328), .B(n8326), .S(n8387), .CO(n8388) );
  FA1A U7394 ( .CI(n8387), .A(n8332), .B(n8385), .S(n8389), .CO(n8390) );
  FA1A U7395 ( .CI(n8334), .A(n8389), .B(n8330), .S(n8391), .CO(n8392) );
  IVP U7396 ( .A(n5784), .Z(n8393) );
  FA1A U7397 ( .CI(n4952), .A(n4056), .B(n8393), .S(n8394), .CO(n8395) );
  FA1A U7398 ( .CI(n8338), .A(n5720), .B(n5016), .S(n8396), .CO(n8397) );
  FA1A U7399 ( .CI(n4184), .A(n4120), .B(n4888), .S(n8398), .CO(n8399) );
  FA1A U7400 ( .CI(n5656), .A(n4248), .B(n5080), .S(n8400), .CO(n8401) );
  FA1A U7401 ( .CI(n4312), .A(n5592), .B(n5144), .S(n8402), .CO(n8403) );
  FA1A U7402 ( .CI(n5528), .A(n4376), .B(n5464), .S(n8404), .CO(n8405) );
  FA1A U7403 ( .CI(n5336), .A(n5400), .B(n4440), .S(n8406), .CO(n8407) );
  FA1A U7404 ( .CI(n5208), .A(n5272), .B(n4504), .S(n8408), .CO(n8409) );
  FA1A U7405 ( .CI(n4760), .A(n4824), .B(n4568), .S(n8410), .CO(n8411) );
  FA1A U7406 ( .CI(n8394), .A(n4632), .B(n4696), .S(n8412), .CO(n8413) );
  FA1A U7407 ( .CI(n8412), .A(n8410), .B(n8352), .S(n8414), .CO(n8415) );
  FA1A U7408 ( .CI(n8408), .A(n8406), .B(n8340), .S(n8416), .CO(n8417) );
  FA1A U7409 ( .CI(n8396), .A(n8404), .B(n8342), .S(n8418), .CO(n8419) );
  FA1A U7410 ( .CI(n8398), .A(n8400), .B(n8344), .S(n8420), .CO(n8421) );
  FA1A U7411 ( .CI(n8402), .A(n8356), .B(n8346), .S(n8422), .CO(n8423) );
  FA1A U7412 ( .CI(n8350), .A(n8354), .B(n8348), .S(n8424), .CO(n8425) );
  FA1A U7413 ( .CI(n8422), .A(n8424), .B(n8358), .S(n8426), .CO(n8427) );
  FA1A U7414 ( .CI(n8370), .A(n8420), .B(n8366), .S(n8428), .CO(n8429) );
  FA1A U7415 ( .CI(n8414), .A(n8418), .B(n8364), .S(n8430), .CO(n8431) );
  FA1A U7416 ( .CI(n8416), .A(n8368), .B(n8360), .S(n8432), .CO(n8433) );
  FA1A U7417 ( .CI(n8372), .A(n8426), .B(n8362), .S(n8434), .CO(n8435) );
  FA1A U7418 ( .CI(n8430), .A(n8432), .B(n8374), .S(n8436), .CO(n8437) );
  FA1A U7419 ( .CI(n8428), .A(n8378), .B(n8376), .S(n8438), .CO(n8439) );
  FA1A U7420 ( .CI(n8438), .A(n8380), .B(n8434), .S(n8440), .CO(n8441) );
  FA1A U7421 ( .CI(n8436), .A(n8384), .B(n8382), .S(n8442), .CO(n8443) );
  FA1A U7422 ( .CI(n8442), .A(n8386), .B(n8440), .S(n8444), .CO(n8445) );
  FA1A U7423 ( .CI(n8390), .A(n8444), .B(n8388), .S(n8446), .CO(n8447) );
  FA1A U7424 ( .CI(n4057), .A(n5785), .B(n5784), .S(n8448), .CO(n8449) );
  FA1A U7425 ( .CI(n8448), .A(n5721), .B(n5017), .S(n8450), .CO(n8451) );
  FA1A U7426 ( .CI(n4185), .A(n5657), .B(n4121), .S(n8452), .CO(n8453) );
  FA1A U7427 ( .CI(n4313), .A(n4249), .B(n4953), .S(n8454), .CO(n8455) );
  FA1A U7428 ( .CI(n5529), .A(n5593), .B(n5145), .S(n8456), .CO(n8457) );
  FA1A U7429 ( .CI(n5401), .A(n5465), .B(n4377), .S(n8458), .CO(n8459) );
  FA1A U7430 ( .CI(n5337), .A(n4441), .B(n4761), .S(n8460), .CO(n8461) );
  FA1A U7431 ( .CI(n5209), .A(n5273), .B(n4505), .S(n8462), .CO(n8463) );
  FA1A U7432 ( .CI(n4889), .A(n5081), .B(n4569), .S(n8464), .CO(n8465) );
  FA1A U7433 ( .CI(n4697), .A(n4825), .B(n4633), .S(n8466), .CO(n8467) );
  FA1A U7434 ( .CI(n8464), .A(n8466), .B(n8395), .S(n8468), .CO(n8469) );
  FA1A U7435 ( .CI(n8413), .A(n8450), .B(n8397), .S(n8470), .CO(n8471) );
  FA1A U7436 ( .CI(n8460), .A(n8462), .B(n8399), .S(n8472), .CO(n8473) );
  FA1A U7437 ( .CI(n8454), .A(n8458), .B(n8407), .S(n8474), .CO(n8475) );
  FA1A U7438 ( .CI(n8452), .A(n8456), .B(n8401), .S(n8476), .CO(n8477) );
  FA1A U7439 ( .CI(n8409), .A(n8411), .B(n8403), .S(n8478), .CO(n8479) );
  FA1A U7440 ( .CI(n8415), .A(n8468), .B(n8405), .S(n8480), .CO(n8481) );
  FA1A U7441 ( .CI(n8476), .A(n8478), .B(n8423), .S(n8482), .CO(n8483) );
  FA1A U7442 ( .CI(n8470), .A(n8474), .B(n8421), .S(n8484), .CO(n8485) );
  FA1A U7443 ( .CI(n8472), .A(n8425), .B(n8417), .S(n8486), .CO(n8487) );
  FA1A U7444 ( .CI(n8427), .A(n8480), .B(n8419), .S(n8488), .CO(n8489) );
  FA1A U7445 ( .CI(n8484), .A(n8486), .B(n8429), .S(n8490), .CO(n8491) );
  FA1A U7446 ( .CI(n8482), .A(n8433), .B(n8431), .S(n8492), .CO(n8493) );
  FA1A U7447 ( .CI(n8492), .A(n8435), .B(n8488), .S(n8494), .CO(n8495) );
  FA1A U7448 ( .CI(n8490), .A(n8439), .B(n8437), .S(n8496), .CO(n8497) );
  FA1A U7449 ( .CI(n8496), .A(n8441), .B(n8494), .S(n8498), .CO(n8499) );
  FA1A U7450 ( .CI(n8445), .A(n8498), .B(n8443), .S(n8500), .CO(n8501) );
  IVP U7451 ( .A(n5786), .Z(n8502) );
  FA1A U7452 ( .CI(n5018), .A(n4122), .B(n8502), .S(n8503), .CO(n8504) );
  FA1A U7453 ( .CI(n8449), .A(n4186), .B(n5082), .S(n8505), .CO(n8506) );
  FA1A U7454 ( .CI(n5722), .A(n4250), .B(n5146), .S(n8507), .CO(n8508) );
  FA1A U7455 ( .CI(n4378), .A(n4314), .B(n4954), .S(n8509), .CO(n8510) );
  FA1A U7456 ( .CI(n5594), .A(n5658), .B(n5274), .S(n8511), .CO(n8512) );
  FA1A U7457 ( .CI(n4506), .A(n4442), .B(n5530), .S(n8513), .CO(n8514) );
  FA1A U7458 ( .CI(n5402), .A(n5466), .B(n4570), .S(n8515), .CO(n8516) );
  FA1A U7459 ( .CI(n5210), .A(n5338), .B(n4634), .S(n8517), .CO(n8518) );
  FA1A U7460 ( .CI(n4826), .A(n4890), .B(n4698), .S(n8519), .CO(n8520) );
  FA1A U7461 ( .CI(n8451), .A(n8503), .B(n4762), .S(n8521), .CO(n8522) );
  FA1A U7462 ( .CI(n8505), .A(n8519), .B(n8465), .S(n8523), .CO(n8524) );
  FA1A U7463 ( .CI(n8515), .A(n8517), .B(n8453), .S(n8525), .CO(n8526) );
  FA1A U7464 ( .CI(n8509), .A(n8513), .B(n8461), .S(n8527), .CO(n8528) );
  FA1A U7465 ( .CI(n8507), .A(n8511), .B(n8455), .S(n8529), .CO(n8530) );
  FA1A U7466 ( .CI(n8463), .A(n8467), .B(n8457), .S(n8531), .CO(n8532) );
  FA1A U7467 ( .CI(n8469), .A(n8521), .B(n8459), .S(n8533), .CO(n8534) );
  FA1A U7468 ( .CI(n8529), .A(n8531), .B(n8477), .S(n8535), .CO(n8536) );
  FA1A U7469 ( .CI(n8523), .A(n8527), .B(n8475), .S(n8537), .CO(n8538) );
  FA1A U7470 ( .CI(n8525), .A(n8479), .B(n8471), .S(n8539), .CO(n8540) );
  FA1A U7471 ( .CI(n8481), .A(n8533), .B(n8473), .S(n8541), .CO(n8542) );
  FA1A U7472 ( .CI(n8537), .A(n8539), .B(n8483), .S(n8543), .CO(n8544) );
  FA1A U7473 ( .CI(n8535), .A(n8487), .B(n8485), .S(n8545), .CO(n8546) );
  FA1A U7474 ( .CI(n8545), .A(n8489), .B(n8541), .S(n8547), .CO(n8548) );
  FA1A U7475 ( .CI(n8543), .A(n8493), .B(n8491), .S(n8549), .CO(n8550) );
  FA1A U7476 ( .CI(n8549), .A(n8495), .B(n8547), .S(n8551), .CO(n8552) );
  FA1A U7477 ( .CI(n8499), .A(n8551), .B(n8497), .S(n8553), .CO(n8554) );
  FA1A U7478 ( .CI(n4123), .A(n5787), .B(n5786), .S(n8555), .CO(n8556) );
  FA1A U7479 ( .CI(n8555), .A(n5723), .B(n5019), .S(n8557), .CO(n8558) );
  FA1A U7480 ( .CI(n4251), .A(n5659), .B(n4187), .S(n8559), .CO(n8560) );
  FA1A U7481 ( .CI(n5595), .A(n4315), .B(n4955), .S(n8561), .CO(n8562) );
  FA1A U7482 ( .CI(n5467), .A(n5531), .B(n5083), .S(n8563), .CO(n8564) );
  FA1A U7483 ( .CI(n4443), .A(n5403), .B(n4379), .S(n8565), .CO(n8566) );
  FA1A U7484 ( .CI(n5275), .A(n5339), .B(n4827), .S(n8567), .CO(n8568) );
  FA1A U7485 ( .CI(n5147), .A(n5211), .B(n4507), .S(n8569), .CO(n8570) );
  FA1A U7486 ( .CI(n4763), .A(n4891), .B(n4571), .S(n8571), .CO(n8572) );
  FA1A U7487 ( .CI(n8504), .A(n4699), .B(n4635), .S(n8573), .CO(n8574) );
  FA1A U7488 ( .CI(n8557), .A(n8571), .B(n8518), .S(n8575), .CO(n8576) );
  FA1A U7489 ( .CI(n8567), .A(n8569), .B(n8506), .S(n8577), .CO(n8578) );
  FA1A U7490 ( .CI(n8561), .A(n8565), .B(n8514), .S(n8579), .CO(n8580) );
  FA1A U7491 ( .CI(n8559), .A(n8563), .B(n8508), .S(n8581), .CO(n8582) );
  FA1A U7492 ( .CI(n8516), .A(n8520), .B(n8510), .S(n8583), .CO(n8584) );
  FA1A U7493 ( .CI(n8522), .A(n8573), .B(n8512), .S(n8585), .CO(n8586) );
  FA1A U7494 ( .CI(n8585), .A(n8583), .B(n8530), .S(n8587), .CO(n8588) );
  FA1A U7495 ( .CI(n8575), .A(n8581), .B(n8528), .S(n8589), .CO(n8590) );
  FA1A U7496 ( .CI(n8579), .A(n8577), .B(n8524), .S(n8591), .CO(n8592) );
  FA1A U7497 ( .CI(n8534), .A(n8532), .B(n8526), .S(n8593), .CO(n8594) );
  FA1A U7498 ( .CI(n8593), .A(n8591), .B(n8536), .S(n8595), .CO(n8596) );
  FA1A U7499 ( .CI(n8589), .A(n8587), .B(n8538), .S(n8597), .CO(n8598) );
  FA1A U7500 ( .CI(n8544), .A(n8542), .B(n8540), .S(n8599), .CO(n8600) );
  FA1A U7501 ( .CI(n8597), .A(n8595), .B(n8546), .S(n8601), .CO(n8602) );
  FA1A U7502 ( .CI(n8601), .A(n8548), .B(n8599), .S(n8603), .CO(n8604) );
  FA1A U7503 ( .CI(n8552), .A(n8603), .B(n8550), .S(n8605), .CO(n8606) );
  IVP U7504 ( .A(n5788), .Z(n8607) );
  FA1A U7505 ( .CI(n4252), .A(n4188), .B(n8607), .S(n8608), .CO(n8609) );
  FA1A U7506 ( .CI(n8556), .A(n4316), .B(n5084), .S(n8610), .CO(n8611) );
  FA1A U7507 ( .CI(n4444), .A(n4380), .B(n5148), .S(n8612), .CO(n8613) );
  FA1A U7508 ( .CI(n5724), .A(n4508), .B(n5276), .S(n8614), .CO(n8615) );
  FA1A U7509 ( .CI(n5596), .A(n5660), .B(n5212), .S(n8616), .CO(n8617) );
  FA1A U7510 ( .CI(n5468), .A(n4572), .B(n5532), .S(n8618), .CO(n8619) );
  FA1A U7511 ( .CI(n5340), .A(n5404), .B(n4636), .S(n8620), .CO(n8621) );
  FA1A U7512 ( .CI(n4956), .A(n5020), .B(n4700), .S(n8622), .CO(n8623) );
  FA1A U7513 ( .CI(n4828), .A(n4892), .B(n4764), .S(n8624), .CO(n8625) );
  FA1A U7514 ( .CI(n8624), .A(n8572), .B(n8608), .S(n8626), .CO(n8627) );
  FA1A U7515 ( .CI(n8620), .A(n8622), .B(n8558), .S(n8628), .CO(n8629) );
  FA1A U7516 ( .CI(n8610), .A(n8618), .B(n8568), .S(n8630), .CO(n8631) );
  FA1A U7517 ( .CI(n8614), .A(n8612), .B(n8560), .S(n8632), .CO(n8633) );
  FA1A U7518 ( .CI(n8616), .A(n8570), .B(n8562), .S(n8634), .CO(n8635) );
  FA1A U7519 ( .CI(n8574), .A(n8566), .B(n8564), .S(n8636), .CO(n8637) );
  FA1A U7520 ( .CI(n8636), .A(n8634), .B(n8626), .S(n8638), .CO(n8639) );
  FA1A U7521 ( .CI(n8586), .A(n8630), .B(n8576), .S(n8640), .CO(n8641) );
  FA1A U7522 ( .CI(n8632), .A(n8628), .B(n8578), .S(n8642), .CO(n8643) );
  FA1A U7523 ( .CI(n8582), .A(n8584), .B(n8580), .S(n8644), .CO(n8645) );
  FA1A U7524 ( .CI(n8594), .A(n8644), .B(n8638), .S(n8646), .CO(n8647) );
  FA1A U7525 ( .CI(n8640), .A(n8642), .B(n8588), .S(n8648), .CO(n8649) );
  FA1A U7526 ( .CI(n8646), .A(n8592), .B(n8590), .S(n8650), .CO(n8651) );
  FA1A U7527 ( .CI(n8650), .A(n8648), .B(n8596), .S(n8652), .CO(n8653) );
  FA1A U7528 ( .CI(n8602), .A(n8600), .B(n8598), .S(n8654), .CO(n8655) );
  FA1A U7529 ( .CI(n8604), .A(n8654), .B(n8652), .S(n8656), .CO(n8657) );
  FA1A U7530 ( .CI(n4189), .A(n5789), .B(n5788), .S(n8658), .CO(n8659) );
  FA1A U7531 ( .CI(n8658), .A(n4253), .B(n5085), .S(n8660), .CO(n8661) );
  FA1A U7532 ( .CI(n5661), .A(n5725), .B(n4317), .S(n8662), .CO(n8663) );
  FA1A U7533 ( .CI(n4381), .A(n5597), .B(n5021), .S(n8664), .CO(n8665) );
  FA1A U7534 ( .CI(n5469), .A(n5533), .B(n5149), .S(n8666), .CO(n8667) );
  FA1A U7535 ( .CI(n4509), .A(n5405), .B(n4445), .S(n8668), .CO(n8669) );
  FA1A U7536 ( .CI(n5277), .A(n5341), .B(n4893), .S(n8670), .CO(n8671) );
  FA1A U7537 ( .CI(n4957), .A(n5213), .B(n4573), .S(n8672), .CO(n8673) );
  FA1A U7538 ( .CI(n4765), .A(n4829), .B(n4637), .S(n8674), .CO(n8675) );
  FA1A U7539 ( .CI(n8611), .A(n8609), .B(n4701), .S(n8676), .CO(n8677) );
  FA1A U7540 ( .CI(n8672), .A(n8674), .B(n8623), .S(n8678), .CO(n8679) );
  FA1A U7541 ( .CI(n8668), .A(n8670), .B(n8621), .S(n8680), .CO(n8681) );
  FA1A U7542 ( .CI(n8660), .A(n8666), .B(n8619), .S(n8682), .CO(n8683) );
  FA1A U7543 ( .CI(n8662), .A(n8664), .B(n8613), .S(n8684), .CO(n8685) );
  FA1A U7544 ( .CI(n8625), .A(n8617), .B(n8615), .S(n8686), .CO(n8687) );
  FA1A U7545 ( .CI(n8686), .A(n8627), .B(n8676), .S(n8688), .CO(n8689) );
  FA1A U7546 ( .CI(n8678), .A(n8684), .B(n8635), .S(n8690), .CO(n8691) );
  FA1A U7547 ( .CI(n8682), .A(n8680), .B(n8629), .S(n8692), .CO(n8693) );
  FA1A U7548 ( .CI(n8637), .A(n8633), .B(n8631), .S(n8694), .CO(n8695) );
  FA1A U7549 ( .CI(n8694), .A(n8639), .B(n8688), .S(n8696), .CO(n8697) );
  FA1A U7550 ( .CI(n8690), .A(n8692), .B(n8641), .S(n8698), .CO(n8699) );
  FA1A U7551 ( .CI(n8696), .A(n8645), .B(n8643), .S(n8700), .CO(n8701) );
  FA1A U7552 ( .CI(n8700), .A(n8698), .B(n8647), .S(n8702), .CO(n8703) );
  FA1A U7553 ( .CI(n8702), .A(n8651), .B(n8649), .S(n8704), .CO(n8705) );
  FA1A U7554 ( .CI(n8655), .A(n8704), .B(n8653), .S(n8706), .CO(n8707) );
  IVP U7555 ( .A(n5790), .Z(n8708) );
  FA1A U7556 ( .CI(n4318), .A(n4254), .B(n8708), .S(n8709), .CO(n8710) );
  FA1A U7557 ( .CI(n8659), .A(n4382), .B(n5150), .S(n8711), .CO(n8712) );
  FA1A U7558 ( .CI(n5726), .A(n4446), .B(n5086), .S(n8713), .CO(n8714) );
  FA1A U7559 ( .CI(n5598), .A(n5662), .B(n5214), .S(n8715), .CO(n8716) );
  FA1A U7560 ( .CI(n5470), .A(n5534), .B(n5022), .S(n8717), .CO(n8718) );
  FA1A U7561 ( .CI(n5342), .A(n5406), .B(n4830), .S(n8719), .CO(n8720) );
  FA1A U7562 ( .CI(n4958), .A(n5278), .B(n4510), .S(n8721), .CO(n8722) );
  FA1A U7563 ( .CI(n4766), .A(n4894), .B(n4574), .S(n8723), .CO(n8724) );
  FA1A U7564 ( .CI(n8709), .A(n4702), .B(n4638), .S(n8725), .CO(n8726) );
  FA1A U7565 ( .CI(n8725), .A(n8723), .B(n8661), .S(n8727), .CO(n8728) );
  FA1A U7566 ( .CI(n8719), .A(n8721), .B(n8673), .S(n8729), .CO(n8730) );
  FA1A U7567 ( .CI(n8713), .A(n8711), .B(n8663), .S(n8731), .CO(n8732) );
  FA1A U7568 ( .CI(n8717), .A(n8715), .B(n8665), .S(n8733), .CO(n8734) );
  FA1A U7569 ( .CI(n8671), .A(n8675), .B(n8667), .S(n8735), .CO(n8736) );
  FA1A U7570 ( .CI(n8679), .A(n8677), .B(n8669), .S(n8737), .CO(n8738) );
  FA1A U7571 ( .CI(n8733), .A(n8735), .B(n8687), .S(n8739), .CO(n8740) );
  FA1A U7572 ( .CI(n8729), .A(n8727), .B(n8683), .S(n8741), .CO(n8742) );
  FA1A U7573 ( .CI(n8731), .A(n8685), .B(n8681), .S(n8743), .CO(n8744) );
  FA1A U7574 ( .CI(n8743), .A(n8689), .B(n8737), .S(n8745), .CO(n8746) );
  FA1A U7575 ( .CI(n8739), .A(n8741), .B(n8691), .S(n8747), .CO(n8748) );
  FA1A U7576 ( .CI(n8745), .A(n8695), .B(n8693), .S(n8749), .CO(n8750) );
  FA1A U7577 ( .CI(n8749), .A(n8747), .B(n8697), .S(n8751), .CO(n8752) );
  FA1A U7578 ( .CI(n8751), .A(n8701), .B(n8699), .S(n8753), .CO(n8754) );
  FA1A U7579 ( .CI(n8705), .A(n8753), .B(n8703), .S(n8755), .CO(n8756) );
  FA1A U7580 ( .CI(n4255), .A(n5791), .B(n5790), .S(n8757), .CO(n8758) );
  FA1A U7581 ( .CI(n8757), .A(n4319), .B(n5087), .S(n8759), .CO(n8760) );
  FA1A U7582 ( .CI(n4447), .A(n5727), .B(n4383), .S(n8761), .CO(n8762) );
  FA1A U7583 ( .CI(n5663), .A(n4511), .B(n5151), .S(n8763), .CO(n8764) );
  FA1A U7584 ( .CI(n5535), .A(n5599), .B(n4575), .S(n8765), .CO(n8766) );
  FA1A U7585 ( .CI(n4703), .A(n4639), .B(n5407), .S(n8767), .CO(n8768) );
  FA1A U7586 ( .CI(n5343), .A(n5471), .B(n4767), .S(n8769), .CO(n8770) );
  FA1A U7587 ( .CI(n5215), .A(n5279), .B(n4831), .S(n8771), .CO(n8772) );
  FA1A U7588 ( .CI(n4959), .A(n5023), .B(n4895), .S(n8773), .CO(n8774) );
  FA1A U7589 ( .CI(n8771), .A(n8773), .B(n8710), .S(n8775), .CO(n8776) );
  FA1A U7590 ( .CI(n8726), .A(n8769), .B(n8722), .S(n8777), .CO(n8778) );
  FA1A U7591 ( .CI(n8759), .A(n8767), .B(n8720), .S(n8779), .CO(n8780) );
  FA1A U7592 ( .CI(n8763), .A(n8761), .B(n8712), .S(n8781), .CO(n8782) );
  FA1A U7593 ( .CI(n8765), .A(n8724), .B(n8714), .S(n8783), .CO(n8784) );
  FA1A U7594 ( .CI(n8775), .A(n8716), .B(n8718), .S(n8785), .CO(n8786) );
  FA1A U7595 ( .CI(n8777), .A(n8783), .B(n8734), .S(n8787), .CO(n8788) );
  FA1A U7596 ( .CI(n8781), .A(n8779), .B(n8728), .S(n8789), .CO(n8790) );
  FA1A U7597 ( .CI(n8732), .A(n8736), .B(n8730), .S(n8791), .CO(n8792) );
  FA1A U7598 ( .CI(n8740), .A(n8738), .B(n8785), .S(n8793), .CO(n8794) );
  FA1A U7599 ( .CI(n8787), .A(n8789), .B(n8742), .S(n8795), .CO(n8796) );
  FA1A U7600 ( .CI(n8793), .A(n8791), .B(n8744), .S(n8797), .CO(n8798) );
  FA1A U7601 ( .CI(n8797), .A(n8748), .B(n8746), .S(n8799), .CO(n8800) );
  FA1A U7602 ( .CI(n8799), .A(n8750), .B(n8795), .S(n8801), .CO(n8802) );
  FA1A U7603 ( .CI(n8754), .A(n8801), .B(n8752), .S(n8803), .CO(n8804) );
  IVP U7604 ( .A(n5792), .Z(n8805) );
  FA1A U7605 ( .CI(n5088), .A(n4320), .B(n8805), .S(n8806), .CO(n8807) );
  FA1A U7606 ( .CI(n8758), .A(n5728), .B(n5152), .S(n8808), .CO(n8809) );
  FA1A U7607 ( .CI(n5664), .A(n4384), .B(n5024), .S(n8810), .CO(n8811) );
  FA1A U7608 ( .CI(n4512), .A(n4448), .B(n5216), .S(n8812), .CO(n8813) );
  FA1A U7609 ( .CI(n4640), .A(n4576), .B(n5280), .S(n8814), .CO(n8815) );
  FA1A U7610 ( .CI(n5536), .A(n5600), .B(n4704), .S(n8816), .CO(n8817) );
  FA1A U7611 ( .CI(n5408), .A(n5472), .B(n4768), .S(n8818), .CO(n8819) );
  FA1A U7612 ( .CI(n4960), .A(n5344), .B(n4832), .S(n8820), .CO(n8821) );
  FA1A U7613 ( .CI(n8760), .A(n8806), .B(n4896), .S(n8822), .CO(n8823) );
  FA1A U7614 ( .CI(n8818), .A(n8820), .B(n8772), .S(n8824), .CO(n8825) );
  FA1A U7615 ( .CI(n8808), .A(n8816), .B(n8770), .S(n8826), .CO(n8827) );
  FA1A U7616 ( .CI(n8812), .A(n8810), .B(n8762), .S(n8828), .CO(n8829) );
  FA1A U7617 ( .CI(n8814), .A(n8774), .B(n8764), .S(n8830), .CO(n8831) );
  FA1A U7618 ( .CI(n8822), .A(n8766), .B(n8768), .S(n8832), .CO(n8833) );
  FA1A U7619 ( .CI(n8832), .A(n8830), .B(n8776), .S(n8834), .CO(n8835) );
  FA1A U7620 ( .CI(n8828), .A(n8826), .B(n8778), .S(n8836), .CO(n8837) );
  FA1A U7621 ( .CI(n8824), .A(n8784), .B(n8780), .S(n8838), .CO(n8839) );
  FA1A U7622 ( .CI(n8834), .A(n8786), .B(n8782), .S(n8840), .CO(n8841) );
  FA1A U7623 ( .CI(n8836), .A(n8838), .B(n8788), .S(n8842), .CO(n8843) );
  FA1A U7624 ( .CI(n8840), .A(n8792), .B(n8790), .S(n8844), .CO(n8845) );
  FA1A U7625 ( .CI(n8844), .A(n8796), .B(n8794), .S(n8846), .CO(n8847) );
  FA1A U7626 ( .CI(n8846), .A(n8798), .B(n8842), .S(n8848), .CO(n8849) );
  FA1A U7627 ( .CI(n8848), .A(n8802), .B(n8800), .S(n8850), .CO(n8851) );
  FA1A U7628 ( .CI(n4321), .A(n5793), .B(n5792), .S(n8852), .CO(n8853) );
  FA1A U7629 ( .CI(n8852), .A(n4385), .B(n5089), .S(n8854), .CO(n8855) );
  FA1A U7630 ( .CI(n4513), .A(n5729), .B(n4449), .S(n8856), .CO(n8857) );
  FA1A U7631 ( .CI(n5665), .A(n4577), .B(n5217), .S(n8858), .CO(n8859) );
  FA1A U7632 ( .CI(n5537), .A(n5601), .B(n4641), .S(n8860), .CO(n8861) );
  FA1A U7633 ( .CI(n4769), .A(n4705), .B(n5473), .S(n8862), .CO(n8863) );
  FA1A U7634 ( .CI(n5345), .A(n5409), .B(n4833), .S(n8864), .CO(n8865) );
  FA1A U7635 ( .CI(n5153), .A(n5281), .B(n4897), .S(n8866), .CO(n8867) );
  FA1A U7636 ( .CI(n8807), .A(n5025), .B(n4961), .S(n8868), .CO(n8869) );
  FA1A U7637 ( .CI(n8864), .A(n8866), .B(n8819), .S(n8870), .CO(n8871) );
  FA1A U7638 ( .CI(n8854), .A(n8862), .B(n8817), .S(n8872), .CO(n8873) );
  FA1A U7639 ( .CI(n8858), .A(n8856), .B(n8809), .S(n8874), .CO(n8875) );
  FA1A U7640 ( .CI(n8860), .A(n8821), .B(n8811), .S(n8876), .CO(n8877) );
  FA1A U7641 ( .CI(n8868), .A(n8813), .B(n8815), .S(n8878), .CO(n8879) );
  FA1A U7642 ( .CI(n8878), .A(n8829), .B(n8823), .S(n8880), .CO(n8881) );
  FA1A U7643 ( .CI(n8833), .A(n8870), .B(n8831), .S(n8882), .CO(n8883) );
  FA1A U7644 ( .CI(n8872), .A(n8874), .B(n8825), .S(n8884), .CO(n8885) );
  FA1A U7645 ( .CI(n8880), .A(n8876), .B(n8827), .S(n8886), .CO(n8887) );
  FA1A U7646 ( .CI(n8882), .A(n8884), .B(n8835), .S(n8888), .CO(n8889) );
  FA1A U7647 ( .CI(n8886), .A(n8839), .B(n8837), .S(n8890), .CO(n8891) );
  FA1A U7648 ( .CI(n8843), .A(n8888), .B(n8841), .S(n8892), .CO(n8893) );
  FA1A U7649 ( .CI(n8892), .A(n8845), .B(n8890), .S(n8894), .CO(n8895) );
  FA1A U7650 ( .CI(n8849), .A(n8894), .B(n8847), .S(n8896), .CO(n8897) );
  IVP U7651 ( .A(n5794), .Z(n8898) );
  FA1A U7652 ( .CI(n4450), .A(n4386), .B(n8898), .S(n8899), .CO(n8900) );
  FA1A U7653 ( .CI(n8853), .A(n5730), .B(n5154), .S(n8901), .CO(n8902) );
  FA1A U7654 ( .CI(n4578), .A(n4514), .B(n5218), .S(n8903), .CO(n8904) );
  FA1A U7655 ( .CI(n5666), .A(n4642), .B(n5282), .S(n8905), .CO(n8906) );
  FA1A U7656 ( .CI(n4770), .A(n4706), .B(n5538), .S(n8907), .CO(n8908) );
  FA1A U7657 ( .CI(n5474), .A(n5602), .B(n4834), .S(n8909), .CO(n8910) );
  FA1A U7658 ( .CI(n5346), .A(n5410), .B(n4898), .S(n8911), .CO(n8912) );
  FA1A U7659 ( .CI(n5026), .A(n5090), .B(n4962), .S(n8913), .CO(n8914) );
  FA1A U7660 ( .CI(n8913), .A(n8867), .B(n8899), .S(n8915), .CO(n8916) );
  FA1A U7661 ( .CI(n8903), .A(n8911), .B(n8863), .S(n8917), .CO(n8918) );
  FA1A U7662 ( .CI(n8905), .A(n8901), .B(n8855), .S(n8919), .CO(n8920) );
  FA1A U7663 ( .CI(n8907), .A(n8909), .B(n8857), .S(n8921), .CO(n8922) );
  FA1A U7664 ( .CI(n8861), .A(n8865), .B(n8859), .S(n8923), .CO(n8924) );
  FA1A U7665 ( .CI(n8871), .A(n8915), .B(n8869), .S(n8925), .CO(n8926) );
  FA1A U7666 ( .CI(n8879), .A(n8919), .B(n8877), .S(n8927), .CO(n8928) );
  FA1A U7667 ( .CI(n8917), .A(n8921), .B(n8873), .S(n8929), .CO(n8930) );
  FA1A U7668 ( .CI(n8925), .A(n8923), .B(n8875), .S(n8931), .CO(n8932) );
  FA1A U7669 ( .CI(n8931), .A(n8929), .B(n8881), .S(n8933), .CO(n8934) );
  FA1A U7670 ( .CI(n8887), .A(n8927), .B(n8883), .S(n8935), .CO(n8936) );
  FA1A U7671 ( .CI(n8889), .A(n8933), .B(n8885), .S(n8937), .CO(n8938) );
  FA1A U7672 ( .CI(n8937), .A(n8935), .B(n8891), .S(n8939), .CO(n8940) );
  FA1A U7673 ( .CI(n8895), .A(n8939), .B(n8893), .S(n8941), .CO(n8942) );
  FA1A U7674 ( .CI(n4387), .A(n5795), .B(n5794), .S(n8943), .CO(n8944) );
  FA1A U7675 ( .CI(n8943), .A(n5731), .B(n5155), .S(n8945), .CO(n8946) );
  FA1A U7676 ( .CI(n4515), .A(n5667), .B(n4451), .S(n8947), .CO(n8948) );
  FA1A U7677 ( .CI(n4643), .A(n4579), .B(n5091), .S(n8949), .CO(n8950) );
  FA1A U7678 ( .CI(n5539), .A(n5603), .B(n4707), .S(n8951), .CO(n8952) );
  FA1A U7679 ( .CI(n5475), .A(n4771), .B(n5027), .S(n8953), .CO(n8954) );
  FA1A U7680 ( .CI(n5347), .A(n5411), .B(n4835), .S(n8955), .CO(n8956) );
  FA1A U7681 ( .CI(n5219), .A(n5283), .B(n4899), .S(n8957), .CO(n8958) );
  FA1A U7682 ( .CI(n8902), .A(n8900), .B(n4963), .S(n8959), .CO(n8960) );
  FA1A U7683 ( .CI(n8955), .A(n8957), .B(n8914), .S(n8961), .CO(n8962) );
  FA1A U7684 ( .CI(n8945), .A(n8953), .B(n8910), .S(n8963), .CO(n8964) );
  FA1A U7685 ( .CI(n8949), .A(n8947), .B(n8904), .S(n8965), .CO(n8966) );
  FA1A U7686 ( .CI(n8951), .A(n8908), .B(n8912), .S(n8967), .CO(n8968) );
  FA1A U7687 ( .CI(n8916), .A(n8959), .B(n8906), .S(n8969), .CO(n8970) );
  FA1A U7688 ( .CI(n8961), .A(n8967), .B(n8922), .S(n8971), .CO(n8972) );
  FA1A U7689 ( .CI(n8965), .A(n8963), .B(n8918), .S(n8973), .CO(n8974) );
  FA1A U7690 ( .CI(n8969), .A(n8924), .B(n8920), .S(n8975), .CO(n8976) );
  FA1A U7691 ( .CI(n8975), .A(n8928), .B(n8926), .S(n8977), .CO(n8978) );
  FA1A U7692 ( .CI(n8932), .A(n8971), .B(n8930), .S(n8979), .CO(n8980) );
  FA1A U7693 ( .CI(n8934), .A(n8977), .B(n8973), .S(n8981), .CO(n8982) );
  FA1A U7694 ( .CI(n8981), .A(n8979), .B(n8936), .S(n8983), .CO(n8984) );
  FA1A U7695 ( .CI(n8940), .A(n8983), .B(n8938), .S(n8985), .CO(n8986) );
  IVP U7696 ( .A(n5796), .Z(n8987) );
  FA1A U7697 ( .CI(n4516), .A(n4452), .B(n8987), .S(n8988), .CO(n8989) );
  FA1A U7698 ( .CI(n8944), .A(n4580), .B(n5220), .S(n8990), .CO(n8991) );
  FA1A U7699 ( .CI(n4708), .A(n4644), .B(n5284), .S(n8992), .CO(n8993) );
  FA1A U7700 ( .CI(n5668), .A(n5732), .B(n5348), .S(n8994), .CO(n8995) );
  FA1A U7701 ( .CI(n4836), .A(n4772), .B(n5604), .S(n8996), .CO(n8997) );
  FA1A U7702 ( .CI(n5476), .A(n5540), .B(n4900), .S(n8998), .CO(n8999) );
  FA1A U7703 ( .CI(n5156), .A(n5412), .B(n4964), .S(n9000), .CO(n9001) );
  FA1A U7704 ( .CI(n8988), .A(n5092), .B(n5028), .S(n9002), .CO(n9003) );
  FA1A U7705 ( .CI(n9002), .A(n9000), .B(n8956), .S(n9004), .CO(n9005) );
  FA1A U7706 ( .CI(n8996), .A(n8998), .B(n8946), .S(n9006), .CO(n9007) );
  FA1A U7707 ( .CI(n8992), .A(n8994), .B(n8948), .S(n9008), .CO(n9009) );
  FA1A U7708 ( .CI(n8990), .A(n8958), .B(n8950), .S(n9010), .CO(n9011) );
  FA1A U7709 ( .CI(n8960), .A(n8954), .B(n8952), .S(n9012), .CO(n9013) );
  FA1A U7710 ( .CI(n9012), .A(n9010), .B(n8966), .S(n9014), .CO(n9015) );
  FA1A U7711 ( .CI(n9006), .A(n9008), .B(n8962), .S(n9016), .CO(n9017) );
  FA1A U7712 ( .CI(n9004), .A(n8968), .B(n8964), .S(n9018), .CO(n9019) );
  FA1A U7713 ( .CI(n9014), .A(n8972), .B(n8970), .S(n9020), .CO(n9021) );
  FA1A U7714 ( .CI(n8976), .A(n9016), .B(n8974), .S(n9022), .CO(n9023) );
  FA1A U7715 ( .CI(n8978), .A(n9020), .B(n9018), .S(n9024), .CO(n9025) );
  FA1A U7716 ( .CI(n9024), .A(n9022), .B(n8980), .S(n9026), .CO(n9027) );
  FA1A U7717 ( .CI(n9026), .A(n8984), .B(n8982), .S(n9028), .CO(n9029) );
  FA1A U7718 ( .CI(n4453), .A(n5797), .B(n5796), .S(n9030), .CO(n9031) );
  FA1A U7719 ( .CI(n9030), .A(n5733), .B(n5157), .S(n9032), .CO(n9033) );
  FA1A U7720 ( .CI(n4517), .A(n5669), .B(n5093), .S(n9034), .CO(n9035) );
  FA1A U7721 ( .CI(n5605), .A(n4581), .B(n5221), .S(n9036), .CO(n9037) );
  FA1A U7722 ( .CI(n4709), .A(n5541), .B(n4645), .S(n9038), .CO(n9039) );
  FA1A U7723 ( .CI(n5413), .A(n5477), .B(n5029), .S(n9040), .CO(n9041) );
  FA1A U7724 ( .CI(n5285), .A(n5349), .B(n4773), .S(n9042), .CO(n9043) );
  FA1A U7725 ( .CI(n4901), .A(n4965), .B(n4837), .S(n9044), .CO(n9045) );
  FA1A U7726 ( .CI(n9042), .A(n9044), .B(n8989), .S(n9046), .CO(n9047) );
  FA1A U7727 ( .CI(n9003), .A(n9034), .B(n8991), .S(n9048), .CO(n9049) );
  FA1A U7728 ( .CI(n9038), .A(n9040), .B(n8993), .S(n9050), .CO(n9051) );
  FA1A U7729 ( .CI(n9036), .A(n9032), .B(n8995), .S(n9052), .CO(n9053) );
  FA1A U7730 ( .CI(n8999), .A(n9001), .B(n8997), .S(n9054), .CO(n9055) );
  FA1A U7731 ( .CI(n9013), .A(n9054), .B(n9046), .S(n9056), .CO(n9057) );
  FA1A U7732 ( .CI(n9050), .A(n9052), .B(n9005), .S(n9058), .CO(n9059) );
  FA1A U7733 ( .CI(n9048), .A(n9011), .B(n9007), .S(n9060), .CO(n9061) );
  FA1A U7734 ( .CI(n9015), .A(n9056), .B(n9009), .S(n9062), .CO(n9063) );
  FA1A U7735 ( .CI(n9060), .A(n9058), .B(n9017), .S(n9064), .CO(n9065) );
  FA1A U7736 ( .CI(n9021), .A(n9062), .B(n9019), .S(n9066), .CO(n9067) );
  FA1A U7737 ( .CI(n9066), .A(n9064), .B(n9023), .S(n9068), .CO(n9069) );
  FA1A U7738 ( .CI(n9027), .A(n9068), .B(n9025), .S(n9070), .CO(n9071) );
  IVP U7739 ( .A(n5798), .Z(n9072) );
  FA1A U7740 ( .CI(n4582), .A(n4518), .B(n9072), .S(n9073), .CO(n9074) );
  FA1A U7741 ( .CI(n9031), .A(n4646), .B(n5286), .S(n9075), .CO(n9076) );
  FA1A U7742 ( .CI(n4774), .A(n4710), .B(n5350), .S(n9077), .CO(n9078) );
  FA1A U7743 ( .CI(n4902), .A(n4838), .B(n5414), .S(n9079), .CO(n9080) );
  FA1A U7744 ( .CI(n5670), .A(n4966), .B(n5734), .S(n9081), .CO(n9082) );
  FA1A U7745 ( .CI(n5542), .A(n5606), .B(n5030), .S(n9083), .CO(n9084) );
  FA1A U7746 ( .CI(n5222), .A(n5478), .B(n5094), .S(n9085), .CO(n9086) );
  FA1A U7747 ( .CI(n9033), .A(n9073), .B(n5158), .S(n9087), .CO(n9088) );
  FA1A U7748 ( .CI(n9075), .A(n9085), .B(n9043), .S(n9089), .CO(n9090) );
  FA1A U7749 ( .CI(n9081), .A(n9083), .B(n9035), .S(n9091), .CO(n9092) );
  FA1A U7750 ( .CI(n9079), .A(n9077), .B(n9037), .S(n9093), .CO(n9094) );
  FA1A U7751 ( .CI(n9041), .A(n9045), .B(n9039), .S(n9095), .CO(n9096) );
  FA1A U7752 ( .CI(n9095), .A(n9047), .B(n9087), .S(n9097), .CO(n9098) );
  FA1A U7753 ( .CI(n9091), .A(n9093), .B(n9049), .S(n9099), .CO(n9100) );
  FA1A U7754 ( .CI(n9089), .A(n9055), .B(n9051), .S(n9101), .CO(n9102) );
  FA1A U7755 ( .CI(n9057), .A(n9097), .B(n9053), .S(n9103), .CO(n9104) );
  FA1A U7756 ( .CI(n9101), .A(n9099), .B(n9059), .S(n9105), .CO(n9106) );
  FA1A U7757 ( .CI(n9063), .A(n9103), .B(n9061), .S(n9107), .CO(n9108) );
  FA1A U7758 ( .CI(n9107), .A(n9105), .B(n9065), .S(n9109), .CO(n9110) );
  FA1A U7759 ( .CI(n9069), .A(n9109), .B(n9067), .S(n9111), .CO(n9112) );
  FA1A U7760 ( .CI(n4519), .A(n5799), .B(n5798), .S(n9113), .CO(n9114) );
  FA1A U7761 ( .CI(n9113), .A(n5735), .B(n5223), .S(n9115), .CO(n9116) );
  FA1A U7762 ( .CI(n4647), .A(n5671), .B(n4583), .S(n9117), .CO(n9118) );
  FA1A U7763 ( .CI(n5543), .A(n5607), .B(n5159), .S(n9119), .CO(n9120) );
  FA1A U7764 ( .CI(n4775), .A(n5479), .B(n4711), .S(n9121), .CO(n9122) );
  FA1A U7765 ( .CI(n5351), .A(n5415), .B(n5095), .S(n9123), .CO(n9124) );
  FA1A U7766 ( .CI(n5031), .A(n5287), .B(n4839), .S(n9125), .CO(n9126) );
  FA1A U7767 ( .CI(n9074), .A(n4967), .B(n4903), .S(n9127), .CO(n9128) );
  FA1A U7768 ( .CI(n9115), .A(n9125), .B(n9084), .S(n9129), .CO(n9130) );
  FA1A U7769 ( .CI(n9121), .A(n9123), .B(n9076), .S(n9131), .CO(n9132) );
  FA1A U7770 ( .CI(n9119), .A(n9117), .B(n9078), .S(n9133), .CO(n9134) );
  FA1A U7771 ( .CI(n9082), .A(n9086), .B(n9080), .S(n9135), .CO(n9136) );
  FA1A U7772 ( .CI(n9090), .A(n9088), .B(n9127), .S(n9137), .CO(n9138) );
  FA1A U7773 ( .CI(n9133), .A(n9135), .B(n9096), .S(n9139), .CO(n9140) );
  FA1A U7774 ( .CI(n9131), .A(n9129), .B(n9092), .S(n9141), .CO(n9142) );
  FA1A U7775 ( .CI(n9098), .A(n9137), .B(n9094), .S(n9143), .CO(n9144) );
  FA1A U7776 ( .CI(n9141), .A(n9139), .B(n9100), .S(n9145), .CO(n9146) );
  FA1A U7777 ( .CI(n9104), .A(n9143), .B(n9102), .S(n9147), .CO(n9148) );
  FA1A U7778 ( .CI(n9147), .A(n9145), .B(n9106), .S(n9149), .CO(n9150) );
  FA1A U7779 ( .CI(n9110), .A(n9149), .B(n9108), .S(n9151), .CO(n9152) );
  IVP U7780 ( .A(n5800), .Z(n9153) );
  FA1A U7781 ( .CI(n4648), .A(n4584), .B(n9153), .S(n9154), .CO(n9155) );
  FA1A U7782 ( .CI(n9114), .A(n5736), .B(n5288), .S(n9156), .CO(n9157) );
  FA1A U7783 ( .CI(n5672), .A(n4712), .B(n5224), .S(n9158), .CO(n9159) );
  FA1A U7784 ( .CI(n5608), .A(n4776), .B(n5160), .S(n9160), .CO(n9161) );
  FA1A U7785 ( .CI(n5480), .A(n5544), .B(n5096), .S(n9162), .CO(n9163) );
  FA1A U7786 ( .CI(n5352), .A(n5416), .B(n4840), .S(n9164), .CO(n9165) );
  FA1A U7787 ( .CI(n4968), .A(n5032), .B(n4904), .S(n9166), .CO(n9167) );
  FA1A U7788 ( .CI(n9166), .A(n9126), .B(n9154), .S(n9168), .CO(n9169) );
  FA1A U7789 ( .CI(n9162), .A(n9164), .B(n9116), .S(n9170), .CO(n9171) );
  FA1A U7790 ( .CI(n9158), .A(n9160), .B(n9122), .S(n9172), .CO(n9173) );
  FA1A U7791 ( .CI(n9156), .A(n9124), .B(n9118), .S(n9174), .CO(n9175) );
  FA1A U7792 ( .CI(n9168), .A(n9128), .B(n9120), .S(n9176), .CO(n9177) );
  FA1A U7793 ( .CI(n9176), .A(n9174), .B(n9130), .S(n9178), .CO(n9179) );
  FA1A U7794 ( .CI(n9170), .A(n9172), .B(n9132), .S(n9180), .CO(n9181) );
  FA1A U7795 ( .CI(n9138), .A(n9136), .B(n9134), .S(n9182), .CO(n9183) );
  FA1A U7796 ( .CI(n9182), .A(n9178), .B(n9140), .S(n9184), .CO(n9185) );
  FA1A U7797 ( .CI(n9144), .A(n9180), .B(n9142), .S(n9186), .CO(n9187) );
  FA1A U7798 ( .CI(n9186), .A(n9184), .B(n9146), .S(n9188), .CO(n9189) );
  FA1A U7799 ( .CI(n9150), .A(n9188), .B(n9148), .S(n9190), .CO(n9191) );
  FA1A U7800 ( .CI(n4585), .A(n5801), .B(n5800), .S(n9192), .CO(n9193) );
  FA1A U7801 ( .CI(n9192), .A(n4649), .B(n5289), .S(n9194), .CO(n9195) );
  FA1A U7802 ( .CI(n4777), .A(n5737), .B(n4713), .S(n9196), .CO(n9197) );
  FA1A U7803 ( .CI(n5673), .A(n4841), .B(n5353), .S(n9198), .CO(n9199) );
  FA1A U7804 ( .CI(n5545), .A(n5609), .B(n4905), .S(n9200), .CO(n9201) );
  FA1A U7805 ( .CI(n5417), .A(n5481), .B(n4969), .S(n9202), .CO(n9203) );
  FA1A U7806 ( .CI(n5161), .A(n5225), .B(n5033), .S(n9204), .CO(n9205) );
  FA1A U7807 ( .CI(n9157), .A(n9155), .B(n5097), .S(n9206), .CO(n9207) );
  FA1A U7808 ( .CI(n9202), .A(n9204), .B(n9167), .S(n9208), .CO(n9209) );
  FA1A U7809 ( .CI(n9198), .A(n9200), .B(n9163), .S(n9210), .CO(n9211) );
  FA1A U7810 ( .CI(n9194), .A(n9196), .B(n9159), .S(n9212), .CO(n9213) );
  FA1A U7811 ( .CI(n9206), .A(n9165), .B(n9161), .S(n9214), .CO(n9215) );
  FA1A U7812 ( .CI(n9214), .A(n9212), .B(n9169), .S(n9216), .CO(n9217) );
  FA1A U7813 ( .CI(n9177), .A(n9210), .B(n9171), .S(n9218), .CO(n9219) );
  FA1A U7814 ( .CI(n9208), .A(n9175), .B(n9173), .S(n9220), .CO(n9221) );
  FA1A U7815 ( .CI(n9183), .A(n9220), .B(n9216), .S(n9222), .CO(n9223) );
  FA1A U7816 ( .CI(n9218), .A(n9181), .B(n9179), .S(n9224), .CO(n9225) );
  FA1A U7817 ( .CI(n9187), .A(n9224), .B(n9222), .S(n9226), .CO(n9227) );
  FA1A U7818 ( .CI(n9189), .A(n9226), .B(n9185), .S(n9228), .CO(n9229) );
  IVP U7819 ( .A(n5802), .Z(n9230) );
  FA1A U7820 ( .CI(n4714), .A(n4650), .B(n9230), .S(n9231), .CO(n9232) );
  FA1A U7821 ( .CI(n9193), .A(n5738), .B(n5354), .S(n9233), .CO(n9234) );
  FA1A U7822 ( .CI(n4778), .A(n5674), .B(n5226), .S(n9235), .CO(n9236) );
  FA1A U7823 ( .CI(n4842), .A(n5610), .B(n5290), .S(n9237), .CO(n9238) );
  FA1A U7824 ( .CI(n5482), .A(n5546), .B(n4906), .S(n9239), .CO(n9240) );
  FA1A U7825 ( .CI(n5162), .A(n5418), .B(n4970), .S(n9241), .CO(n9242) );
  FA1A U7826 ( .CI(n9231), .A(n5098), .B(n5034), .S(n9243), .CO(n9244) );
  FA1A U7827 ( .CI(n9243), .A(n9241), .B(n9195), .S(n9245), .CO(n9246) );
  FA1A U7828 ( .CI(n9237), .A(n9239), .B(n9203), .S(n9247), .CO(n9248) );
  FA1A U7829 ( .CI(n9235), .A(n9233), .B(n9197), .S(n9249), .CO(n9250) );
  FA1A U7830 ( .CI(n9201), .A(n9205), .B(n9199), .S(n9251), .CO(n9252) );
  FA1A U7831 ( .CI(n9249), .A(n9251), .B(n9207), .S(n9253), .CO(n9254) );
  FA1A U7832 ( .CI(n9215), .A(n9247), .B(n9209), .S(n9255), .CO(n9256) );
  FA1A U7833 ( .CI(n9245), .A(n9213), .B(n9211), .S(n9257), .CO(n9258) );
  FA1A U7834 ( .CI(n9255), .A(n9257), .B(n9253), .S(n9259), .CO(n9260) );
  FA1A U7835 ( .CI(n9219), .A(n9221), .B(n9217), .S(n9261), .CO(n9262) );
  FA1A U7836 ( .CI(n9225), .A(n9261), .B(n9259), .S(n9263), .CO(n9264) );
  FA1A U7837 ( .CI(n9227), .A(n9263), .B(n9223), .S(n9265), .CO(n9266) );
  FA1A U7838 ( .CI(n4651), .A(n5803), .B(n5802), .S(n9267), .CO(n9268) );
  FA1A U7839 ( .CI(n9267), .A(n5739), .B(n5291), .S(n9269), .CO(n9270) );
  FA1A U7840 ( .CI(n4779), .A(n4715), .B(n5227), .S(n9271), .CO(n9272) );
  FA1A U7841 ( .CI(n5611), .A(n5675), .B(n4843), .S(n9273), .CO(n9274) );
  FA1A U7842 ( .CI(n4971), .A(n4907), .B(n5547), .S(n9275), .CO(n9276) );
  FA1A U7843 ( .CI(n5419), .A(n5483), .B(n5035), .S(n9277), .CO(n9278) );
  FA1A U7844 ( .CI(n5163), .A(n5355), .B(n5099), .S(n9279), .CO(n9280) );
  FA1A U7845 ( .CI(n9277), .A(n9279), .B(n9232), .S(n9281), .CO(n9282) );
  FA1A U7846 ( .CI(n9244), .A(n9275), .B(n9240), .S(n9283), .CO(n9284) );
  FA1A U7847 ( .CI(n9269), .A(n9273), .B(n9238), .S(n9285), .CO(n9286) );
  FA1A U7848 ( .CI(n9271), .A(n9242), .B(n9234), .S(n9287), .CO(n9288) );
  FA1A U7849 ( .CI(n9246), .A(n9281), .B(n9236), .S(n9289), .CO(n9290) );
  FA1A U7850 ( .CI(n9285), .A(n9287), .B(n9248), .S(n9291), .CO(n9292) );
  FA1A U7851 ( .CI(n9283), .A(n9252), .B(n9250), .S(n9293), .CO(n9294) );
  FA1A U7852 ( .CI(n9293), .A(n9254), .B(n9289), .S(n9295), .CO(n9296) );
  FA1A U7853 ( .CI(n9291), .A(n9258), .B(n9256), .S(n9297), .CO(n9298) );
  FA1A U7854 ( .CI(n9297), .A(n9262), .B(n9295), .S(n9299), .CO(n9300) );
  FA1A U7855 ( .CI(n9264), .A(n9299), .B(n9260), .S(n9301), .CO(n9302) );
  IVP U7856 ( .A(n5804), .Z(n9303) );
  FA1A U7857 ( .CI(n4780), .A(n4716), .B(n9303), .S(n9304), .CO(n9305) );
  FA1A U7858 ( .CI(n9268), .A(n4844), .B(n5356), .S(n9306), .CO(n9307) );
  FA1A U7859 ( .CI(n5740), .A(n4908), .B(n5420), .S(n9308), .CO(n9309) );
  FA1A U7860 ( .CI(n4972), .A(n5676), .B(n5292), .S(n9310), .CO(n9311) );
  FA1A U7861 ( .CI(n5548), .A(n5612), .B(n5036), .S(n9312), .CO(n9313) );
  FA1A U7862 ( .CI(n5228), .A(n5484), .B(n5100), .S(n9314), .CO(n9315) );
  FA1A U7863 ( .CI(n9270), .A(n9304), .B(n5164), .S(n9316), .CO(n9317) );
  FA1A U7864 ( .CI(n9312), .A(n9314), .B(n9278), .S(n9318), .CO(n9319) );
  FA1A U7865 ( .CI(n9306), .A(n9310), .B(n9276), .S(n9320), .CO(n9321) );
  FA1A U7866 ( .CI(n9308), .A(n9280), .B(n9272), .S(n9322), .CO(n9323) );
  FA1A U7867 ( .CI(n9282), .A(n9316), .B(n9274), .S(n9324), .CO(n9325) );
  FA1A U7868 ( .CI(n9320), .A(n9322), .B(n9284), .S(n9326), .CO(n9327) );
  FA1A U7869 ( .CI(n9318), .A(n9288), .B(n9286), .S(n9328), .CO(n9329) );
  FA1A U7870 ( .CI(n9328), .A(n9290), .B(n9324), .S(n9330), .CO(n9331) );
  FA1A U7871 ( .CI(n9326), .A(n9294), .B(n9292), .S(n9332), .CO(n9333) );
  FA1A U7872 ( .CI(n9332), .A(n9296), .B(n9330), .S(n9334), .CO(n9335) );
  FA1A U7873 ( .CI(n9300), .A(n9334), .B(n9298), .S(n9336), .CO(n9337) );
  FA1A U7874 ( .CI(n4717), .A(n5805), .B(n5804), .S(n9338), .CO(n9339) );
  FA1A U7875 ( .CI(n9338), .A(n5741), .B(n5293), .S(n9340), .CO(n9341) );
  FA1A U7876 ( .CI(n4781), .A(n5677), .B(n5229), .S(n9342), .CO(n9343) );
  FA1A U7877 ( .CI(n5549), .A(n5613), .B(n4845), .S(n9344), .CO(n9345) );
  FA1A U7878 ( .CI(n5421), .A(n4909), .B(n5485), .S(n9346), .CO(n9347) );
  FA1A U7879 ( .CI(n5165), .A(n5357), .B(n4973), .S(n9348), .CO(n9349) );
  FA1A U7880 ( .CI(n9305), .A(n5101), .B(n5037), .S(n9350), .CO(n9351) );
  FA1A U7881 ( .CI(n9346), .A(n9348), .B(n9313), .S(n9352), .CO(n9353) );
  FA1A U7882 ( .CI(n9340), .A(n9344), .B(n9311), .S(n9354), .CO(n9355) );
  FA1A U7883 ( .CI(n9342), .A(n9315), .B(n9307), .S(n9356), .CO(n9357) );
  FA1A U7884 ( .CI(n9317), .A(n9350), .B(n9309), .S(n9358), .CO(n9359) );
  FA1A U7885 ( .CI(n9358), .A(n9356), .B(n9319), .S(n9360), .CO(n9361) );
  FA1A U7886 ( .CI(n9354), .A(n9352), .B(n9321), .S(n9362), .CO(n9363) );
  FA1A U7887 ( .CI(n9327), .A(n9325), .B(n9323), .S(n9364), .CO(n9365) );
  FA1A U7888 ( .CI(n9362), .A(n9360), .B(n9329), .S(n9366), .CO(n9367) );
  FA1A U7889 ( .CI(n9366), .A(n9331), .B(n9364), .S(n9368), .CO(n9369) );
  FA1A U7890 ( .CI(n9335), .A(n9368), .B(n9333), .S(n9370), .CO(n9371) );
  IVP U7891 ( .A(n5806), .Z(n9372) );
  FA1A U7892 ( .CI(n4846), .A(n4782), .B(n9372), .S(n9373), .CO(n9374) );
  FA1A U7893 ( .CI(n9339), .A(n5742), .B(n5422), .S(n9375), .CO(n9376) );
  FA1A U7894 ( .CI(n5678), .A(n4910), .B(n5294), .S(n9377), .CO(n9378) );
  FA1A U7895 ( .CI(n5038), .A(n4974), .B(n5550), .S(n9379), .CO(n9380) );
  FA1A U7896 ( .CI(n5486), .A(n5614), .B(n5102), .S(n9381), .CO(n9382) );
  FA1A U7897 ( .CI(n5358), .A(n5230), .B(n5166), .S(n9383), .CO(n9384) );
  FA1A U7898 ( .CI(n9383), .A(n9349), .B(n9373), .S(n9385), .CO(n9386) );
  FA1A U7899 ( .CI(n9377), .A(n9381), .B(n9345), .S(n9387), .CO(n9388) );
  FA1A U7900 ( .CI(n9379), .A(n9375), .B(n9341), .S(n9389), .CO(n9390) );
  FA1A U7901 ( .CI(n9351), .A(n9347), .B(n9343), .S(n9391), .CO(n9392) );
  FA1A U7902 ( .CI(n9391), .A(n9389), .B(n9385), .S(n9393), .CO(n9394) );
  FA1A U7903 ( .CI(n9359), .A(n9387), .B(n9353), .S(n9395), .CO(n9396) );
  FA1A U7904 ( .CI(n9393), .A(n9357), .B(n9355), .S(n9397), .CO(n9398) );
  FA1A U7905 ( .CI(n9397), .A(n9395), .B(n9361), .S(n9399), .CO(n9400) );
  FA1A U7906 ( .CI(n9367), .A(n9365), .B(n9363), .S(n9401), .CO(n9402) );
  FA1A U7907 ( .CI(n9369), .A(n9401), .B(n9399), .S(n9403), .CO(n9404) );
  FA1A U7908 ( .CI(n4783), .A(n5807), .B(n5806), .S(n9405), .CO(n9406) );
  FA1A U7909 ( .CI(n9405), .A(n4847), .B(n5359), .S(n9407), .CO(n9408) );
  FA1A U7910 ( .CI(n4975), .A(n5743), .B(n4911), .S(n9409), .CO(n9410) );
  FA1A U7911 ( .CI(n5615), .A(n5679), .B(n5039), .S(n9411), .CO(n9412) );
  FA1A U7912 ( .CI(n5487), .A(n5551), .B(n5295), .S(n9413), .CO(n9414) );
  FA1A U7913 ( .CI(n5231), .A(n5423), .B(n5103), .S(n9415), .CO(n9416) );
  FA1A U7914 ( .CI(n9376), .A(n9374), .B(n5167), .S(n9417), .CO(n9418) );
  FA1A U7915 ( .CI(n9413), .A(n9415), .B(n9384), .S(n9419), .CO(n9420) );
  FA1A U7916 ( .CI(n9409), .A(n9407), .B(n9380), .S(n9421), .CO(n9422) );
  FA1A U7917 ( .CI(n9411), .A(n9382), .B(n9378), .S(n9423), .CO(n9424) );
  FA1A U7918 ( .CI(n9423), .A(n9386), .B(n9417), .S(n9425), .CO(n9426) );
  FA1A U7919 ( .CI(n9419), .A(n9421), .B(n9388), .S(n9427), .CO(n9428) );
  FA1A U7920 ( .CI(n9425), .A(n9392), .B(n9390), .S(n9429), .CO(n9430) );
  FA1A U7921 ( .CI(n9429), .A(n9427), .B(n9394), .S(n9431), .CO(n9432) );
  FA1A U7922 ( .CI(n9431), .A(n9398), .B(n9396), .S(n9433), .CO(n9434) );
  FA1A U7923 ( .CI(n9402), .A(n9433), .B(n9400), .S(n9435), .CO(n9436) );
  IVP U7924 ( .A(n5808), .Z(n9437) );
  FA1A U7925 ( .CI(n4912), .A(n4848), .B(n9437), .S(n9438), .CO(n9439) );
  FA1A U7926 ( .CI(n9406), .A(n4976), .B(n5424), .S(n9440), .CO(n9441) );
  FA1A U7927 ( .CI(n5744), .A(n5040), .B(n5360), .S(n9442), .CO(n9443) );
  FA1A U7928 ( .CI(n5616), .A(n5104), .B(n5680), .S(n9444), .CO(n9445) );
  FA1A U7929 ( .CI(n5488), .A(n5552), .B(n5168), .S(n9446), .CO(n9447) );
  FA1A U7930 ( .CI(n9438), .A(n5232), .B(n5296), .S(n9448), .CO(n9449) );
  FA1A U7931 ( .CI(n9448), .A(n9446), .B(n9414), .S(n9450), .CO(n9451) );
  FA1A U7932 ( .CI(n9442), .A(n9440), .B(n9408), .S(n9452), .CO(n9453) );
  FA1A U7933 ( .CI(n9444), .A(n9416), .B(n9410), .S(n9454), .CO(n9455) );
  FA1A U7934 ( .CI(n9420), .A(n9418), .B(n9412), .S(n9456), .CO(n9457) );
  FA1A U7935 ( .CI(n9450), .A(n9452), .B(n9422), .S(n9458), .CO(n9459) );
  FA1A U7936 ( .CI(n9456), .A(n9454), .B(n9424), .S(n9460), .CO(n9461) );
  FA1A U7937 ( .CI(n9460), .A(n9458), .B(n9426), .S(n9462), .CO(n9463) );
  FA1A U7938 ( .CI(n9462), .A(n9430), .B(n9428), .S(n9464), .CO(n9465) );
  FA1A U7939 ( .CI(n9434), .A(n9464), .B(n9432), .S(n9466), .CO(n9467) );
  FA1A U7940 ( .CI(n4849), .A(n5809), .B(n5808), .S(n9468), .CO(n9469) );
  FA1A U7941 ( .CI(n9468), .A(n5745), .B(n5361), .S(n9470), .CO(n9471) );
  FA1A U7942 ( .CI(n5681), .A(n4913), .B(n5297), .S(n9472), .CO(n9473) );
  FA1A U7943 ( .CI(n5041), .A(n5617), .B(n4977), .S(n9474), .CO(n9475) );
  FA1A U7944 ( .CI(n5489), .A(n5553), .B(n5105), .S(n9476), .CO(n9477) );
  FA1A U7945 ( .CI(n5233), .A(n5425), .B(n5169), .S(n9478), .CO(n9479) );
  FA1A U7946 ( .CI(n9476), .A(n9478), .B(n9439), .S(n9480), .CO(n9481) );
  FA1A U7947 ( .CI(n9449), .A(n9472), .B(n9441), .S(n9482), .CO(n9483) );
  FA1A U7948 ( .CI(n9474), .A(n9470), .B(n9443), .S(n9484), .CO(n9485) );
  FA1A U7949 ( .CI(n9480), .A(n9447), .B(n9445), .S(n9486), .CO(n9487) );
  FA1A U7950 ( .CI(n9482), .A(n9484), .B(n9451), .S(n9488), .CO(n9489) );
  FA1A U7951 ( .CI(n9486), .A(n9455), .B(n9453), .S(n9490), .CO(n9491) );
  FA1A U7952 ( .CI(n9490), .A(n9459), .B(n9457), .S(n9492), .CO(n9493) );
  FA1A U7953 ( .CI(n9492), .A(n9461), .B(n9488), .S(n9494), .CO(n9495) );
  FA1A U7954 ( .CI(n9465), .A(n9494), .B(n9463), .S(n9496), .CO(n9497) );
  IVP U7955 ( .A(n5810), .Z(n9498) );
  FA1A U7956 ( .CI(n4978), .A(n4914), .B(n9498), .S(n9499), .CO(n9500) );
  FA1A U7957 ( .CI(n9469), .A(n5746), .B(n5426), .S(n9501), .CO(n9502) );
  FA1A U7958 ( .CI(n5618), .A(n5682), .B(n5362), .S(n9503), .CO(n9504) );
  FA1A U7959 ( .CI(n5298), .A(n5490), .B(n5554), .S(n9505), .CO(n9506) );
  FA1A U7960 ( .CI(n5170), .A(n5234), .B(n5042), .S(n9507), .CO(n9508) );
  FA1A U7961 ( .CI(n9471), .A(n9499), .B(n5106), .S(n9509), .CO(n9510) );
  FA1A U7962 ( .CI(n9501), .A(n9507), .B(n9477), .S(n9511), .CO(n9512) );
  FA1A U7963 ( .CI(n9505), .A(n9503), .B(n9473), .S(n9513), .CO(n9514) );
  FA1A U7964 ( .CI(n9509), .A(n9479), .B(n9475), .S(n9515), .CO(n9516) );
  FA1A U7965 ( .CI(n9515), .A(n9513), .B(n9481), .S(n9517), .CO(n9518) );
  FA1A U7966 ( .CI(n9511), .A(n9485), .B(n9483), .S(n9519), .CO(n9520) );
  FA1A U7967 ( .CI(n9489), .A(n9517), .B(n9487), .S(n9521), .CO(n9522) );
  FA1A U7968 ( .CI(n9521), .A(n9491), .B(n9519), .S(n9523), .CO(n9524) );
  FA1A U7969 ( .CI(n9495), .A(n9523), .B(n9493), .S(n9525), .CO(n9526) );
  FA1A U7970 ( .CI(n4915), .A(n5811), .B(n5810), .S(n9527), .CO(n9528) );
  FA1A U7971 ( .CI(n9527), .A(n4979), .B(n5427), .S(n9529), .CO(n9530) );
  FA1A U7972 ( .CI(n5747), .A(n5043), .B(n5363), .S(n9531), .CO(n9532) );
  FA1A U7973 ( .CI(n5171), .A(n5683), .B(n5107), .S(n9533), .CO(n9534) );
  FA1A U7974 ( .CI(n5555), .A(n5619), .B(n5235), .S(n9535), .CO(n9536) );
  FA1A U7975 ( .CI(n9500), .A(n5491), .B(n5299), .S(n9537), .CO(n9538) );
  FA1A U7976 ( .CI(n9529), .A(n9535), .B(n9506), .S(n9539), .CO(n9540) );
  FA1A U7977 ( .CI(n9533), .A(n9531), .B(n9502), .S(n9541), .CO(n9542) );
  FA1A U7978 ( .CI(n9537), .A(n9508), .B(n9504), .S(n9543), .CO(n9544) );
  FA1A U7979 ( .CI(n9543), .A(n9512), .B(n9510), .S(n9545), .CO(n9546) );
  FA1A U7980 ( .CI(n9516), .A(n9539), .B(n9514), .S(n9547), .CO(n9548) );
  FA1A U7981 ( .CI(n9518), .A(n9545), .B(n9541), .S(n9549), .CO(n9550) );
  FA1A U7982 ( .CI(n9549), .A(n9547), .B(n9520), .S(n9551), .CO(n9552) );
  FA1A U7983 ( .CI(n9524), .A(n9551), .B(n9522), .S(n9553), .CO(n9554) );
  IVP U7984 ( .A(n5812), .Z(n9555) );
  FA1A U7985 ( .CI(n5044), .A(n4980), .B(n9555), .S(n9556), .CO(n9557) );
  FA1A U7986 ( .CI(n9528), .A(n5108), .B(n5492), .S(n9558), .CO(n9559) );
  FA1A U7987 ( .CI(n5684), .A(n5748), .B(n5556), .S(n9560), .CO(n9561) );
  FA1A U7988 ( .CI(n5428), .A(n5620), .B(n5172), .S(n9562), .CO(n9563) );
  FA1A U7989 ( .CI(n5300), .A(n5364), .B(n5236), .S(n9564), .CO(n9565) );
  FA1A U7990 ( .CI(n9564), .A(n9536), .B(n9556), .S(n9566), .CO(n9567) );
  FA1A U7991 ( .CI(n9560), .A(n9562), .B(n9530), .S(n9568), .CO(n9569) );
  FA1A U7992 ( .CI(n9558), .A(n9534), .B(n9532), .S(n9570), .CO(n9571) );
  FA1A U7993 ( .CI(n9540), .A(n9566), .B(n9538), .S(n9572), .CO(n9573) );
  FA1A U7994 ( .CI(n9544), .A(n9568), .B(n9542), .S(n9574), .CO(n9575) );
  FA1A U7995 ( .CI(n9546), .A(n9572), .B(n9570), .S(n9576), .CO(n9577) );
  FA1A U7996 ( .CI(n9576), .A(n9574), .B(n9548), .S(n9578), .CO(n9579) );
  FA1A U7997 ( .CI(n9552), .A(n9578), .B(n9550), .S(n9580), .CO(n9581) );
  FA1A U7998 ( .CI(n4981), .A(n5813), .B(n5812), .S(n9582), .CO(n9583) );
  FA1A U7999 ( .CI(n9582), .A(n5749), .B(n5429), .S(n9584), .CO(n9585) );
  FA1A U8000 ( .CI(n5621), .A(n5685), .B(n5365), .S(n9586), .CO(n9587) );
  FA1A U8001 ( .CI(n5493), .A(n5557), .B(n5045), .S(n9588), .CO(n9589) );
  FA1A U8002 ( .CI(n5237), .A(n5301), .B(n5109), .S(n9590), .CO(n9591) );
  FA1A U8003 ( .CI(n9559), .A(n9557), .B(n5173), .S(n9592), .CO(n9593) );
  FA1A U8004 ( .CI(n9588), .A(n9590), .B(n9565), .S(n9594), .CO(n9595) );
  FA1A U8005 ( .CI(n9586), .A(n9584), .B(n9561), .S(n9596), .CO(n9597) );
  FA1A U8006 ( .CI(n9567), .A(n9592), .B(n9563), .S(n9598), .CO(n9599) );
  FA1A U8007 ( .CI(n9596), .A(n9594), .B(n9569), .S(n9600), .CO(n9601) );
  FA1A U8008 ( .CI(n9573), .A(n9598), .B(n9571), .S(n9602), .CO(n9603) );
  FA1A U8009 ( .CI(n9602), .A(n9600), .B(n9575), .S(n9604), .CO(n9605) );
  FA1A U8010 ( .CI(n9579), .A(n9604), .B(n9577), .S(n9606), .CO(n9607) );
  IVP U8011 ( .A(n5814), .Z(n9608) );
  FA1A U8012 ( .CI(n5110), .A(n5046), .B(n9608), .S(n9609), .CO(n9610) );
  FA1A U8013 ( .CI(n9583), .A(n5750), .B(n5494), .S(n9611), .CO(n9612) );
  FA1A U8014 ( .CI(n5238), .A(n5174), .B(n5430), .S(n9613), .CO(n9614) );
  FA1A U8015 ( .CI(n5622), .A(n5686), .B(n5302), .S(n9615), .CO(n9616) );
  FA1A U8016 ( .CI(n9609), .A(n5558), .B(n5366), .S(n9617), .CO(n9618) );
  FA1A U8017 ( .CI(n9617), .A(n9615), .B(n9585), .S(n9619), .CO(n9620) );
  FA1A U8018 ( .CI(n9611), .A(n9613), .B(n9587), .S(n9621), .CO(n9622) );
  FA1A U8019 ( .CI(n9593), .A(n9591), .B(n9589), .S(n9623), .CO(n9624) );
  FA1A U8020 ( .CI(n9623), .A(n9619), .B(n9595), .S(n9625), .CO(n9626) );
  FA1A U8021 ( .CI(n9599), .A(n9621), .B(n9597), .S(n9627), .CO(n9628) );
  FA1A U8022 ( .CI(n9627), .A(n9625), .B(n9601), .S(n9629), .CO(n9630) );
  FA1A U8023 ( .CI(n9605), .A(n9629), .B(n9603), .S(n9631), .CO(n9632) );
  FA1A U8024 ( .CI(n5047), .A(n5815), .B(n5814), .S(n9633), .CO(n9634) );
  FA1A U8025 ( .CI(n9633), .A(n5111), .B(n5495), .S(n9635), .CO(n9636) );
  FA1A U8026 ( .CI(n5687), .A(n5751), .B(n5175), .S(n9637), .CO(n9638) );
  FA1A U8027 ( .CI(n5559), .A(n5239), .B(n5623), .S(n9639), .CO(n9640) );
  FA1A U8028 ( .CI(n5367), .A(n5431), .B(n5303), .S(n9641), .CO(n9642) );
  FA1A U8029 ( .CI(n9639), .A(n9641), .B(n9610), .S(n9643), .CO(n9644) );
  FA1A U8030 ( .CI(n9618), .A(n9637), .B(n9612), .S(n9645), .CO(n9646) );
  FA1A U8031 ( .CI(n9635), .A(n9616), .B(n9614), .S(n9647), .CO(n9648) );
  FA1A U8032 ( .CI(n9624), .A(n9647), .B(n9643), .S(n9649), .CO(n9650) );
  FA1A U8033 ( .CI(n9645), .A(n9622), .B(n9620), .S(n9651), .CO(n9652) );
  FA1A U8034 ( .CI(n9628), .A(n9651), .B(n9649), .S(n9653), .CO(n9654) );
  FA1A U8035 ( .CI(n9630), .A(n9653), .B(n9626), .S(n9655), .CO(n9656) );
  IVP U8036 ( .A(n5816), .Z(n9657) );
  FA1A U8037 ( .CI(n5176), .A(n5112), .B(n9657), .S(n9658), .CO(n9659) );
  FA1A U8038 ( .CI(n9634), .A(n5240), .B(n5560), .S(n9660), .CO(n9661) );
  FA1A U8039 ( .CI(n5304), .A(n5752), .B(n5624), .S(n9662), .CO(n9663) );
  FA1A U8040 ( .CI(n5496), .A(n5688), .B(n5368), .S(n9664), .CO(n9665) );
  FA1A U8041 ( .CI(n9636), .A(n9658), .B(n5432), .S(n9666), .CO(n9667) );
  FA1A U8042 ( .CI(n9662), .A(n9664), .B(n9638), .S(n9668), .CO(n9669) );
  FA1A U8043 ( .CI(n9660), .A(n9642), .B(n9640), .S(n9670), .CO(n9671) );
  FA1A U8044 ( .CI(n9670), .A(n9644), .B(n9666), .S(n9672), .CO(n9673) );
  FA1A U8045 ( .CI(n9668), .A(n9648), .B(n9646), .S(n9674), .CO(n9675) );
  FA1A U8046 ( .CI(n9674), .A(n9650), .B(n9672), .S(n9676), .CO(n9677) );
  FA1A U8047 ( .CI(n9654), .A(n9676), .B(n9652), .S(n9678), .CO(n9679) );
  FA1A U8048 ( .CI(n5113), .A(n5817), .B(n5816), .S(n9680), .CO(n9681) );
  FA1A U8049 ( .CI(n9680), .A(n5753), .B(n5497), .S(n9682), .CO(n9683) );
  FA1A U8050 ( .CI(n5625), .A(n5689), .B(n5177), .S(n9684), .CO(n9685) );
  FA1A U8051 ( .CI(n5433), .A(n5561), .B(n5369), .S(n9686), .CO(n9687) );
  FA1A U8052 ( .CI(n9659), .A(n5305), .B(n5241), .S(n9688), .CO(n9689) );
  FA1A U8053 ( .CI(n9684), .A(n9686), .B(n9661), .S(n9690), .CO(n9691) );
  FA1A U8054 ( .CI(n9682), .A(n9665), .B(n9663), .S(n9692), .CO(n9693) );
  FA1A U8055 ( .CI(n9669), .A(n9667), .B(n9688), .S(n9694), .CO(n9695) );
  FA1A U8056 ( .CI(n9692), .A(n9690), .B(n9671), .S(n9696), .CO(n9697) );
  FA1A U8057 ( .CI(n9696), .A(n9673), .B(n9694), .S(n9698), .CO(n9699) );
  FA1A U8058 ( .CI(n9677), .A(n9698), .B(n9675), .S(n9700), .CO(n9701) );
  IVP U8059 ( .A(n5818), .Z(n9702) );
  FA1A U8060 ( .CI(n5242), .A(n5178), .B(n9702), .S(n9703), .CO(n9704) );
  FA1A U8061 ( .CI(n9681), .A(n5306), .B(n5626), .S(n9705), .CO(n9706) );
  FA1A U8062 ( .CI(n5690), .A(n5370), .B(n5754), .S(n9707), .CO(n9708) );
  FA1A U8063 ( .CI(n5498), .A(n5562), .B(n5434), .S(n9709), .CO(n9710) );
  FA1A U8064 ( .CI(n9709), .A(n9687), .B(n9703), .S(n9711), .CO(n9712) );
  FA1A U8065 ( .CI(n9707), .A(n9705), .B(n9683), .S(n9713), .CO(n9714) );
  FA1A U8066 ( .CI(n9711), .A(n9689), .B(n9685), .S(n9715), .CO(n9716) );
  FA1A U8067 ( .CI(n9715), .A(n9713), .B(n9691), .S(n9717), .CO(n9718) );
  FA1A U8068 ( .CI(n9697), .A(n9695), .B(n9693), .S(n9719), .CO(n9720) );
  FA1A U8069 ( .CI(n9699), .A(n9719), .B(n9717), .S(n9721), .CO(n9722) );
  FA1A U8070 ( .CI(n5179), .A(n5819), .B(n5818), .S(n9723), .CO(n9724) );
  FA1A U8071 ( .CI(n9723), .A(n5243), .B(n5563), .S(n9725), .CO(n9726) );
  FA1A U8072 ( .CI(n5691), .A(n5755), .B(n5307), .S(n9727), .CO(n9728) );
  FA1A U8073 ( .CI(n5499), .A(n5627), .B(n5371), .S(n9729), .CO(n9730) );
  FA1A U8074 ( .CI(n9706), .A(n9704), .B(n5435), .S(n9731), .CO(n9732) );
  FA1A U8075 ( .CI(n9725), .A(n9727), .B(n9708), .S(n9733), .CO(n9734) );
  FA1A U8076 ( .CI(n9731), .A(n9729), .B(n9710), .S(n9735), .CO(n9736) );
  FA1A U8077 ( .CI(n9735), .A(n9733), .B(n9712), .S(n9737), .CO(n9738) );
  FA1A U8078 ( .CI(n9737), .A(n9716), .B(n9714), .S(n9739), .CO(n9740) );
  FA1A U8079 ( .CI(n9720), .A(n9739), .B(n9718), .S(n9741), .CO(n9742) );
  IVP U8080 ( .A(n5820), .Z(n9743) );
  FA1A U8081 ( .CI(n5308), .A(n5244), .B(n9743), .S(n9744), .CO(n9745) );
  FA1A U8082 ( .CI(n9724), .A(n5756), .B(n5628), .S(n9746), .CO(n9747) );
  FA1A U8083 ( .CI(n5500), .A(n5564), .B(n5692), .S(n9748), .CO(n9749) );
  FA1A U8084 ( .CI(n9744), .A(n5436), .B(n5372), .S(n9750), .CO(n9751) );
  FA1A U8085 ( .CI(n9750), .A(n9748), .B(n9726), .S(n9752), .CO(n9753) );
  FA1A U8086 ( .CI(n9746), .A(n9730), .B(n9728), .S(n9754), .CO(n9755) );
  FA1A U8087 ( .CI(n9752), .A(n9754), .B(n9732), .S(n9756), .CO(n9757) );
  FA1A U8088 ( .CI(n9756), .A(n9736), .B(n9734), .S(n9758), .CO(n9759) );
  FA1A U8089 ( .CI(n9740), .A(n9758), .B(n9738), .S(n9760), .CO(n9761) );
  FA1A U8090 ( .CI(n5245), .A(n5821), .B(n5820), .S(n9762), .CO(n9763) );
  FA1A U8091 ( .CI(n9762), .A(n5757), .B(n5565), .S(n9764), .CO(n9765) );
  FA1A U8092 ( .CI(n5373), .A(n5693), .B(n5309), .S(n9766), .CO(n9767) );
  FA1A U8093 ( .CI(n5501), .A(n5629), .B(n5437), .S(n9768), .CO(n9769) );
  FA1A U8094 ( .CI(n9766), .A(n9768), .B(n9745), .S(n9770), .CO(n9771) );
  FA1A U8095 ( .CI(n9751), .A(n9764), .B(n9747), .S(n9772), .CO(n9773) );
  FA1A U8096 ( .CI(n9753), .A(n9770), .B(n9749), .S(n9774), .CO(n9775) );
  FA1A U8097 ( .CI(n9774), .A(n9772), .B(n9755), .S(n9776), .CO(n9777) );
  FA1A U8098 ( .CI(n9759), .A(n9776), .B(n9757), .S(n9778), .CO(n9779) );
  IVP U8099 ( .A(n5822), .Z(n9780) );
  FA1A U8100 ( .CI(n5374), .A(n5310), .B(n9780), .S(n9781), .CO(n9782) );
  FA1A U8101 ( .CI(n9763), .A(n5438), .B(n5694), .S(n9783), .CO(n9784) );
  FA1A U8102 ( .CI(n5630), .A(n5758), .B(n5502), .S(n9785), .CO(n9786) );
  FA1A U8103 ( .CI(n9765), .A(n9781), .B(n5566), .S(n9787), .CO(n9788) );
  FA1A U8104 ( .CI(n9785), .A(n9783), .B(n9767), .S(n9789), .CO(n9790) );
  FA1A U8105 ( .CI(n9771), .A(n9787), .B(n9769), .S(n9791), .CO(n9792) );
  FA1A U8106 ( .CI(n9791), .A(n9789), .B(n9773), .S(n9793), .CO(n9794) );
  FA1A U8107 ( .CI(n9777), .A(n9793), .B(n9775), .S(n9795), .CO(n9796) );
  FA1A U8108 ( .CI(n5311), .A(n5823), .B(n5822), .S(n9797), .CO(n9798) );
  FA1A U8109 ( .CI(n9797), .A(n5375), .B(n5631), .S(n9799), .CO(n9800) );
  FA1A U8110 ( .CI(n5695), .A(n5759), .B(n5439), .S(n9801), .CO(n9802) );
  FA1A U8111 ( .CI(n9782), .A(n5567), .B(n5503), .S(n9803), .CO(n9804) );
  FA1A U8112 ( .CI(n9801), .A(n9799), .B(n9784), .S(n9805), .CO(n9806) );
  FA1A U8113 ( .CI(n9788), .A(n9803), .B(n9786), .S(n9807), .CO(n9808) );
  FA1A U8114 ( .CI(n9807), .A(n9805), .B(n9790), .S(n9809), .CO(n9810) );
  FA1A U8115 ( .CI(n9794), .A(n9809), .B(n9792), .S(n9811), .CO(n9812) );
  IVP U8116 ( .A(n5824), .Z(n9813) );
  FA1A U8117 ( .CI(n5440), .A(n5376), .B(n9813), .S(n9814), .CO(n9815) );
  FA1A U8118 ( .CI(n9798), .A(n5760), .B(n5696), .S(n9816), .CO(n9817) );
  FA1A U8119 ( .CI(n5568), .A(n5632), .B(n5504), .S(n9818), .CO(n9819) );
  FA1A U8120 ( .CI(n9816), .A(n9802), .B(n9814), .S(n9820), .CO(n9821) );
  FA1A U8121 ( .CI(n9804), .A(n9818), .B(n9800), .S(n9822), .CO(n9823) );
  FA1A U8122 ( .CI(n9822), .A(n9806), .B(n9820), .S(n9824), .CO(n9825) );
  FA1A U8123 ( .CI(n9810), .A(n9824), .B(n9808), .S(n9826), .CO(n9827) );
  FA1A U8124 ( .CI(n5377), .A(n5825), .B(n5824), .S(n9828), .CO(n9829) );
  FA1A U8125 ( .CI(n9828), .A(n5441), .B(n5633), .S(n9830), .CO(n9831) );
  FA1A U8126 ( .CI(n5569), .A(n5761), .B(n5505), .S(n9832), .CO(n9833) );
  FA1A U8127 ( .CI(n9817), .A(n9815), .B(n5697), .S(n9834), .CO(n9835) );
  FA1A U8128 ( .CI(n9832), .A(n9830), .B(n9819), .S(n9836), .CO(n9837) );
  FA1A U8129 ( .CI(n9836), .A(n9821), .B(n9834), .S(n9838), .CO(n9839) );
  FA1A U8130 ( .CI(n9825), .A(n9838), .B(n9823), .S(n9840), .CO(n9841) );
  IVP U8131 ( .A(n5826), .Z(n9842) );
  FA1A U8132 ( .CI(n5506), .A(n5442), .B(n9842), .S(n9843), .CO(n9844) );
  FA1A U8133 ( .CI(n9829), .A(n5570), .B(n5698), .S(n9845), .CO(n9846) );
  FA1A U8134 ( .CI(n9843), .A(n5762), .B(n5634), .S(n9847), .CO(n9848) );
  FA1A U8135 ( .CI(n9847), .A(n9845), .B(n9831), .S(n9849), .CO(n9850) );
  FA1A U8136 ( .CI(n9837), .A(n9835), .B(n9833), .S(n9851), .CO(n9852) );
  FA1A U8137 ( .CI(n9839), .A(n9851), .B(n9849), .S(n9853), .CO(n9854) );
  FA1A U8138 ( .CI(n5443), .A(n5827), .B(n5826), .S(n9855), .CO(n9856) );
  FA1A U8139 ( .CI(n9855), .A(n5507), .B(n5699), .S(n9857), .CO(n9858) );
  FA1A U8140 ( .CI(n5571), .A(n5635), .B(n5763), .S(n9859), .CO(n9860) );
  FA1A U8141 ( .CI(n9857), .A(n9859), .B(n9844), .S(n9861), .CO(n9862) );
  FA1A U8142 ( .CI(n9861), .A(n9848), .B(n9846), .S(n9863), .CO(n9864) );
  FA1A U8143 ( .CI(n9852), .A(n9863), .B(n9850), .S(n9865), .CO(n9866) );
  IVP U8144 ( .A(n5828), .Z(n9867) );
  FA1A U8145 ( .CI(n5572), .A(n5508), .B(n9867), .S(n9868), .CO(n9869) );
  FA1A U8146 ( .CI(n9856), .A(n5636), .B(n5764), .S(n9870), .CO(n9871) );
  FA1A U8147 ( .CI(n9858), .A(n9868), .B(n5700), .S(n9872), .CO(n9873) );
  FA1A U8148 ( .CI(n9872), .A(n9870), .B(n9860), .S(n9874), .CO(n9875) );
  FA1A U8149 ( .CI(n9864), .A(n9874), .B(n9862), .S(n9876), .CO(n9877) );
  FA1A U8150 ( .CI(n5509), .A(n5829), .B(n5828), .S(n9878), .CO(n9879) );
  FA1A U8151 ( .CI(n9878), .A(n5573), .B(n5701), .S(n9880), .CO(n9881) );
  FA1A U8152 ( .CI(n9869), .A(n5765), .B(n5637), .S(n9882), .CO(n9883) );
  FA1A U8153 ( .CI(n9882), .A(n9880), .B(n9871), .S(n9884), .CO(n9885) );
  FA1A U8154 ( .CI(n9875), .A(n9884), .B(n9873), .S(n9886), .CO(n9887) );
  IVP U8155 ( .A(n5830), .Z(n9888) );
  FA1A U8156 ( .CI(n5638), .A(n5574), .B(n9888), .S(n9889), .CO(n9890) );
  FA1A U8157 ( .CI(n9879), .A(n5766), .B(n5702), .S(n9891), .CO(n9892) );
  FA1A U8158 ( .CI(n9891), .A(n9881), .B(n9889), .S(n9893), .CO(n9894) );
  FA1A U8159 ( .CI(n9885), .A(n9893), .B(n9883), .S(n9895), .CO(n9896) );
  FA1A U8160 ( .CI(n5575), .A(n5831), .B(n5830), .S(n9897), .CO(n9898) );
  FA1A U8161 ( .CI(n9897), .A(n5703), .B(n5767), .S(n9899), .CO(n9900) );
  FA1A U8162 ( .CI(n9892), .A(n9890), .B(n5639), .S(n9901), .CO(n9902) );
  FA1A U8163 ( .CI(n9894), .A(n9901), .B(n9899), .S(n9903), .CO(n9904) );
  IVP U8164 ( .A(n5832), .Z(n9905) );
  FA1A U8165 ( .CI(n5704), .A(n5640), .B(n9905), .S(n9906), .CO(n9907) );
  FA1A U8166 ( .CI(n9906), .A(n9898), .B(n5768), .S(n9908), .CO(n9909) );
  FA1A U8167 ( .CI(n9902), .A(n9908), .B(n9900), .S(n9910), .CO(n9911) );
  FA1A U8168 ( .CI(n5641), .A(n5833), .B(n5832), .S(n9912), .CO(n9913) );
  FA1A U8169 ( .CI(n9912), .A(n5769), .B(n5705), .S(n9914), .CO(n9915) );
  FA1A U8170 ( .CI(n9909), .A(n9914), .B(n9907), .S(n9916), .CO(n9917) );
  IVP U8171 ( .A(n5834), .Z(n9918) );
  FA1A U8172 ( .CI(n5770), .A(n5706), .B(n9918), .S(n9919), .CO(n9920) );
  FA1A U8173 ( .CI(n9915), .A(n9919), .B(n9913), .S(n9921), .CO(n9922) );
  FA1A U8174 ( .CI(n5707), .A(n5835), .B(n5834), .S(n9923), .CO(n9924) );
  FA1A U8175 ( .CI(n9920), .A(n9923), .B(n5771), .S(n9925), .CO(n9926) );
  IVP U8176 ( .A(n5836), .Z(n9927) );
  FA1A U8177 ( .CI(n9924), .A(n5772), .B(n9927), .S(n9928), .CO(n9929) );
  EO3 U8178 ( .A(n5773), .B(n5836), .C(n5837), .Z(n9930) );
  HA1 U8179 ( .A(n3663), .B(n5838), .S(product[1]), .CO(n9931) );
  FA1A U8180 ( .CI(n9931), .A(n3664), .B(n10866), .S(product[2]), .CO(n9932)
         );
  FA1A U8181 ( .CI(n9932), .A(n5870), .B(n5839), .S(product[3]), .CO(n9933) );
  FA1A U8182 ( .CI(n9933), .A(n5872), .B(n5871), .S(product[4]), .CO(n9934) );
  FA1A U8183 ( .CI(n9934), .A(n5876), .B(n5873), .S(product[5]), .CO(n9935) );
  FA1A U8184 ( .CI(n9935), .A(n5880), .B(n5877), .S(product[6]), .CO(n9936) );
  FA1A U8185 ( .CI(n9936), .A(n5886), .B(n5881), .S(product[7]), .CO(n9937) );
  FA1A U8186 ( .CI(n9937), .A(n5892), .B(n5887), .S(product[8]), .CO(n9938) );
  FA1A U8187 ( .CI(n9938), .A(n5900), .B(n5893), .S(product[9]), .CO(n9939) );
  FA1A U8188 ( .CI(n9939), .A(n5908), .B(n5901), .S(product[10]), .CO(n9940)
         );
  FA1A U8189 ( .CI(n9940), .A(n5918), .B(n5909), .S(product[11]), .CO(n9941)
         );
  FA1A U8190 ( .CI(n9941), .A(n5928), .B(n5919), .S(product[12]), .CO(n9942)
         );
  FA1A U8191 ( .CI(n9942), .A(n5929), .B(n5940), .S(product[13]), .CO(n9943)
         );
  FA1A U8192 ( .CI(n9943), .A(n5952), .B(n5941), .S(product[14]), .CO(n9944)
         );
  FA1A U8193 ( .CI(n9944), .A(n5966), .B(n5953), .S(product[15]), .CO(n9945)
         );
  FA1A U8194 ( .CI(n9945), .A(n5980), .B(n5967), .S(product[16]), .CO(n9946)
         );
  FA1A U8195 ( .CI(n9946), .A(n5996), .B(n5981), .S(product[17]), .CO(n9947)
         );
  FA1A U8196 ( .CI(n9947), .A(n6012), .B(n5997), .S(product[18]), .CO(n9948)
         );
  FA1A U8197 ( .CI(n9948), .A(n6013), .B(n6030), .S(product[19]), .CO(n9949)
         );
  FA1A U8198 ( .CI(n9949), .A(n6031), .B(n6048), .S(product[20]), .CO(n9950)
         );
  FA1A U8199 ( .CI(n9950), .A(n6049), .B(n6068), .S(product[21]), .CO(n9951)
         );
  FA1A U8200 ( .CI(n9951), .A(n6088), .B(n6069), .S(product[22]), .CO(n9952)
         );
  FA1A U8201 ( .CI(n9952), .A(n6089), .B(n6110), .S(product[23]), .CO(n9953)
         );
  FA1A U8202 ( .CI(n9953), .A(n6132), .B(n6111), .S(product[24]), .CO(n9954)
         );
  FA1A U8203 ( .CI(n9954), .A(n6133), .B(n6156), .S(product[25]), .CO(n9955)
         );
  FA1A U8204 ( .CI(n9955), .A(n6180), .B(n6157), .S(product[26]), .CO(n9956)
         );
  FA1A U8205 ( .CI(n9956), .A(n6206), .B(n6181), .S(product[27]), .CO(n9957)
         );
  FA1A U8206 ( .CI(n9957), .A(n6232), .B(n6207), .S(product[28]), .CO(n9958)
         );
  FA1A U8207 ( .CI(n9958), .A(n6233), .B(n6260), .S(product[29]), .CO(n9959)
         );
  FA1A U8208 ( .CI(n9959), .A(n6261), .B(n6288), .S(product[30]), .CO(n9960)
         );
  FA1A U8209 ( .CI(n9960), .A(n6318), .B(n6289), .S(product[31]), .CO(n9961)
         );
  FA1A U8210 ( .CI(n9961), .A(n6348), .B(n6319), .S(product[32]), .CO(n9962)
         );
  FA1A U8211 ( .CI(n9962), .A(n6380), .B(n6349), .S(product[33]), .CO(n9963)
         );
  FA1A U8212 ( .CI(n9963), .A(n6381), .B(n6412), .S(product[34]), .CO(n9964)
         );
  FA1A U8213 ( .CI(n9964), .A(n6413), .B(n6446), .S(product[35]), .CO(n9965)
         );
  FA1A U8214 ( .CI(n9965), .A(n6447), .B(n6480), .S(product[36]), .CO(n9966)
         );
  FA1A U8215 ( .CI(n9966), .A(n6516), .B(n6481), .S(product[37]), .CO(n9967)
         );
  FA1A U8216 ( .CI(n9967), .A(n6517), .B(n6552), .S(product[38]), .CO(n9968)
         );
  FA1A U8217 ( .CI(n9968), .A(n6590), .B(n6553), .S(product[39]), .CO(n9969)
         );
  FA1A U8218 ( .CI(n9969), .A(n6628), .B(n6591), .S(product[40]), .CO(n9970)
         );
  FA1A U8219 ( .CI(n9970), .A(n6668), .B(n6629), .S(product[41]), .CO(n9971)
         );
  FA1A U8220 ( .CI(n9971), .A(n6708), .B(n6669), .S(product[42]), .CO(n9972)
         );
  FA1A U8221 ( .CI(n9972), .A(n6709), .B(n6750), .S(product[43]), .CO(n9973)
         );
  FA1A U8222 ( .CI(n9973), .A(n6751), .B(n6792), .S(product[44]), .CO(n9974)
         );
  FA1A U8223 ( .CI(n9974), .A(n6793), .B(n6836), .S(product[45]), .CO(n9975)
         );
  FA1A U8224 ( .CI(n9975), .A(n6837), .B(n6880), .S(product[46]), .CO(n9976)
         );
  FA1A U8225 ( .CI(n9976), .A(n6926), .B(n6881), .S(product[47]), .CO(n9977)
         );
  FA1A U8226 ( .CI(n9977), .A(n6972), .B(n6927), .S(product[48]), .CO(n9978)
         );
  FA1A U8227 ( .CI(n9978), .A(n6973), .B(n7020), .S(product[49]), .CO(n9979)
         );
  FA1A U8228 ( .CI(n9979), .A(n7021), .B(n7068), .S(product[50]), .CO(n9980)
         );
  FA1A U8229 ( .CI(n9980), .A(n7069), .B(n7118), .S(product[51]), .CO(n9981)
         );
  FA1A U8230 ( .CI(n9981), .A(n7119), .B(n7168), .S(product[52]), .CO(n9982)
         );
  FA1A U8231 ( .CI(n9982), .A(n7169), .B(n7220), .S(product[53]), .CO(n9983)
         );
  FA1A U8232 ( .CI(n9983), .A(n7221), .B(n7272), .S(product[54]), .CO(n9984)
         );
  FA1A U8233 ( .CI(n9984), .A(n7273), .B(n7326), .S(product[55]), .CO(n9985)
         );
  FA1A U8234 ( .CI(n9985), .A(n7327), .B(n7380), .S(product[56]), .CO(n9986)
         );
  FA1A U8235 ( .CI(n9986), .A(n7381), .B(n7436), .S(product[57]), .CO(n9987)
         );
  FA1A U8236 ( .CI(n9987), .A(n7492), .B(n7437), .S(product[58]), .CO(n9988)
         );
  FA1A U8237 ( .CI(n9988), .A(n7550), .B(n7493), .S(product[59]), .CO(n9989)
         );
  FA1A U8238 ( .CI(n9989), .A(n7608), .B(n7551), .S(product[60]), .CO(n9990)
         );
  FA1A U8239 ( .CI(n9990), .A(n7609), .B(n7668), .S(product[61]), .CO(n9991)
         );
  FA1A U8240 ( .CI(n9991), .A(n7669), .B(n7728), .S(product[62]), .CO(n9992)
         );
  FA1A U8241 ( .CI(n9992), .A(n7790), .B(n7729), .S(product[63]), .CO(n9993)
         );
  FA1A U8242 ( .CI(n9993), .A(n7791), .B(n7852), .S(product[64]), .CO(n9994)
         );
  FA1A U8243 ( .CI(n9994), .A(n7853), .B(n7915), .S(product[65]), .CO(n9995)
         );
  FA1A U8244 ( .CI(n9995), .A(n7916), .B(n7978), .S(product[66]), .CO(n9996)
         );
  FA1A U8245 ( .CI(n9996), .A(n7979), .B(n8040), .S(product[67]), .CO(n9997)
         );
  FA1A U8246 ( .CI(n9997), .A(n8041), .B(n8101), .S(product[68]), .CO(n9998)
         );
  FA1A U8247 ( .CI(n9998), .A(n8102), .B(n8161), .S(product[69]), .CO(n9999)
         );
  FA1A U8248 ( .CI(n9999), .A(n8162), .B(n8220), .S(product[70]), .CO(n10000)
         );
  FA1A U8249 ( .CI(n10000), .A(n8221), .B(n8278), .S(product[71]), .CO(n10001)
         );
  FA1A U8250 ( .CI(n10001), .A(n8279), .B(n8335), .S(product[72]), .CO(n10002)
         );
  FA1A U8251 ( .CI(n10002), .A(n8336), .B(n8391), .S(product[73]), .CO(n10003)
         );
  FA1A U8252 ( .CI(n10003), .A(n8392), .B(n8446), .S(product[74]), .CO(n10004)
         );
  FA1A U8253 ( .CI(n10004), .A(n8447), .B(n8500), .S(product[75]), .CO(n10005)
         );
  FA1A U8254 ( .CI(n10005), .A(n8501), .B(n8553), .S(product[76]), .CO(n10006)
         );
  FA1A U8255 ( .CI(n10006), .A(n8554), .B(n8605), .S(product[77]), .CO(n10007)
         );
  FA1A U8256 ( .CI(n10007), .A(n8606), .B(n8656), .S(product[78]), .CO(n10008)
         );
  FA1A U8257 ( .CI(n10008), .A(n8657), .B(n8706), .S(product[79]), .CO(n10009)
         );
  FA1A U8258 ( .CI(n10009), .A(n8707), .B(n8755), .S(product[80]), .CO(n10010)
         );
  FA1A U8259 ( .CI(n10010), .A(n8756), .B(n8803), .S(product[81]), .CO(n10011)
         );
  FA1A U8260 ( .CI(n10011), .A(n8804), .B(n8850), .S(product[82]), .CO(n10012)
         );
  FA1A U8261 ( .CI(n10012), .A(n8851), .B(n8896), .S(product[83]), .CO(n10013)
         );
  FA1A U8262 ( .CI(n10013), .A(n8897), .B(n8941), .S(product[84]), .CO(n10014)
         );
  FA1A U8263 ( .CI(n10014), .A(n8942), .B(n8985), .S(product[85]), .CO(n10015)
         );
  FA1A U8264 ( .CI(n10015), .A(n8986), .B(n9028), .S(product[86]), .CO(n10016)
         );
  FA1A U8265 ( .CI(n10016), .A(n9029), .B(n9070), .S(product[87]), .CO(n10017)
         );
  FA1A U8266 ( .CI(n10017), .A(n9071), .B(n9111), .S(product[88]), .CO(n10018)
         );
  FA1A U8267 ( .CI(n10018), .A(n9112), .B(n9151), .S(product[89]), .CO(n10019)
         );
  FA1A U8268 ( .CI(n10019), .A(n9152), .B(n9190), .S(product[90]), .CO(n10020)
         );
  FA1A U8269 ( .CI(n10020), .A(n9191), .B(n9228), .S(product[91]), .CO(n10021)
         );
  FA1A U8270 ( .CI(n10021), .A(n9229), .B(n9265), .S(product[92]), .CO(n10022)
         );
  FA1A U8271 ( .CI(n10022), .A(n9266), .B(n9301), .S(product[93]), .CO(n10023)
         );
  FA1A U8272 ( .CI(n10023), .A(n9302), .B(n9336), .S(product[94]), .CO(n10024)
         );
  FA1A U8273 ( .CI(n10024), .A(n9337), .B(n9370), .S(product[95]), .CO(n10025)
         );
  FA1A U8274 ( .CI(n10025), .A(n9371), .B(n9403), .S(product[96]), .CO(n10026)
         );
  FA1A U8275 ( .CI(n10026), .A(n9404), .B(n9435), .S(product[97]), .CO(n10027)
         );
  FA1A U8276 ( .CI(n10027), .A(n9436), .B(n9466), .S(product[98]), .CO(n10028)
         );
  FA1A U8277 ( .CI(n10028), .A(n9467), .B(n9496), .S(product[99]), .CO(n10029)
         );
  FA1A U8278 ( .CI(n10029), .A(n9497), .B(n9525), .S(product[100]), .CO(n10030) );
  FA1A U8279 ( .CI(n10030), .A(n9526), .B(n9553), .S(product[101]), .CO(n10031) );
  FA1A U8280 ( .CI(n10031), .A(n9554), .B(n9580), .S(product[102]), .CO(n10032) );
  FA1A U8281 ( .CI(n10032), .A(n9581), .B(n9606), .S(product[103]), .CO(n10033) );
  FA1A U8282 ( .CI(n10033), .A(n9607), .B(n9631), .S(product[104]), .CO(n10034) );
  FA1A U8283 ( .CI(n10034), .A(n9632), .B(n9655), .S(product[105]), .CO(n10035) );
  FA1A U8284 ( .CI(n10035), .A(n9656), .B(n9678), .S(product[106]), .CO(n10036) );
  FA1A U8285 ( .CI(n10036), .A(n9679), .B(n9700), .S(product[107]), .CO(n10037) );
  FA1A U8286 ( .CI(n10037), .A(n9701), .B(n9721), .S(product[108]), .CO(n10038) );
  FA1A U8287 ( .CI(n10038), .A(n9722), .B(n9741), .S(product[109]), .CO(n10039) );
  FA1A U8288 ( .CI(n10039), .A(n9742), .B(n9760), .S(product[110]), .CO(n10040) );
  FA1A U8289 ( .CI(n10040), .A(n9761), .B(n9778), .S(product[111]), .CO(n10041) );
  FA1A U8290 ( .CI(n10041), .A(n9779), .B(n9795), .S(product[112]), .CO(n10042) );
  FA1A U8291 ( .CI(n10042), .A(n9796), .B(n9811), .S(product[113]), .CO(n10043) );
  FA1A U8292 ( .CI(n10043), .A(n9812), .B(n9826), .S(product[114]), .CO(n10044) );
  FA1A U8293 ( .CI(n10044), .A(n9827), .B(n9840), .S(product[115]), .CO(n10045) );
  FA1A U8294 ( .CI(n10045), .A(n9841), .B(n9853), .S(product[116]), .CO(n10046) );
  FA1A U8295 ( .CI(n10046), .A(n9854), .B(n9865), .S(product[117]), .CO(n10047) );
  FA1A U8296 ( .CI(n10047), .A(n9866), .B(n9876), .S(product[118]), .CO(n10048) );
  FA1A U8297 ( .CI(n10048), .A(n9877), .B(n9886), .S(product[119]), .CO(n10049) );
  FA1A U8298 ( .CI(n10049), .A(n9887), .B(n9895), .S(product[120]), .CO(n10050) );
  FA1A U8299 ( .CI(n10050), .A(n9896), .B(n9903), .S(product[121]), .CO(n10051) );
  FA1A U8300 ( .CI(n10051), .A(n9904), .B(n9910), .S(product[122]), .CO(n10052) );
  FA1A U8301 ( .CI(n10052), .A(n9911), .B(n9916), .S(product[123]), .CO(n10053) );
  FA1A U8302 ( .CI(n10053), .A(n9917), .B(n9921), .S(product[124]), .CO(n10054) );
  FA1A U8303 ( .CI(n10054), .A(n9922), .B(n9925), .S(product[125]), .CO(n10055) );
  FA1A U8304 ( .CI(n10055), .A(n9926), .B(n9928), .S(product[126]), .CO(n10056) );
  EO U8305 ( .A(n9929), .B(n9930), .Z(n10057) );
  EO U8306 ( .A(n10056), .B(n10057), .Z(product[127]) );
  AN2P U8307 ( .A(n10251), .B(n1060), .Z(n10866) );
  AN2P U8308 ( .A(n10247), .B(n875), .Z(n10867) );
  AN2P U8309 ( .A(n10247), .B(n880), .Z(n10868) );
  AN2P U8310 ( .A(n10247), .B(n886), .Z(n10869) );
  AN2P U8311 ( .A(n10247), .B(n892), .Z(n10870) );
  AN2P U8312 ( .A(n10247), .B(n898), .Z(n10871) );
  AN2P U8313 ( .A(n10247), .B(n904), .Z(n10872) );
  AN2P U8314 ( .A(n10247), .B(n910), .Z(n10873) );
  AN2P U8315 ( .A(n10247), .B(n916), .Z(n10874) );
  AN2P U8316 ( .A(n10248), .B(n922), .Z(n10875) );
  AN2P U8317 ( .A(n10248), .B(n928), .Z(n10876) );
  AN2P U8318 ( .A(n10248), .B(n934), .Z(n10877) );
  AN2P U8319 ( .A(n10248), .B(n940), .Z(n10878) );
  AN2P U8320 ( .A(n10248), .B(n946), .Z(n10879) );
  AN2P U8321 ( .A(n10248), .B(n952), .Z(n10880) );
  AN2P U8322 ( .A(n10248), .B(n958), .Z(n10881) );
  AN2P U8323 ( .A(n10249), .B(n964), .Z(n10882) );
  AN2P U8324 ( .A(n10249), .B(n970), .Z(n10883) );
  AN2P U8325 ( .A(n10249), .B(n976), .Z(n10884) );
  AN2P U8326 ( .A(n10249), .B(n982), .Z(n10885) );
  AN2P U8327 ( .A(n10249), .B(n988), .Z(n10886) );
  AN2P U8328 ( .A(n10249), .B(n994), .Z(n10887) );
  AN2P U8329 ( .A(n10249), .B(n1000), .Z(n10888) );
  AN2P U8330 ( .A(n10250), .B(n1006), .Z(n10889) );
  AN2P U8331 ( .A(n10250), .B(n1012), .Z(n10890) );
  AN2P U8332 ( .A(n10250), .B(n1018), .Z(n10891) );
  AN2P U8333 ( .A(n10250), .B(n1024), .Z(n10892) );
  AN2P U8334 ( .A(n10250), .B(n1030), .Z(n10893) );
  AN2P U8335 ( .A(n10250), .B(n1036), .Z(n10894) );
  AN2P U8336 ( .A(n10250), .B(n1042), .Z(n10895) );
  AN2P U8337 ( .A(n10251), .B(n1048), .Z(n10896) );
  AN2P U8338 ( .A(n10251), .B(n1054), .Z(n10897) );
  AN2P U8339 ( .A(n10251), .B(n1066), .Z(product[0]) );
  IVP U8340 ( .A(n243), .Z(n10535) );
  IVP U8341 ( .A(n253), .Z(n10525) );
  IVP U8342 ( .A(n248), .Z(n10530) );
  IVP U8343 ( .A(n214), .Z(n10564) );
  IVP U8344 ( .A(n282), .Z(n10496) );
  IVP U8345 ( .A(n219), .Z(n10559) );
  IVP U8346 ( .A(n263), .Z(n10515) );
  IVP U8347 ( .A(n287), .Z(n10491) );
  IVP U8348 ( .A(n258), .Z(n10520) );
  IVP U8349 ( .A(n268), .Z(n10510) );
  IVP U8350 ( .A(n224), .Z(n10554) );
  IVP U8351 ( .A(n292), .Z(n10486) );
  IVP U8352 ( .A(n302), .Z(n10476) );
  IVP U8353 ( .A(n273), .Z(n10505) );
  IVP U8354 ( .A(n234), .Z(n10544) );
  IVP U8355 ( .A(n229), .Z(n10549) );
  IVP U8356 ( .A(n297), .Z(n10481) );
  IVP U8357 ( .A(n239), .Z(n10539) );
  IVP U8358 ( .A(n307), .Z(n10471) );
  IVP U8359 ( .A(n244), .Z(n10534) );
  IVP U8360 ( .A(n312), .Z(n10466) );
  IVP U8361 ( .A(n278), .Z(n10500) );
  IVP U8362 ( .A(n283), .Z(n10495) );
  IVP U8363 ( .A(n249), .Z(n10529) );
  IVP U8364 ( .A(n317), .Z(n10461) );
  IVP U8365 ( .A(n254), .Z(n10524) );
  IVP U8366 ( .A(n322), .Z(n10456) );
  IVP U8367 ( .A(n288), .Z(n10490) );
  IVP U8368 ( .A(n293), .Z(n10485) );
  IVP U8369 ( .A(n327), .Z(n10451) );
  IVP U8370 ( .A(n308), .Z(n10470) );
  IVP U8371 ( .A(n259), .Z(n10519) );
  IVP U8372 ( .A(n274), .Z(n10504) );
  IVP U8373 ( .A(n264), .Z(n10514) );
  IVP U8374 ( .A(n342), .Z(n10436) );
  IVP U8375 ( .A(n332), .Z(n10446) );
  IVP U8376 ( .A(n269), .Z(n10509) );
  IVP U8377 ( .A(n337), .Z(n10441) );
  IVP U8378 ( .A(n298), .Z(n10480) );
  IVP U8379 ( .A(n303), .Z(n10475) );
  IVP U8380 ( .A(n313), .Z(n10465) );
  IVP U8381 ( .A(n279), .Z(n10499) );
  IVP U8382 ( .A(n347), .Z(n10431) );
  IVP U8383 ( .A(n352), .Z(n10426) );
  IVP U8384 ( .A(n318), .Z(n10460) );
  IVP U8385 ( .A(n284), .Z(n10494) );
  IVP U8386 ( .A(n289), .Z(n10489) );
  IVP U8387 ( .A(n250), .Z(n10528) );
  IVP U8388 ( .A(n255), .Z(n10523) );
  IVP U8389 ( .A(n260), .Z(n10518) );
  IVP U8390 ( .A(n238), .Z(n10540) );
  IVP U8391 ( .A(n228), .Z(n10550) );
  IVP U8392 ( .A(n233), .Z(n10545) );
  IVP U8393 ( .A(n252), .Z(n10526) );
  IVP U8394 ( .A(n262), .Z(n10516) );
  IVP U8395 ( .A(n267), .Z(n10511) );
  IVP U8396 ( .A(n223), .Z(n10555) );
  IVP U8397 ( .A(n277), .Z(n10501) );
  IVP U8398 ( .A(n257), .Z(n10521) );
  IVP U8399 ( .A(n218), .Z(n10560) );
  IVP U8400 ( .A(n272), .Z(n10506) );
  IVP U8401 ( .A(n213), .Z(n10565) );
  IVP U8402 ( .A(n209), .Z(n10569) );
  IVP U8403 ( .A(n204), .Z(n10574) );
  IVP U8404 ( .A(n323), .Z(n10455) );
  IVP U8405 ( .A(n357), .Z(n10421) );
  IVP U8406 ( .A(n265), .Z(n10513) );
  IVP U8407 ( .A(n294), .Z(n10484) );
  IVP U8408 ( .A(n275), .Z(n10503) );
  IVP U8409 ( .A(n270), .Z(n10508) );
  IVP U8410 ( .A(n328), .Z(n10450) );
  IVP U8411 ( .A(n333), .Z(n10445) );
  IVP U8412 ( .A(n299), .Z(n10479) );
  IVP U8413 ( .A(n280), .Z(n10498) );
  IVP U8414 ( .A(n304), .Z(n10474) );
  IVP U8415 ( .A(n338), .Z(n10440) );
  IVP U8416 ( .A(n314), .Z(n10464) );
  IVP U8417 ( .A(n343), .Z(n10435) );
  IVP U8418 ( .A(n290), .Z(n10488) );
  IVP U8419 ( .A(n348), .Z(n10430) );
  IVP U8420 ( .A(n309), .Z(n10469) );
  IVP U8421 ( .A(n285), .Z(n10493) );
  IVP U8422 ( .A(n319), .Z(n10459) );
  IVP U8423 ( .A(n353), .Z(n10425) );
  IVP U8424 ( .A(n295), .Z(n10483) );
  IVP U8425 ( .A(n324), .Z(n10454) );
  IVP U8426 ( .A(n300), .Z(n10478) );
  IVP U8427 ( .A(n240), .Z(n10538) );
  IVP U8428 ( .A(n245), .Z(n10533) );
  IVP U8429 ( .A(n212), .Z(n10566) );
  IVP U8430 ( .A(n237), .Z(n10541) );
  IVP U8431 ( .A(n242), .Z(n10536) );
  IVP U8432 ( .A(n227), .Z(n10551) );
  IVP U8433 ( .A(n222), .Z(n10556) );
  IVP U8434 ( .A(n208), .Z(n10570) );
  IVP U8435 ( .A(n232), .Z(n10546) );
  IVP U8436 ( .A(n203), .Z(n10575) );
  IVP U8437 ( .A(n247), .Z(n10531) );
  IVP U8438 ( .A(n358), .Z(n10420) );
  IVP U8439 ( .A(n329), .Z(n10449) );
  IVP U8440 ( .A(n305), .Z(n10473) );
  IVP U8441 ( .A(n320), .Z(n10458) );
  IVP U8442 ( .A(n334), .Z(n10444) );
  IVP U8443 ( .A(n339), .Z(n10439) );
  IVP U8444 ( .A(n315), .Z(n10463) );
  IVP U8445 ( .A(n310), .Z(n10468) );
  IVP U8446 ( .A(n344), .Z(n10434) );
  IVP U8447 ( .A(n349), .Z(n10429) );
  IVP U8448 ( .A(n325), .Z(n10453) );
  IVP U8449 ( .A(n230), .Z(n10548) );
  IVP U8450 ( .A(n235), .Z(n10543) );
  IVP U8451 ( .A(n207), .Z(n10571) );
  IVP U8452 ( .A(n217), .Z(n10561) );
  IVP U8453 ( .A(n354), .Z(n10424) );
  IVP U8454 ( .A(n359), .Z(n10419) );
  IVP U8455 ( .A(n330), .Z(n10448) );
  IVP U8456 ( .A(n335), .Z(n10443) );
  IVP U8457 ( .A(n340), .Z(n10438) );
  IVP U8458 ( .A(n220), .Z(n10558) );
  IVP U8459 ( .A(n225), .Z(n10553) );
  IVP U8460 ( .A(n202), .Z(n10576) );
  IVP U8461 ( .A(n345), .Z(n10433) );
  IVP U8462 ( .A(n350), .Z(n10428) );
  IVP U8463 ( .A(n210), .Z(n10568) );
  IVP U8464 ( .A(n215), .Z(n10563) );
  IVP U8465 ( .A(n360), .Z(n10418) );
  IVP U8466 ( .A(n355), .Z(n10423) );
  IVP U8467 ( .A(n205), .Z(n10573) );
  IVP U8468 ( .A(n301), .Z(n10477) );
  IVP U8469 ( .A(n306), .Z(n10472) );
  IVP U8470 ( .A(n311), .Z(n10467) );
  IVP U8471 ( .A(n316), .Z(n10462) );
  IVP U8472 ( .A(n321), .Z(n10457) );
  IVP U8473 ( .A(n326), .Z(n10452) );
  IVP U8474 ( .A(n331), .Z(n10447) );
  IVP U8475 ( .A(n336), .Z(n10442) );
  IVP U8476 ( .A(n341), .Z(n10437) );
  IVP U8477 ( .A(n346), .Z(n10432) );
  IVP U8478 ( .A(n351), .Z(n10427) );
  IVP U8479 ( .A(n356), .Z(n10422) );
  IVP U8480 ( .A(n266), .Z(n10512) );
  IVP U8481 ( .A(n271), .Z(n10507) );
  IVP U8482 ( .A(n276), .Z(n10502) );
  IVP U8483 ( .A(n296), .Z(n10482) );
  IVP U8484 ( .A(n291), .Z(n10487) );
  IVP U8485 ( .A(n281), .Z(n10497) );
  IVP U8486 ( .A(n286), .Z(n10492) );
  IVP U8487 ( .A(n246), .Z(n10532) );
  IVP U8488 ( .A(n261), .Z(n10517) );
  IVP U8489 ( .A(n251), .Z(n10527) );
  IVP U8490 ( .A(n256), .Z(n10522) );
  IVP U8491 ( .A(n226), .Z(n10552) );
  IVP U8492 ( .A(n231), .Z(n10547) );
  IVP U8493 ( .A(n236), .Z(n10542) );
  IVP U8494 ( .A(n241), .Z(n10537) );
  IVP U8495 ( .A(n216), .Z(n10562) );
  IVP U8496 ( .A(n221), .Z(n10557) );
  IVP U8497 ( .A(n211), .Z(n10567) );
  IVP U8498 ( .A(n206), .Z(n10572) );
  IVP U8499 ( .A(n201), .Z(n10577) );
  IVP U8500 ( .A(n143), .Z(n10635) );
  IVP U8501 ( .A(n60), .Z(n10700) );
  IVP U8502 ( .A(n117), .Z(n10661) );
  IVP U8503 ( .A(n88), .Z(n10690) );
  IVP U8504 ( .A(n108), .Z(n10670) );
  IVP U8505 ( .A(n103), .Z(n10675) );
  IVP U8506 ( .A(n142), .Z(n10636) );
  IVP U8507 ( .A(n147), .Z(n10631) );
  IVP U8508 ( .A(n113), .Z(n10665) );
  IVP U8509 ( .A(n70), .Z(n10699) );
  IVP U8510 ( .A(n84), .Z(n10694) );
  IVP U8511 ( .A(n157), .Z(n10621) );
  IVP U8512 ( .A(n182), .Z(n10596) );
  IVP U8513 ( .A(n114), .Z(n10664) );
  IVP U8514 ( .A(n148), .Z(n10630) );
  IVP U8515 ( .A(n119), .Z(n10659) );
  IVP U8516 ( .A(n187), .Z(n10591) );
  IVP U8517 ( .A(n153), .Z(n10625) );
  IVP U8518 ( .A(n197), .Z(n10581) );
  IVP U8519 ( .A(n31), .Z(n10711) );
  IVP U8520 ( .A(n36), .Z(n10706) );
  IVP U8521 ( .A(n92), .Z(n10686) );
  IVP U8522 ( .A(n27), .Z(n10715) );
  IVP U8523 ( .A(n97), .Z(n10681) );
  IVP U8524 ( .A(n102), .Z(n10676) );
  IVP U8525 ( .A(n32), .Z(n10710) );
  IVP U8526 ( .A(n112), .Z(n10666) );
  IVP U8527 ( .A(n107), .Z(n10671) );
  IVP U8528 ( .A(n83), .Z(n10695) );
  IVP U8529 ( .A(n37), .Z(n10705) );
  IVP U8530 ( .A(n8), .Z(n10734) );
  IVP U8531 ( .A(n13), .Z(n10729) );
  IVP U8532 ( .A(n18), .Z(n10724) );
  IVP U8533 ( .A(n122), .Z(n10656) );
  IVP U8534 ( .A(n127), .Z(n10651) );
  IVP U8535 ( .A(n93), .Z(n10685) );
  IVP U8536 ( .A(n23), .Z(n10719) );
  IVP U8537 ( .A(n28), .Z(n10714) );
  IVP U8538 ( .A(n132), .Z(n10646) );
  IVP U8539 ( .A(n98), .Z(n10680) );
  IVP U8540 ( .A(n137), .Z(n10641) );
  IVP U8541 ( .A(n33), .Z(n10709) );
  IVP U8542 ( .A(n38), .Z(n10704) );
  IVP U8543 ( .A(n152), .Z(n10626) );
  IVP U8544 ( .A(n118), .Z(n10660) );
  IVP U8545 ( .A(n94), .Z(n10684) );
  IVP U8546 ( .A(n123), .Z(n10655) );
  IVP U8547 ( .A(n89), .Z(n10689) );
  IVP U8548 ( .A(n128), .Z(n10650) );
  IVP U8549 ( .A(n162), .Z(n10616) );
  IVP U8550 ( .A(n167), .Z(n10611) );
  IVP U8551 ( .A(n133), .Z(n10645) );
  IVP U8552 ( .A(n138), .Z(n10640) );
  IVP U8553 ( .A(n99), .Z(n10679) );
  IVP U8554 ( .A(n172), .Z(n10606) );
  IVP U8555 ( .A(n104), .Z(n10674) );
  IVP U8556 ( .A(n109), .Z(n10669) );
  IVP U8557 ( .A(n177), .Z(n10601) );
  IVP U8558 ( .A(n124), .Z(n10654) );
  IVP U8559 ( .A(n158), .Z(n10620) );
  IVP U8560 ( .A(n192), .Z(n10586) );
  IVP U8561 ( .A(n129), .Z(n10649) );
  IVP U8562 ( .A(n163), .Z(n10615) );
  IVP U8563 ( .A(n134), .Z(n10644) );
  IVP U8564 ( .A(n193), .Z(n10585) );
  IVP U8565 ( .A(n159), .Z(n10619) );
  IVP U8566 ( .A(n26), .Z(n10716) );
  IVP U8567 ( .A(n50), .Z(n10701) );
  IVP U8568 ( .A(n12), .Z(n10730) );
  IVP U8569 ( .A(n3), .Z(n10735) );
  IVP U8570 ( .A(n82), .Z(n10696) );
  IVP U8571 ( .A(n87), .Z(n10691) );
  IVP U8572 ( .A(n17), .Z(n10725) );
  IVP U8573 ( .A(n22), .Z(n10720) );
  IVP U8574 ( .A(n168), .Z(n10610) );
  IVP U8575 ( .A(n144), .Z(n10634) );
  IVP U8576 ( .A(n139), .Z(n10639) );
  IVP U8577 ( .A(n173), .Z(n10605) );
  IVP U8578 ( .A(n178), .Z(n10600) );
  IVP U8579 ( .A(n183), .Z(n10595) );
  IVP U8580 ( .A(n154), .Z(n10624) );
  IVP U8581 ( .A(n149), .Z(n10629) );
  IVP U8582 ( .A(n188), .Z(n10590) );
  IVP U8583 ( .A(n164), .Z(n10614) );
  IVP U8584 ( .A(n198), .Z(n10580) );
  IVP U8585 ( .A(n169), .Z(n10609) );
  IVP U8586 ( .A(n2), .Z(n10736) );
  IVP U8587 ( .A(n11), .Z(n10731) );
  IVP U8588 ( .A(n16), .Z(n10726) );
  IVP U8589 ( .A(n21), .Z(n10721) );
  IVP U8590 ( .A(n174), .Z(n10604) );
  IVP U8591 ( .A(n179), .Z(n10599) );
  IVP U8592 ( .A(n184), .Z(n10594) );
  IVP U8593 ( .A(n189), .Z(n10589) );
  IVP U8594 ( .A(n194), .Z(n10584) );
  IVP U8595 ( .A(n199), .Z(n10579) );
  IVP U8596 ( .A(n9), .Z(n10733) );
  IVP U8597 ( .A(n90), .Z(n10688) );
  IVP U8598 ( .A(n95), .Z(n10683) );
  IVP U8599 ( .A(n100), .Z(n10678) );
  IVP U8600 ( .A(n105), .Z(n10673) );
  IVP U8601 ( .A(n115), .Z(n10663) );
  IVP U8602 ( .A(n110), .Z(n10668) );
  IVP U8603 ( .A(n120), .Z(n10658) );
  IVP U8604 ( .A(n130), .Z(n10648) );
  IVP U8605 ( .A(n125), .Z(n10653) );
  IVP U8606 ( .A(n140), .Z(n10638) );
  IVP U8607 ( .A(n135), .Z(n10643) );
  IVP U8608 ( .A(n160), .Z(n10618) );
  IVP U8609 ( .A(n80), .Z(n10698) );
  IVP U8610 ( .A(n85), .Z(n10693) );
  IVP U8611 ( .A(n145), .Z(n10633) );
  IVP U8612 ( .A(n150), .Z(n10628) );
  IVP U8613 ( .A(n155), .Z(n10623) );
  IVP U8614 ( .A(n170), .Z(n10608) );
  IVP U8615 ( .A(n165), .Z(n10613) );
  IVP U8616 ( .A(n34), .Z(n10708) );
  IVP U8617 ( .A(n39), .Z(n10703) );
  IVP U8618 ( .A(n175), .Z(n10603) );
  IVP U8619 ( .A(n185), .Z(n10593) );
  IVP U8620 ( .A(n180), .Z(n10598) );
  IVP U8621 ( .A(n24), .Z(n10718) );
  IVP U8622 ( .A(n29), .Z(n10713) );
  IVP U8623 ( .A(n19), .Z(n10723) );
  IVP U8624 ( .A(n190), .Z(n10588) );
  IVP U8625 ( .A(n195), .Z(n10583) );
  IVP U8626 ( .A(n200), .Z(n10578) );
  IVP U8627 ( .A(n14), .Z(n10728) );
  IVP U8628 ( .A(n1137), .Z(n1431) );
  IVP U8629 ( .A(n1134), .Z(n1432) );
  IVP U8630 ( .A(n1125), .Z(n1435) );
  IVP U8631 ( .A(n1119), .Z(n1437) );
  IVP U8632 ( .A(n1116), .Z(n1438) );
  IVP U8633 ( .A(n1131), .Z(n1433) );
  IVP U8634 ( .A(n1113), .Z(n1439) );
  IVP U8635 ( .A(n1122), .Z(n1436) );
  IVP U8636 ( .A(n1104), .Z(n1442) );
  IVP U8637 ( .A(n1098), .Z(n1444) );
  IVP U8638 ( .A(n1101), .Z(n1443) );
  IVP U8639 ( .A(n1095), .Z(n1445) );
  IVP U8640 ( .A(n1110), .Z(n1440) );
  IVP U8641 ( .A(n1092), .Z(n1446) );
  IVP U8642 ( .A(n1107), .Z(n1441) );
  IVP U8643 ( .A(n1143), .Z(n1429) );
  IVP U8644 ( .A(n1140), .Z(n1430) );
  IVP U8645 ( .A(n1128), .Z(n1434) );
  IVP U8646 ( .A(n1089), .Z(n1447) );
  IVP U8647 ( .A(n1086), .Z(n1448) );
  IVP U8648 ( .A(n1083), .Z(n1449) );
  IVP U8649 ( .A(n1080), .Z(n1450) );
  IVP U8650 ( .A(n1077), .Z(n1451) );
  IVP U8651 ( .A(n1149), .Z(n1427) );
  IVP U8652 ( .A(n1161), .Z(n1423) );
  IVP U8653 ( .A(n1146), .Z(n1428) );
  IVP U8654 ( .A(n1074), .Z(n1452) );
  IVP U8655 ( .A(n1071), .Z(n1453) );
  IVP U8656 ( .A(n1155), .Z(n1425) );
  IVP U8657 ( .A(n1152), .Z(n1426) );
  IVP U8658 ( .A(n1158), .Z(n1424) );
  IVP U8659 ( .A(n1164), .Z(n1422) );
  IVP U8660 ( .A(n146), .Z(n10632) );
  IVP U8661 ( .A(n181), .Z(n10597) );
  IVP U8662 ( .A(n136), .Z(n10642) );
  IVP U8663 ( .A(n141), .Z(n10637) );
  IVP U8664 ( .A(n151), .Z(n10627) );
  IVP U8665 ( .A(n156), .Z(n10622) );
  IVP U8666 ( .A(n161), .Z(n10617) );
  IVP U8667 ( .A(n166), .Z(n10612) );
  IVP U8668 ( .A(n171), .Z(n10607) );
  IVP U8669 ( .A(n186), .Z(n10592) );
  IVP U8670 ( .A(n176), .Z(n10602) );
  IVP U8671 ( .A(n191), .Z(n10587) );
  IVP U8672 ( .A(n196), .Z(n10582) );
  IVP U8673 ( .A(n131), .Z(n10647) );
  IVP U8674 ( .A(n106), .Z(n10672) );
  IVP U8675 ( .A(n101), .Z(n10677) );
  IVP U8676 ( .A(n111), .Z(n10667) );
  IVP U8677 ( .A(n116), .Z(n10662) );
  IVP U8678 ( .A(n121), .Z(n10657) );
  IVP U8679 ( .A(n126), .Z(n10652) );
  IVP U8680 ( .A(n35), .Z(n10707) );
  IVP U8681 ( .A(n40), .Z(n10702) );
  IVP U8682 ( .A(n81), .Z(n10697) );
  IVP U8683 ( .A(n86), .Z(n10692) );
  IVP U8684 ( .A(n91), .Z(n10687) );
  IVP U8685 ( .A(n96), .Z(n10682) );
  IVP U8686 ( .A(n25), .Z(n10717) );
  IVP U8687 ( .A(n30), .Z(n10712) );
  IVP U8688 ( .A(n15), .Z(n10727) );
  IVP U8689 ( .A(n20), .Z(n10722) );
  IVP U8690 ( .A(n10), .Z(n10732) );
  IVP U8691 ( .A(n1), .Z(n10737) );
  IVP U8692 ( .A(n361), .Z(n10417) );
  IVP U8693 ( .A(n362), .Z(n10416) );
  IVP U8694 ( .A(n363), .Z(n10415) );
  IVP U8695 ( .A(n364), .Z(n10414) );
  IVP U8696 ( .A(n662), .Z(n10248) );
  IVP U8697 ( .A(n661), .Z(n10249) );
  IVP U8698 ( .A(n658), .Z(n10252) );
  IVP U8699 ( .A(n663), .Z(n10247) );
  IVP U8700 ( .A(n660), .Z(n10250) );
  IVP U8701 ( .A(n467), .Z(n10366) );
  IVP U8702 ( .A(n407), .Z(n10371) );
  IVP U8703 ( .A(n501), .Z(n10332) );
  IVP U8704 ( .A(n378), .Z(n10400) );
  IVP U8705 ( .A(n383), .Z(n10395) );
  IVP U8706 ( .A(n472), .Z(n10361) );
  IVP U8707 ( .A(n482), .Z(n10351) );
  IVP U8708 ( .A(n506), .Z(n10327) );
  IVP U8709 ( .A(n477), .Z(n10356) );
  IVP U8710 ( .A(n487), .Z(n10346) );
  IVP U8711 ( .A(n388), .Z(n10390) );
  IVP U8712 ( .A(n566), .Z(n10322) );
  IVP U8713 ( .A(n576), .Z(n10312) );
  IVP U8714 ( .A(n374), .Z(n10404) );
  IVP U8715 ( .A(n492), .Z(n10341) );
  IVP U8716 ( .A(n398), .Z(n10380) );
  IVP U8717 ( .A(n393), .Z(n10385) );
  IVP U8718 ( .A(n571), .Z(n10317) );
  IVP U8719 ( .A(n403), .Z(n10375) );
  IVP U8720 ( .A(n581), .Z(n10307) );
  IVP U8721 ( .A(n586), .Z(n10302) );
  IVP U8722 ( .A(n591), .Z(n10297) );
  IVP U8723 ( .A(n408), .Z(n10370) );
  IVP U8724 ( .A(n497), .Z(n10336) );
  IVP U8725 ( .A(n507), .Z(n10326) );
  IVP U8726 ( .A(n502), .Z(n10331) );
  IVP U8727 ( .A(n468), .Z(n10365) );
  IVP U8728 ( .A(n596), .Z(n10292) );
  IVP U8729 ( .A(n473), .Z(n10360) );
  IVP U8730 ( .A(n567), .Z(n10321) );
  IVP U8731 ( .A(n601), .Z(n10287) );
  IVP U8732 ( .A(n478), .Z(n10355) );
  IVP U8733 ( .A(n582), .Z(n10306) );
  IVP U8734 ( .A(n493), .Z(n10340) );
  IVP U8735 ( .A(n587), .Z(n10301) );
  IVP U8736 ( .A(n483), .Z(n10350) );
  IVP U8737 ( .A(n638), .Z(n10272) );
  IVP U8738 ( .A(n606), .Z(n10282) );
  IVP U8739 ( .A(n488), .Z(n10345) );
  IVP U8740 ( .A(n633), .Z(n10277) );
  IVP U8741 ( .A(n572), .Z(n10316) );
  IVP U8742 ( .A(n577), .Z(n10311) );
  IVP U8743 ( .A(n498), .Z(n10335) );
  IVP U8744 ( .A(n643), .Z(n10267) );
  IVP U8745 ( .A(n648), .Z(n10262) );
  IVP U8746 ( .A(n503), .Z(n10330) );
  IVP U8747 ( .A(n592), .Z(n10296) );
  IVP U8748 ( .A(n508), .Z(n10325) );
  IVP U8749 ( .A(n469), .Z(n10364) );
  IVP U8750 ( .A(n474), .Z(n10359) );
  IVP U8751 ( .A(n479), .Z(n10354) );
  IVP U8752 ( .A(n402), .Z(n10376) );
  IVP U8753 ( .A(n392), .Z(n10386) );
  IVP U8754 ( .A(n397), .Z(n10381) );
  IVP U8755 ( .A(n481), .Z(n10352) );
  IVP U8756 ( .A(n471), .Z(n10362) );
  IVP U8757 ( .A(n486), .Z(n10347) );
  IVP U8758 ( .A(n387), .Z(n10391) );
  IVP U8759 ( .A(n496), .Z(n10337) );
  IVP U8760 ( .A(n476), .Z(n10357) );
  IVP U8761 ( .A(n382), .Z(n10396) );
  IVP U8762 ( .A(n491), .Z(n10342) );
  IVP U8763 ( .A(n377), .Z(n10401) );
  IVP U8764 ( .A(n373), .Z(n10405) );
  IVP U8765 ( .A(n368), .Z(n10410) );
  IVP U8766 ( .A(n597), .Z(n10291) );
  IVP U8767 ( .A(n653), .Z(n10257) );
  IVP U8768 ( .A(n484), .Z(n10349) );
  IVP U8769 ( .A(n602), .Z(n10286) );
  IVP U8770 ( .A(n573), .Z(n10315) );
  IVP U8771 ( .A(n568), .Z(n10320) );
  IVP U8772 ( .A(n494), .Z(n10339) );
  IVP U8773 ( .A(n489), .Z(n10344) );
  IVP U8774 ( .A(n607), .Z(n10281) );
  IVP U8775 ( .A(n578), .Z(n10310) );
  IVP U8776 ( .A(n634), .Z(n10276) );
  IVP U8777 ( .A(n639), .Z(n10271) );
  IVP U8778 ( .A(n499), .Z(n10334) );
  IVP U8779 ( .A(n588), .Z(n10300) );
  IVP U8780 ( .A(n583), .Z(n10305) );
  IVP U8781 ( .A(n509), .Z(n10324) );
  IVP U8782 ( .A(n644), .Z(n10266) );
  IVP U8783 ( .A(n504), .Z(n10329) );
  IVP U8784 ( .A(n593), .Z(n10295) );
  IVP U8785 ( .A(n649), .Z(n10261) );
  IVP U8786 ( .A(n654), .Z(n10256) );
  IVP U8787 ( .A(n569), .Z(n10319) );
  IVP U8788 ( .A(n598), .Z(n10290) );
  IVP U8789 ( .A(n574), .Z(n10314) );
  IVP U8790 ( .A(n404), .Z(n10374) );
  IVP U8791 ( .A(n409), .Z(n10369) );
  IVP U8792 ( .A(n401), .Z(n10377) );
  IVP U8793 ( .A(n406), .Z(n10372) );
  IVP U8794 ( .A(n391), .Z(n10387) );
  IVP U8795 ( .A(n372), .Z(n10406) );
  IVP U8796 ( .A(n396), .Z(n10382) );
  IVP U8797 ( .A(n367), .Z(n10411) );
  IVP U8798 ( .A(n466), .Z(n10367) );
  IVP U8799 ( .A(n603), .Z(n10285) );
  IVP U8800 ( .A(n579), .Z(n10309) );
  IVP U8801 ( .A(n608), .Z(n10280) );
  IVP U8802 ( .A(n594), .Z(n10294) );
  IVP U8803 ( .A(n635), .Z(n10275) );
  IVP U8804 ( .A(n640), .Z(n10270) );
  IVP U8805 ( .A(n589), .Z(n10299) );
  IVP U8806 ( .A(n584), .Z(n10304) );
  IVP U8807 ( .A(n645), .Z(n10265) );
  IVP U8808 ( .A(n650), .Z(n10260) );
  IVP U8809 ( .A(n599), .Z(n10289) );
  IVP U8810 ( .A(n394), .Z(n10384) );
  IVP U8811 ( .A(n399), .Z(n10379) );
  IVP U8812 ( .A(n381), .Z(n10397) );
  IVP U8813 ( .A(n376), .Z(n10402) );
  IVP U8814 ( .A(n386), .Z(n10392) );
  IVP U8815 ( .A(n655), .Z(n10255) );
  IVP U8816 ( .A(n604), .Z(n10284) );
  IVP U8817 ( .A(n609), .Z(n10279) );
  IVP U8818 ( .A(n636), .Z(n10274) );
  IVP U8819 ( .A(n384), .Z(n10394) );
  IVP U8820 ( .A(n389), .Z(n10389) );
  IVP U8821 ( .A(n371), .Z(n10407) );
  IVP U8822 ( .A(n366), .Z(n10412) );
  IVP U8823 ( .A(n641), .Z(n10269) );
  IVP U8824 ( .A(n646), .Z(n10264) );
  IVP U8825 ( .A(n379), .Z(n10399) );
  IVP U8826 ( .A(n656), .Z(n10254) );
  IVP U8827 ( .A(n651), .Z(n10259) );
  IVP U8828 ( .A(n657), .Z(n10253) );
  IVP U8829 ( .A(n369), .Z(n10409) );
  IVP U8830 ( .A(n659), .Z(n10251) );
  IVP U8831 ( .A(n580), .Z(n10308) );
  IVP U8832 ( .A(n575), .Z(n10313) );
  IVP U8833 ( .A(n585), .Z(n10303) );
  IVP U8834 ( .A(n590), .Z(n10298) );
  IVP U8835 ( .A(n595), .Z(n10293) );
  IVP U8836 ( .A(n600), .Z(n10288) );
  IVP U8837 ( .A(n605), .Z(n10283) );
  IVP U8838 ( .A(n632), .Z(n10278) );
  IVP U8839 ( .A(n637), .Z(n10273) );
  IVP U8840 ( .A(n642), .Z(n10268) );
  IVP U8841 ( .A(n647), .Z(n10263) );
  IVP U8842 ( .A(n652), .Z(n10258) );
  IVP U8843 ( .A(n485), .Z(n10348) );
  IVP U8844 ( .A(n490), .Z(n10343) );
  IVP U8845 ( .A(n495), .Z(n10338) );
  IVP U8846 ( .A(n570), .Z(n10318) );
  IVP U8847 ( .A(n565), .Z(n10323) );
  IVP U8848 ( .A(n500), .Z(n10333) );
  IVP U8849 ( .A(n505), .Z(n10328) );
  IVP U8850 ( .A(n465), .Z(n10368) );
  IVP U8851 ( .A(n480), .Z(n10353) );
  IVP U8852 ( .A(n470), .Z(n10363) );
  IVP U8853 ( .A(n475), .Z(n10358) );
  IVP U8854 ( .A(n390), .Z(n10388) );
  IVP U8855 ( .A(n395), .Z(n10383) );
  IVP U8856 ( .A(n400), .Z(n10378) );
  IVP U8857 ( .A(n405), .Z(n10373) );
  IVP U8858 ( .A(n380), .Z(n10398) );
  IVP U8859 ( .A(n385), .Z(n10393) );
  IVP U8860 ( .A(n375), .Z(n10403) );
  IVP U8861 ( .A(n370), .Z(n10408) );
  IVP U8862 ( .A(n365), .Z(n10413) );
  IVP U8863 ( .A(n1069), .Z(n1518) );
  IVP U8864 ( .A(n1165), .Z(n1358) );
  IVP U8865 ( .A(n1096), .Z(n1381) );
  IVP U8866 ( .A(n1111), .Z(n1376) );
  IVP U8867 ( .A(n1135), .Z(n1368) );
  IVP U8868 ( .A(n1132), .Z(n1369) );
  IVP U8869 ( .A(n1126), .Z(n1371) );
  IVP U8870 ( .A(n1129), .Z(n1370) );
  IVP U8871 ( .A(n1123), .Z(n1372) );
  IVP U8872 ( .A(n1120), .Z(n1373) );
  IVP U8873 ( .A(n1117), .Z(n1374) );
  IVP U8874 ( .A(n1138), .Z(n1367) );
  IVP U8875 ( .A(n1114), .Z(n1375) );
  IVP U8876 ( .A(n1105), .Z(n1378) );
  IVP U8877 ( .A(n1099), .Z(n1380) );
  IVP U8878 ( .A(n1102), .Z(n1379) );
  IVP U8879 ( .A(n1093), .Z(n1382) );
  IVP U8880 ( .A(n1108), .Z(n1377) );
  IVP U8881 ( .A(n1090), .Z(n1383) );
  IVP U8882 ( .A(n1136), .Z(n1463) );
  IVP U8883 ( .A(n1147), .Z(n1364) );
  IVP U8884 ( .A(n1144), .Z(n1365) );
  IVP U8885 ( .A(n1141), .Z(n1366) );
  IVP U8886 ( .A(n1133), .Z(n1464) );
  IVP U8887 ( .A(n1124), .Z(n1467) );
  IVP U8888 ( .A(n1118), .Z(n1469) );
  IVP U8889 ( .A(n1115), .Z(n1470) );
  IVP U8890 ( .A(n1130), .Z(n1465) );
  IVP U8891 ( .A(n1112), .Z(n1471) );
  IVP U8892 ( .A(n1121), .Z(n1468) );
  IVP U8893 ( .A(n1160), .Z(n1455) );
  IVP U8894 ( .A(n1103), .Z(n1474) );
  IVP U8895 ( .A(n1097), .Z(n1476) );
  IVP U8896 ( .A(n1100), .Z(n1475) );
  IVP U8897 ( .A(n1094), .Z(n1477) );
  IVP U8898 ( .A(n1109), .Z(n1472) );
  IVP U8899 ( .A(n1091), .Z(n1478) );
  IVP U8900 ( .A(n1087), .Z(n1384) );
  IVP U8901 ( .A(n1106), .Z(n1473) );
  IVP U8902 ( .A(n1084), .Z(n1385) );
  IVP U8903 ( .A(n1081), .Z(n1386) );
  IVP U8904 ( .A(n1078), .Z(n1387) );
  IVP U8905 ( .A(n1075), .Z(n1388) );
  IVP U8906 ( .A(n1153), .Z(n1362) );
  IVP U8907 ( .A(n1150), .Z(n1363) );
  IVP U8908 ( .A(n1142), .Z(n1461) );
  IVP U8909 ( .A(n1139), .Z(n1462) );
  IVP U8910 ( .A(n1127), .Z(n1466) );
  IVP U8911 ( .A(n1088), .Z(n1479) );
  IVP U8912 ( .A(n1085), .Z(n1480) );
  IVP U8913 ( .A(n1082), .Z(n1481) );
  IVP U8914 ( .A(n1079), .Z(n1482) );
  IVP U8915 ( .A(n1076), .Z(n1483) );
  IVP U8916 ( .A(n1073), .Z(n1484) );
  IVP U8917 ( .A(n1072), .Z(n1389) );
  IVP U8918 ( .A(n1159), .Z(n1360) );
  IVP U8919 ( .A(n1156), .Z(n1361) );
  IVP U8920 ( .A(n1148), .Z(n1459) );
  IVP U8921 ( .A(n1145), .Z(n1460) );
  IVP U8922 ( .A(n1070), .Z(n1485) );
  IVP U8923 ( .A(n1154), .Z(n1457) );
  IVP U8924 ( .A(n1151), .Z(n1458) );
  IVP U8925 ( .A(n1162), .Z(n1359) );
  IVP U8926 ( .A(n1157), .Z(n1456) );
  IVP U8927 ( .A(n1163), .Z(n1454) );
  IVP U8928 ( .A(n699), .Z(n10211) );
  IVP U8929 ( .A(n736), .Z(n10196) );
  IVP U8930 ( .A(n739), .Z(n10193) );
  IVP U8931 ( .A(n666), .Z(n10244) );
  IVP U8932 ( .A(n669), .Z(n10241) );
  IVP U8933 ( .A(n702), .Z(n10208) );
  IVP U8934 ( .A(n705), .Z(n10205) );
  IVP U8935 ( .A(n687), .Z(n10223) );
  IVP U8936 ( .A(n693), .Z(n10217) );
  IVP U8937 ( .A(n708), .Z(n10202) );
  IVP U8938 ( .A(n675), .Z(n10235) );
  IVP U8939 ( .A(n678), .Z(n10232) );
  IVP U8940 ( .A(n696), .Z(n10214) );
  IVP U8941 ( .A(n684), .Z(n10226) );
  IVP U8942 ( .A(n681), .Z(n10229) );
  IVP U8943 ( .A(n733), .Z(n10199) );
  IVP U8944 ( .A(n742), .Z(n10190) );
  IVP U8945 ( .A(n672), .Z(n10238) );
  IVP U8946 ( .A(n690), .Z(n10220) );
  IVP U8947 ( .A(n751), .Z(n10181) );
  IVP U8948 ( .A(n754), .Z(n10178) );
  IVP U8949 ( .A(n790), .Z(n10142) );
  IVP U8950 ( .A(n748), .Z(n10184) );
  IVP U8951 ( .A(n745), .Z(n10187) );
  IVP U8952 ( .A(n760), .Z(n10172) );
  IVP U8953 ( .A(n757), .Z(n10175) );
  IVP U8954 ( .A(n769), .Z(n10163) );
  IVP U8955 ( .A(n763), .Z(n10169) );
  IVP U8956 ( .A(n778), .Z(n10154) );
  IVP U8957 ( .A(n772), .Z(n10160) );
  IVP U8958 ( .A(n787), .Z(n10145) );
  IVP U8959 ( .A(n781), .Z(n10151) );
  IVP U8960 ( .A(n775), .Z(n10157) );
  IVP U8961 ( .A(n793), .Z(n10139) );
  IVP U8962 ( .A(n766), .Z(n10166) );
  IVP U8963 ( .A(n784), .Z(n10148) );
  IVP U8964 ( .A(n796), .Z(n10136) );
  IVP U8965 ( .A(n805), .Z(n10127) );
  IVP U8966 ( .A(n814), .Z(n10118) );
  IVP U8967 ( .A(n823), .Z(n10109) );
  IVP U8968 ( .A(n817), .Z(n10115) );
  IVP U8969 ( .A(n799), .Z(n10133) );
  IVP U8970 ( .A(n802), .Z(n10130) );
  IVP U8971 ( .A(n808), .Z(n10124) );
  IVP U8972 ( .A(n811), .Z(n10121) );
  IVP U8973 ( .A(n820), .Z(n10112) );
  IVP U8974 ( .A(n826), .Z(n10106) );
  IVP U8975 ( .A(n829), .Z(n10103) );
  IVP U8976 ( .A(n838), .Z(n10094) );
  IVP U8977 ( .A(n832), .Z(n10100) );
  IVP U8978 ( .A(n835), .Z(n10097) );
  IVP U8979 ( .A(n844), .Z(n10088) );
  IVP U8980 ( .A(n841), .Z(n10091) );
  IVP U8981 ( .A(n847), .Z(n10085) );
  IVP U8982 ( .A(n850), .Z(n10082) );
  IVP U8983 ( .A(n853), .Z(n10079) );
  IVP U8984 ( .A(n859), .Z(n10073) );
  IVP U8985 ( .A(n856), .Z(n10076) );
  IVP U8986 ( .A(n862), .Z(n10070) );
  IVP U8987 ( .A(n865), .Z(n10067) );
  IVP U8988 ( .A(n868), .Z(n10064) );
  IVP U8989 ( .A(n874), .Z(n10058) );
  IVP U8990 ( .A(n871), .Z(n10061) );
  IVP U8991 ( .A(n804), .Z(n10128) );
  IVP U8992 ( .A(n801), .Z(n10131) );
  IVP U8993 ( .A(n665), .Z(n10245) );
  IVP U8994 ( .A(n668), .Z(n10242) );
  IVP U8995 ( .A(n671), .Z(n10239) );
  IVP U8996 ( .A(n770), .Z(n10162) );
  IVP U8997 ( .A(n773), .Z(n10159) );
  IVP U8998 ( .A(n686), .Z(n10224) );
  IVP U8999 ( .A(n689), .Z(n10221) );
  IVP U9000 ( .A(n797), .Z(n10135) );
  IVP U9001 ( .A(n800), .Z(n10132) );
  IVP U9002 ( .A(n812), .Z(n10120) );
  IVP U9003 ( .A(n803), .Z(n10129) );
  IVP U9004 ( .A(n809), .Z(n10123) );
  IVP U9005 ( .A(n806), .Z(n10126) );
  IVP U9006 ( .A(n750), .Z(n10182) );
  IVP U9007 ( .A(n792), .Z(n10140) );
  IVP U9008 ( .A(n753), .Z(n10179) );
  IVP U9009 ( .A(n789), .Z(n10143) );
  IVP U9010 ( .A(n824), .Z(n10108) );
  IVP U9011 ( .A(n830), .Z(n10102) );
  IVP U9012 ( .A(n827), .Z(n10105) );
  IVP U9013 ( .A(n786), .Z(n10146) );
  IVP U9014 ( .A(n795), .Z(n10137) );
  IVP U9015 ( .A(n854), .Z(n10078) );
  IVP U9016 ( .A(n857), .Z(n10075) );
  IVP U9017 ( .A(n798), .Z(n10134) );
  IVP U9018 ( .A(n860), .Z(n10072) );
  IVP U9019 ( .A(n807), .Z(n10125) );
  IVP U9020 ( .A(n700), .Z(n10210) );
  IVP U9021 ( .A(n749), .Z(n10183) );
  IVP U9022 ( .A(n755), .Z(n10177) );
  IVP U9023 ( .A(n752), .Z(n10180) );
  IVP U9024 ( .A(n776), .Z(n10156) );
  IVP U9025 ( .A(n758), .Z(n10174) );
  IVP U9026 ( .A(n674), .Z(n10236) );
  IVP U9027 ( .A(n761), .Z(n10171) );
  IVP U9028 ( .A(n677), .Z(n10233) );
  IVP U9029 ( .A(n767), .Z(n10165) );
  IVP U9030 ( .A(n764), .Z(n10168) );
  IVP U9031 ( .A(n788), .Z(n10144) );
  IVP U9032 ( .A(n695), .Z(n10215) );
  IVP U9033 ( .A(n692), .Z(n10218) );
  IVP U9034 ( .A(n683), .Z(n10227) );
  IVP U9035 ( .A(n680), .Z(n10230) );
  IVP U9036 ( .A(n779), .Z(n10153) );
  IVP U9037 ( .A(n791), .Z(n10141) );
  IVP U9038 ( .A(n698), .Z(n10212) );
  IVP U9039 ( .A(n782), .Z(n10150) );
  IVP U9040 ( .A(n794), .Z(n10138) );
  IVP U9041 ( .A(n701), .Z(n10209) );
  IVP U9042 ( .A(n785), .Z(n10147) );
  IVP U9043 ( .A(n704), .Z(n10206) );
  IVP U9044 ( .A(n707), .Z(n10203) );
  IVP U9045 ( .A(n732), .Z(n10200) );
  IVP U9046 ( .A(n735), .Z(n10197) );
  IVP U9047 ( .A(n741), .Z(n10191) );
  IVP U9048 ( .A(n738), .Z(n10194) );
  IVP U9049 ( .A(n759), .Z(n10173) );
  IVP U9050 ( .A(n756), .Z(n10176) );
  IVP U9051 ( .A(n747), .Z(n10185) );
  IVP U9052 ( .A(n744), .Z(n10188) );
  IVP U9053 ( .A(n821), .Z(n10111) );
  IVP U9054 ( .A(n815), .Z(n10117) );
  IVP U9055 ( .A(n818), .Z(n10114) );
  IVP U9056 ( .A(n768), .Z(n10164) );
  IVP U9057 ( .A(n771), .Z(n10161) );
  IVP U9058 ( .A(n762), .Z(n10170) );
  IVP U9059 ( .A(n765), .Z(n10167) );
  IVP U9060 ( .A(n833), .Z(n10099) );
  IVP U9061 ( .A(n836), .Z(n10096) );
  IVP U9062 ( .A(n842), .Z(n10090) );
  IVP U9063 ( .A(n839), .Z(n10093) );
  IVP U9064 ( .A(n780), .Z(n10152) );
  IVP U9065 ( .A(n777), .Z(n10155) );
  IVP U9066 ( .A(n774), .Z(n10158) );
  IVP U9067 ( .A(n783), .Z(n10149) );
  IVP U9068 ( .A(n845), .Z(n10087) );
  IVP U9069 ( .A(n866), .Z(n10066) );
  IVP U9070 ( .A(n869), .Z(n10063) );
  IVP U9071 ( .A(n863), .Z(n10069) );
  IVP U9072 ( .A(n851), .Z(n10081) );
  IVP U9073 ( .A(n848), .Z(n10084) );
  IVP U9074 ( .A(n872), .Z(n10060) );
  IVP U9075 ( .A(n813), .Z(n10119) );
  IVP U9076 ( .A(n810), .Z(n10122) );
  IVP U9077 ( .A(n819), .Z(n10113) );
  IVP U9078 ( .A(n816), .Z(n10116) );
  IVP U9079 ( .A(n843), .Z(n10089) );
  IVP U9080 ( .A(n846), .Z(n10086) );
  IVP U9081 ( .A(n855), .Z(n10077) );
  IVP U9082 ( .A(n664), .Z(n10246) );
  IVP U9083 ( .A(n697), .Z(n10213) );
  IVP U9084 ( .A(n694), .Z(n10216) );
  IVP U9085 ( .A(n703), .Z(n10207) );
  IVP U9086 ( .A(n740), .Z(n10192) );
  IVP U9087 ( .A(n709), .Z(n10201) );
  IVP U9088 ( .A(n706), .Z(n10204) );
  IVP U9089 ( .A(n737), .Z(n10195) );
  IVP U9090 ( .A(n734), .Z(n10198) );
  IVP U9091 ( .A(n743), .Z(n10189) );
  IVP U9092 ( .A(n746), .Z(n10186) );
  IVP U9093 ( .A(n831), .Z(n10101) );
  IVP U9094 ( .A(n828), .Z(n10104) );
  IVP U9095 ( .A(n825), .Z(n10107) );
  IVP U9096 ( .A(n822), .Z(n10110) );
  IVP U9097 ( .A(n837), .Z(n10095) );
  IVP U9098 ( .A(n834), .Z(n10098) );
  IVP U9099 ( .A(n840), .Z(n10092) );
  IVP U9100 ( .A(n852), .Z(n10080) );
  IVP U9101 ( .A(n849), .Z(n10083) );
  IVP U9102 ( .A(n858), .Z(n10074) );
  IVP U9103 ( .A(n861), .Z(n10071) );
  IVP U9104 ( .A(n870), .Z(n10062) );
  IVP U9105 ( .A(n670), .Z(n10240) );
  IVP U9106 ( .A(n667), .Z(n10243) );
  IVP U9107 ( .A(n673), .Z(n10237) );
  IVP U9108 ( .A(n676), .Z(n10234) );
  IVP U9109 ( .A(n679), .Z(n10231) );
  IVP U9110 ( .A(n685), .Z(n10225) );
  IVP U9111 ( .A(n682), .Z(n10228) );
  IVP U9112 ( .A(n691), .Z(n10219) );
  IVP U9113 ( .A(n688), .Z(n10222) );
  IVP U9114 ( .A(n867), .Z(n10065) );
  IVP U9115 ( .A(n864), .Z(n10068) );
  IVP U9116 ( .A(n873), .Z(n10059) );
endmodule


module tx_DW01_add_64_0 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   \carry[63] , \carry[62] , \carry[61] , \carry[60] , \carry[59] ,
         \carry[58] , \carry[57] , \carry[56] , \carry[55] , \carry[54] ,
         \carry[53] , \carry[52] , \carry[51] , \carry[50] , \carry[49] ,
         \carry[48] , \carry[47] , \carry[46] , \carry[45] , \carry[44] ,
         \carry[43] , \carry[42] , \carry[41] , \carry[40] , \carry[39] ,
         \carry[38] , \carry[37] , \carry[36] , \carry[35] , \carry[34] ,
         \carry[33] , \carry[32] , \carry[31] , \carry[30] , \carry[29] ,
         \carry[28] , \carry[27] , \carry[26] , \carry[25] , \carry[24] ,
         \carry[23] , \carry[22] , \carry[21] , \carry[20] , \carry[19] ,
         \carry[18] , \carry[17] , \carry[16] , \carry[15] , \carry[14] ,
         \carry[13] , \carry[12] , \carry[11] , \carry[10] , \carry[9] ,
         \carry[8] , \carry[7] , \carry[6] , \carry[5] , \carry[4] ,
         \carry[3] , \carry[2] , \carry[1] ;

  FA1A U1_1 ( .CI(\carry[1] ), .A(A[1]), .B(B[1]), .S(SUM[1]), .CO(\carry[2] )
         );
  FA1A U1_2 ( .CI(\carry[2] ), .A(A[2]), .B(B[2]), .S(SUM[2]), .CO(\carry[3] )
         );
  FA1A U1_3 ( .CI(\carry[3] ), .A(A[3]), .B(B[3]), .S(SUM[3]), .CO(\carry[4] )
         );
  FA1A U1_4 ( .CI(\carry[4] ), .A(A[4]), .B(B[4]), .S(SUM[4]), .CO(\carry[5] )
         );
  FA1A U1_5 ( .CI(\carry[5] ), .A(A[5]), .B(B[5]), .S(SUM[5]), .CO(\carry[6] )
         );
  FA1A U1_6 ( .CI(\carry[6] ), .A(A[6]), .B(B[6]), .S(SUM[6]), .CO(\carry[7] )
         );
  FA1A U1_7 ( .CI(\carry[7] ), .A(A[7]), .B(B[7]), .S(SUM[7]), .CO(\carry[8] )
         );
  FA1A U1_8 ( .CI(\carry[8] ), .A(A[8]), .B(B[8]), .S(SUM[8]), .CO(\carry[9] )
         );
  FA1A U1_9 ( .CI(\carry[9] ), .A(A[9]), .B(B[9]), .S(SUM[9]), .CO(\carry[10] ) );
  FA1A U1_10 ( .CI(\carry[10] ), .A(A[10]), .B(B[10]), .S(SUM[10]), .CO(
        \carry[11] ) );
  FA1A U1_11 ( .CI(\carry[11] ), .A(A[11]), .B(B[11]), .S(SUM[11]), .CO(
        \carry[12] ) );
  FA1A U1_12 ( .CI(\carry[12] ), .A(A[12]), .B(B[12]), .S(SUM[12]), .CO(
        \carry[13] ) );
  FA1A U1_13 ( .CI(\carry[13] ), .A(A[13]), .B(B[13]), .S(SUM[13]), .CO(
        \carry[14] ) );
  FA1A U1_14 ( .CI(\carry[14] ), .A(A[14]), .B(B[14]), .S(SUM[14]), .CO(
        \carry[15] ) );
  FA1A U1_15 ( .CI(\carry[15] ), .A(A[15]), .B(B[15]), .S(SUM[15]), .CO(
        \carry[16] ) );
  FA1A U1_16 ( .CI(\carry[16] ), .A(A[16]), .B(B[16]), .S(SUM[16]), .CO(
        \carry[17] ) );
  FA1A U1_17 ( .CI(\carry[17] ), .A(A[17]), .B(B[17]), .S(SUM[17]), .CO(
        \carry[18] ) );
  FA1A U1_18 ( .CI(\carry[18] ), .A(A[18]), .B(B[18]), .S(SUM[18]), .CO(
        \carry[19] ) );
  FA1A U1_19 ( .CI(\carry[19] ), .A(A[19]), .B(B[19]), .S(SUM[19]), .CO(
        \carry[20] ) );
  FA1A U1_20 ( .CI(\carry[20] ), .A(A[20]), .B(B[20]), .S(SUM[20]), .CO(
        \carry[21] ) );
  FA1A U1_21 ( .CI(\carry[21] ), .A(A[21]), .B(B[21]), .S(SUM[21]), .CO(
        \carry[22] ) );
  FA1A U1_22 ( .CI(\carry[22] ), .A(A[22]), .B(B[22]), .S(SUM[22]), .CO(
        \carry[23] ) );
  FA1A U1_23 ( .CI(\carry[23] ), .A(A[23]), .B(B[23]), .S(SUM[23]), .CO(
        \carry[24] ) );
  FA1A U1_24 ( .CI(\carry[24] ), .A(A[24]), .B(B[24]), .S(SUM[24]), .CO(
        \carry[25] ) );
  FA1A U1_25 ( .CI(\carry[25] ), .A(A[25]), .B(B[25]), .S(SUM[25]), .CO(
        \carry[26] ) );
  FA1A U1_26 ( .CI(\carry[26] ), .A(A[26]), .B(B[26]), .S(SUM[26]), .CO(
        \carry[27] ) );
  FA1A U1_27 ( .CI(\carry[27] ), .A(A[27]), .B(B[27]), .S(SUM[27]), .CO(
        \carry[28] ) );
  FA1A U1_28 ( .CI(\carry[28] ), .A(A[28]), .B(B[28]), .S(SUM[28]), .CO(
        \carry[29] ) );
  FA1A U1_29 ( .CI(\carry[29] ), .A(A[29]), .B(B[29]), .S(SUM[29]), .CO(
        \carry[30] ) );
  FA1A U1_30 ( .CI(\carry[30] ), .A(A[30]), .B(B[30]), .S(SUM[30]), .CO(
        \carry[31] ) );
  FA1A U1_31 ( .CI(\carry[31] ), .A(A[31]), .B(B[31]), .S(SUM[31]), .CO(
        \carry[32] ) );
  FA1A U1_32 ( .CI(\carry[32] ), .A(A[32]), .B(B[32]), .S(SUM[32]), .CO(
        \carry[33] ) );
  FA1A U1_33 ( .CI(\carry[33] ), .A(A[33]), .B(B[33]), .S(SUM[33]), .CO(
        \carry[34] ) );
  FA1A U1_34 ( .CI(\carry[34] ), .A(A[34]), .B(B[34]), .S(SUM[34]), .CO(
        \carry[35] ) );
  FA1A U1_35 ( .CI(\carry[35] ), .A(A[35]), .B(B[35]), .S(SUM[35]), .CO(
        \carry[36] ) );
  FA1A U1_36 ( .CI(\carry[36] ), .A(A[36]), .B(B[36]), .S(SUM[36]), .CO(
        \carry[37] ) );
  FA1A U1_37 ( .CI(\carry[37] ), .A(A[37]), .B(B[37]), .S(SUM[37]), .CO(
        \carry[38] ) );
  FA1A U1_38 ( .CI(\carry[38] ), .A(A[38]), .B(B[38]), .S(SUM[38]), .CO(
        \carry[39] ) );
  FA1A U1_39 ( .CI(\carry[39] ), .A(A[39]), .B(B[39]), .S(SUM[39]), .CO(
        \carry[40] ) );
  FA1A U1_40 ( .CI(\carry[40] ), .A(A[40]), .B(B[40]), .S(SUM[40]), .CO(
        \carry[41] ) );
  FA1A U1_41 ( .CI(\carry[41] ), .A(A[41]), .B(B[41]), .S(SUM[41]), .CO(
        \carry[42] ) );
  FA1A U1_42 ( .CI(\carry[42] ), .A(A[42]), .B(B[42]), .S(SUM[42]), .CO(
        \carry[43] ) );
  FA1A U1_43 ( .CI(\carry[43] ), .A(A[43]), .B(B[43]), .S(SUM[43]), .CO(
        \carry[44] ) );
  FA1A U1_44 ( .CI(\carry[44] ), .A(A[44]), .B(B[44]), .S(SUM[44]), .CO(
        \carry[45] ) );
  FA1A U1_45 ( .CI(\carry[45] ), .A(A[45]), .B(B[45]), .S(SUM[45]), .CO(
        \carry[46] ) );
  FA1A U1_46 ( .CI(\carry[46] ), .A(A[46]), .B(B[46]), .S(SUM[46]), .CO(
        \carry[47] ) );
  FA1A U1_47 ( .CI(\carry[47] ), .A(A[47]), .B(B[47]), .S(SUM[47]), .CO(
        \carry[48] ) );
  FA1A U1_48 ( .CI(\carry[48] ), .A(A[48]), .B(B[48]), .S(SUM[48]), .CO(
        \carry[49] ) );
  FA1A U1_49 ( .CI(\carry[49] ), .A(A[49]), .B(B[49]), .S(SUM[49]), .CO(
        \carry[50] ) );
  FA1A U1_50 ( .CI(\carry[50] ), .A(A[50]), .B(B[50]), .S(SUM[50]), .CO(
        \carry[51] ) );
  FA1A U1_51 ( .CI(\carry[51] ), .A(A[51]), .B(B[51]), .S(SUM[51]), .CO(
        \carry[52] ) );
  FA1A U1_52 ( .CI(\carry[52] ), .A(A[52]), .B(B[52]), .S(SUM[52]), .CO(
        \carry[53] ) );
  FA1A U1_53 ( .CI(\carry[53] ), .A(A[53]), .B(B[53]), .S(SUM[53]), .CO(
        \carry[54] ) );
  FA1A U1_54 ( .CI(\carry[54] ), .A(A[54]), .B(B[54]), .S(SUM[54]), .CO(
        \carry[55] ) );
  FA1A U1_55 ( .CI(\carry[55] ), .A(A[55]), .B(B[55]), .S(SUM[55]), .CO(
        \carry[56] ) );
  FA1A U1_56 ( .CI(\carry[56] ), .A(A[56]), .B(B[56]), .S(SUM[56]), .CO(
        \carry[57] ) );
  FA1A U1_57 ( .CI(\carry[57] ), .A(A[57]), .B(B[57]), .S(SUM[57]), .CO(
        \carry[58] ) );
  FA1A U1_58 ( .CI(\carry[58] ), .A(A[58]), .B(B[58]), .S(SUM[58]), .CO(
        \carry[59] ) );
  FA1A U1_59 ( .CI(\carry[59] ), .A(A[59]), .B(B[59]), .S(SUM[59]), .CO(
        \carry[60] ) );
  FA1A U1_60 ( .CI(\carry[60] ), .A(A[60]), .B(B[60]), .S(SUM[60]), .CO(
        \carry[61] ) );
  FA1A U1_61 ( .CI(\carry[61] ), .A(A[61]), .B(B[61]), .S(SUM[61]), .CO(
        \carry[62] ) );
  FA1A U1_62 ( .CI(\carry[62] ), .A(A[62]), .B(B[62]), .S(SUM[62]), .CO(
        \carry[63] ) );
  EO3P U1_63 ( .A(A[63]), .B(B[63]), .C(\carry[63] ), .Z(SUM[63]) );
  AN2 U4 ( .A(B[0]), .B(A[0]), .Z(\carry[1] ) );
  EO U5 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
endmodule


module tx ( in1, in2, mult_out, add_out );
  input [63:0] in1;
  input [63:0] in2;
  output [127:0] mult_out;
  output [63:0] add_out;


  tx_DW_mult_uns_1 mult_12 ( .a(in1), .b(in2), .product(mult_out) );
  tx_DW01_add_64_0 add_13 ( .A(in1), .B(in2), .CI(1'b0), .SUM(add_out) );
endmodule


module hierA ( sum_0, dec_tap_1, sum_1, in1, in2, mult_out, add_out );
  input [9:0] sum_0;
  input [9:0] dec_tap_1;
  output [9:0] sum_1;
  input [63:0] in1;
  input [63:0] in2;
  output [127:0] mult_out;
  output [63:0] add_out;


  rx U1 ( .sum_0(sum_0), .dec_tap_1(dec_tap_1), .sum_1(sum_1) );
  tx U2 ( .in1(in1), .in2(in2), .mult_out(mult_out), .add_out(add_out) );
endmodule


module hierB ( sum_0, dec_tap_1, sum_1, in1, in2, mult_out, add_out );
  input [9:0] sum_0;
  input [9:0] dec_tap_1;
  output [9:0] sum_1;
  input [63:0] in1;
  input [63:0] in2;
  output [127:0] mult_out;
  output [63:0] add_out;


  hierA U1 ( .sum_0(sum_0), .dec_tap_1(dec_tap_1), .sum_1(sum_1), .in1(in1), 
        .in2(in2), .mult_out(mult_out), .add_out(add_out) );
endmodule


module hierC ( sum_0, dec_tap_1, sum_1, in1, in2, mult_out, add_out );
  input [9:0] sum_0;
  input [9:0] dec_tap_1;
  output [9:0] sum_1;
  input [63:0] in1;
  input [63:0] in2;
  output [127:0] mult_out;
  output [63:0] add_out;


  hierB U1 ( .sum_0(sum_0), .dec_tap_1(dec_tap_1), .sum_1(sum_1), .in1(in1), 
        .in2(in2), .mult_out(mult_out), .add_out(add_out) );
endmodule


module top ( sum_0, dec_tap_1, sum_1, in1, in2, mult_out, add_out );
  input [9:0] sum_0;
  input [9:0] dec_tap_1;
  output [9:0] sum_1;
  input [63:0] in1;
  input [63:0] in2;
  output [127:0] mult_out;
  output [63:0] add_out;


  hierC U1 ( .sum_0(sum_0), .dec_tap_1(dec_tap_1), .sum_1(sum_1), .in1(in1), 
        .in2(in2), .mult_out(mult_out), .add_out(add_out) );
endmodule

