library verilog;
use verilog.vl_types.all;
entity routines is
end routines;
