
module BIST_AWid5_DWid32_DW01_inc_5 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_4 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_2 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32 ( DataO, Addr, ReadCmd, WriteCmd, Testing, TestOK, 
        DataI, DoSelfTest, ParityErr, Clk, Reset );
  output [31:0] DataO;
  output [4:0] Addr;
  input [31:0] DataI;
  input DoSelfTest, ParityErr, Clk, Reset;
  output ReadCmd, WriteCmd, Testing, TestOK;
  wire   n519, TDone5, TDone3, TDone1, TRes5, TRes3, TRes1, AllDoner, N132,
         N138, N145, N151, N158, N165, N170, N172, N184, N185, N186, N203,
         N204, N205, N206, N208, N210, N211, N212, N214, N216, N217, N218,
         N219, N220, N221, N226, N227, N228, N229, N230, N231, N233, N279,
         N280, N281, N282, N284, N285, N286, N287, N288, N289, N319, N320,
         N321, N322, N323, N324, N326, N364, N370, N371, N372, N373, N374,
         N375, N404, N405, N406, N407, N408, N409, N411, N449, N455, N456,
         N457, N458, N459, N460, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n176, n177, n178, n179, n180, n181, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n237, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n175, n182, n225,
         n236, n238, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518;
  wire   [6:1] TestDone;
  wire   [2:0] TestNo;
  wire   [4:0] Addr1;
  wire   [4:0] Addr3;
  wire   [4:0] Addr5;
  wire   [31:0] DataO1;
  wire   [2:0] State;
  wire   [4:0] i1;
  wire   [4:0] i2;
  wire   [4:0] i3;
  wire   [4:0] i4;
  wire   [4:0] i5;
  wire   [4:0] i6;

  DFND1 \Addr2_reg[3]  ( .D(n282), .CPN(Clk), .QN(n235) );
  DFND1 \Addr2_reg[0]  ( .D(n280), .CPN(Clk), .QN(n233) );
  DFND1 \Addr2_reg[1]  ( .D(n278), .CPN(Clk), .QN(n231) );
  DFND1 \Addr2_reg[2]  ( .D(n276), .CPN(Clk), .QN(n229) );
  DFND1 \Addr2_reg[4]  ( .D(n274), .CPN(Clk), .QN(n227) );
  DFND1 \Addr4_reg[3]  ( .D(n269), .CPN(Clk), .QN(n223) );
  DFND1 \Addr4_reg[0]  ( .D(n267), .CPN(Clk), .QN(n221) );
  DFND1 \Addr4_reg[1]  ( .D(n265), .CPN(Clk), .QN(n219) );
  DFND1 \Addr4_reg[2]  ( .D(n263), .CPN(Clk), .QN(n217) );
  DFND1 \Addr4_reg[4]  ( .D(n261), .CPN(Clk), .QN(n215) );
  DFND1 \Addr6_reg[3]  ( .D(n250), .CPN(Clk), .QN(n211) );
  DFND1 \Addr6_reg[0]  ( .D(n248), .CPN(Clk), .QN(n209) );
  DFND1 \Addr6_reg[1]  ( .D(n246), .CPN(Clk), .QN(n207) );
  DFND1 \Addr6_reg[2]  ( .D(n244), .CPN(Clk), .QN(n205) );
  DFND1 \Addr6_reg[4]  ( .D(n242), .CPN(Clk), .QN(n203) );
  MOAI22D1 U6 ( .A1(n202), .A2(n72), .B1(n73), .B2(N460), .ZN(n241) );
  MOAI22D1 U9 ( .A1(n204), .A2(n73), .B1(N459), .B2(n73), .ZN(n243) );
  MOAI22D1 U11 ( .A1(n206), .A2(n73), .B1(N457), .B2(n73), .ZN(n245) );
  MOAI22D1 U13 ( .A1(n208), .A2(n73), .B1(N456), .B2(n73), .ZN(n247) );
  MOAI22D1 U15 ( .A1(n210), .A2(n73), .B1(N455), .B2(n73), .ZN(n249) );
  MOAI22D1 U47 ( .A1(n212), .A2(n73), .B1(N458), .B2(n73), .ZN(n251) );
  AO21D1 U51 ( .A1(N411), .A2(N409), .B(TDone5), .Z(n253) );
  AO21D1 U52 ( .A1(N411), .A2(N409), .B(TRes5), .Z(n254) );
  AO21D1 U53 ( .A1(N326), .A2(N324), .B(TDone3), .Z(n255) );
  AO21D1 U55 ( .A1(N233), .A2(N231), .B(TDone1), .Z(n257) );
  AO21D1 U56 ( .A1(N233), .A2(N231), .B(TRes1), .Z(n258) );
  MOAI22D1 U59 ( .A1(n214), .A2(n85), .B1(n86), .B2(N375), .ZN(n260) );
  MOAI22D1 U62 ( .A1(n216), .A2(n86), .B1(N374), .B2(n86), .ZN(n262) );
  MOAI22D1 U64 ( .A1(n218), .A2(n86), .B1(N372), .B2(n86), .ZN(n264) );
  MOAI22D1 U66 ( .A1(n220), .A2(n86), .B1(N371), .B2(n86), .ZN(n266) );
  MOAI22D1 U68 ( .A1(n222), .A2(n86), .B1(N370), .B2(n86), .ZN(n268) );
  MOAI22D1 U72 ( .A1(n224), .A2(n86), .B1(N373), .B2(n86), .ZN(n270) );
  MOAI22D1 U90 ( .A1(n226), .A2(n103), .B1(n104), .B2(N289), .ZN(n272) );
  MOAI22D1 U95 ( .A1(n228), .A2(n104), .B1(N288), .B2(n104), .ZN(n275) );
  MOAI22D1 U97 ( .A1(n230), .A2(n104), .B1(N286), .B2(n104), .ZN(n277) );
  MOAI22D1 U99 ( .A1(n232), .A2(n104), .B1(N285), .B2(n104), .ZN(n279) );
  MOAI22D1 U101 ( .A1(n234), .A2(n104), .B1(N284), .B2(n104), .ZN(n281) );
  MOAI22D1 U105 ( .A1(n237), .A2(n104), .B1(N287), .B2(n104), .ZN(n283) );
  OR4D1 U118 ( .A1(DataI[24]), .A2(DataI[25]), .A3(DataI[26]), .A4(DataI[27]), 
        .Z(n118) );
  OR4D1 U119 ( .A1(DataI[28]), .A2(DataI[29]), .A3(DataI[2]), .A4(DataI[30]), 
        .Z(n117) );
  OR4D1 U120 ( .A1(DataI[31]), .A2(DataI[3]), .A3(DataI[4]), .A4(DataI[5]), 
        .Z(n116) );
  OR4D1 U121 ( .A1(DataI[6]), .A2(DataI[7]), .A3(DataI[8]), .A4(DataI[9]), .Z(
        n115) );
  OR4D1 U123 ( .A1(DataI[0]), .A2(DataI[10]), .A3(DataI[11]), .A4(DataI[12]), 
        .Z(n122) );
  OR4D1 U124 ( .A1(DataI[13]), .A2(DataI[14]), .A3(DataI[15]), .A4(DataI[16]), 
        .Z(n121) );
  OR4D1 U125 ( .A1(DataI[17]), .A2(DataI[18]), .A3(DataI[19]), .A4(DataI[1]), 
        .Z(n120) );
  OR4D1 U126 ( .A1(DataI[20]), .A2(DataI[21]), .A3(DataI[22]), .A4(DataI[23]), 
        .Z(n119) );
  OR3D1 U137 ( .A1(n214), .A2(n202), .A3(n226), .Z(n129) );
  IAO21D1 U144 ( .A1(n226), .A2(n457), .B(n145), .ZN(n144) );
  IAO21D1 U163 ( .A1(n168), .A2(n130), .B(n169), .ZN(n165) );
  OA222D1 U188 ( .A1(n145), .A2(TestDone[2]), .B1(n180), .B2(TestDone[4]), 
        .C1(n152), .C2(TestDone[6]), .Z(n179) );
  BIST_AWid5_DWid32_DW01_inc_0 \TestPhase06/DelayedSample/add_551  ( .A(i6), 
        .SUM({N459, N458, N457, N456, N455}) );
  BIST_AWid5_DWid32_DW01_inc_1 \TestPhase05/add_513  ( .A(i5), .SUM({N408, 
        N407, N406, N405, N404}) );
  BIST_AWid5_DWid32_DW01_inc_2 \TestPhase04/DelayedSample/add_483  ( .A(i4), 
        .SUM({N374, N373, N372, N371, N370}) );
  BIST_AWid5_DWid32_DW01_inc_3 \TestPhase03/add_445  ( .A(i3), .SUM({N323, 
        N322, N321, N320, N319}) );
  BIST_AWid5_DWid32_DW01_inc_4 \TestPhase02/DelayedSample/add_415  ( .A(i2), 
        .SUM({N288, N287, N286, N285, N284}) );
  BIST_AWid5_DWid32_DW01_inc_5 \TestPhase01/add_373  ( .A(i1), .SUM({N230, 
        N229, N228, N227, N226}) );
  EDFCNQD1 TestOKr_reg ( .D(N220), .E(N219), .CP(Clk), .CDN(n460), .Q(n519) );
  EDFQD1 \DataO1_reg[9]  ( .D(i1[1]), .E(n1), .CP(Clk), .Q(DataO1[9]) );
  EDFQD1 \DataO1_reg[3]  ( .D(i1[3]), .E(n1), .CP(Clk), .Q(DataO1[3]) );
  EDFQD1 \DataO1_reg[1]  ( .D(i1[1]), .E(n1), .CP(Clk), .Q(DataO1[1]) );
  EDFQD1 \DataO1_reg[0]  ( .D(i1[0]), .E(n1), .CP(Clk), .Q(DataO1[0]) );
  EDFQD1 \DataO1_reg[2]  ( .D(i1[2]), .E(n1), .CP(Clk), .Q(DataO1[2]) );
  EDFQD1 \DataO1_reg[4]  ( .D(i1[4]), .E(n1), .CP(Clk), .Q(DataO1[4]) );
  EDFQD1 \DataO1_reg[8]  ( .D(i1[0]), .E(n1), .CP(Clk), .Q(DataO1[8]) );
  DFNSND1 Wait2_reg ( .D(n273), .CPN(Clk), .SDN(n35), .QN(n106) );
  DFNSND1 Wait4_reg ( .D(n271), .CPN(Clk), .SDN(n35), .QN(n90) );
  DFNSND1 Wait6_reg ( .D(n252), .CPN(Clk), .SDN(n35), .QN(n79) );
  DFNCND1 \i4_reg[4]  ( .D(n262), .CPN(Clk), .CDN(n461), .Q(i4[4]), .QN(n216)
         );
  DFNCND1 \i6_reg[4]  ( .D(n243), .CPN(Clk), .CDN(n4), .Q(i6[4]), .QN(n204) );
  EDFCNQD1 WriteCmdr_reg ( .D(N186), .E(N221), .CP(Clk), .CDN(n460), .Q(
        WriteCmd) );
  EDFCNQD1 ReadCmdr_reg ( .D(N185), .E(N221), .CP(Clk), .CDN(n460), .Q(ReadCmd) );
  EDFCNQD1 \i3_reg[4]  ( .D(N323), .E(N326), .CP(Clk), .CDN(n461), .Q(i3[4])
         );
  EDFCNQD1 \i5_reg[4]  ( .D(N408), .E(N411), .CP(Clk), .CDN(n461), .Q(i5[4])
         );
  DFCNQD1 TDone3_reg ( .D(n255), .CP(Clk), .CDN(n461), .Q(TDone3) );
  DFCNQD1 TDone5_reg ( .D(n253), .CP(Clk), .CDN(n461), .Q(TDone5) );
  DFNCND1 \i4_reg[3]  ( .D(n270), .CPN(Clk), .CDN(n461), .Q(i4[3]), .QN(n224)
         );
  DFNCND1 \i4_reg[1]  ( .D(n266), .CPN(Clk), .CDN(n461), .Q(i4[1]), .QN(n220)
         );
  DFNCND1 \i4_reg[2]  ( .D(n264), .CPN(Clk), .CDN(n461), .Q(i4[2]), .QN(n218)
         );
  DFNCND1 \i6_reg[3]  ( .D(n251), .CPN(Clk), .CDN(n4), .Q(i6[3]), .QN(n212) );
  DFNCND1 \i6_reg[1]  ( .D(n247), .CPN(Clk), .CDN(n4), .Q(i6[1]), .QN(n208) );
  DFNCND1 \i6_reg[2]  ( .D(n245), .CPN(Clk), .CDN(n4), .Q(i6[2]), .QN(n206) );
  DFCNQD1 TRes1_reg ( .D(n258), .CP(Clk), .CDN(n460), .Q(TRes1) );
  DFCNQD1 TDone1_reg ( .D(n257), .CP(Clk), .CDN(n461), .Q(TDone1) );
  DFCNQD1 TRes5_reg ( .D(n254), .CP(Clk), .CDN(n461), .Q(TRes5) );
  DFNCND1 \i4_reg[0]  ( .D(n268), .CPN(Clk), .CDN(n461), .Q(i4[0]), .QN(n222)
         );
  DFNCND1 \i6_reg[0]  ( .D(n249), .CPN(Clk), .CDN(n4), .Q(i6[0]), .QN(n210) );
  EDFCNQD1 \i3_reg[1]  ( .D(N320), .E(N326), .CP(Clk), .CDN(n461), .Q(i3[1])
         );
  EDFCNQD1 \i3_reg[2]  ( .D(N321), .E(N326), .CP(Clk), .CDN(n461), .Q(i3[2])
         );
  EDFCNQD1 \i3_reg[3]  ( .D(N322), .E(N326), .CP(Clk), .CDN(n461), .Q(i3[3])
         );
  EDFCNQD1 \i5_reg[1]  ( .D(N405), .E(N411), .CP(Clk), .CDN(n461), .Q(i5[1])
         );
  EDFCNQD1 \i5_reg[2]  ( .D(N406), .E(N411), .CP(Clk), .CDN(n461), .Q(i5[2])
         );
  EDFCNQD1 \i5_reg[3]  ( .D(N407), .E(N411), .CP(Clk), .CDN(n461), .Q(i5[3])
         );
  EDFCNQD1 \i3_reg[0]  ( .D(N319), .E(N326), .CP(Clk), .CDN(n35), .Q(i3[0]) );
  EDFCNQD1 \i5_reg[0]  ( .D(N404), .E(N411), .CP(Clk), .CDN(n461), .Q(i5[0])
         );
  EDFCNQD1 AllDoner_reg ( .D(N206), .E(N205), .CP(Clk), .CDN(n4), .Q(AllDoner)
         );
  DFCNQD1 TRes3_reg ( .D(n256), .CP(Clk), .CDN(n461), .Q(TRes3) );
  DFNCND1 \i2_reg[2]  ( .D(n277), .CPN(Clk), .CDN(n461), .Q(i2[2]), .QN(n230)
         );
  DFNCND1 \i2_reg[1]  ( .D(n279), .CPN(Clk), .CDN(n461), .Q(i2[1]), .QN(n232)
         );
  EDFCNQD1 \i1_reg[4]  ( .D(N230), .E(N233), .CP(Clk), .CDN(n461), .Q(i1[4])
         );
  DFNCND1 \i2_reg[4]  ( .D(n275), .CPN(Clk), .CDN(n461), .Q(i2[4]), .QN(n228)
         );
  EDFCNQD1 \i1_reg[1]  ( .D(N227), .E(N233), .CP(Clk), .CDN(n35), .Q(i1[1]) );
  EDFCNQD1 \i1_reg[2]  ( .D(N228), .E(N233), .CP(Clk), .CDN(n35), .Q(i1[2]) );
  EDFCNQD1 \i1_reg[3]  ( .D(N229), .E(N233), .CP(Clk), .CDN(n35), .Q(i1[3]) );
  EDFCNQD1 \i1_reg[0]  ( .D(N226), .E(N233), .CP(Clk), .CDN(n35), .Q(i1[0]) );
  DFNCND1 \i2_reg[0]  ( .D(n281), .CPN(Clk), .CDN(n461), .Q(i2[0]), .QN(n234)
         );
  EDFCNQD1 \State_reg[1]  ( .D(N216), .E(N217), .CP(Clk), .CDN(n461), .Q(
        State[1]) );
  EDFCNQD1 \State_reg[2]  ( .D(N218), .E(N217), .CP(Clk), .CDN(n460), .Q(
        State[2]) );
  EDFCNQD1 \State_reg[0]  ( .D(N214), .E(N217), .CP(Clk), .CDN(n460), .Q(
        State[0]) );
  EDFQD1 \DataO1_reg[27]  ( .D(i1[3]), .E(n1), .CP(Clk), .Q(DataO1[27]) );
  EDFQD1 \DataO1_reg[25]  ( .D(i1[1]), .E(n1), .CP(Clk), .Q(DataO1[25]) );
  EDFQD1 \DataO1_reg[19]  ( .D(i1[3]), .E(n1), .CP(Clk), .Q(DataO1[19]) );
  EDFQD1 \DataO1_reg[17]  ( .D(i1[1]), .E(n1), .CP(Clk), .Q(DataO1[17]) );
  EDFQD1 \DataO1_reg[11]  ( .D(i1[3]), .E(n1), .CP(Clk), .Q(DataO1[11]) );
  EDFQD1 \DataO1_reg[10]  ( .D(i1[2]), .E(n1), .CP(Clk), .Q(DataO1[10]) );
  EDFQD1 \DataO1_reg[12]  ( .D(i1[4]), .E(n1), .CP(Clk), .Q(DataO1[12]) );
  EDFQD1 \DataO1_reg[16]  ( .D(i1[0]), .E(n1), .CP(Clk), .Q(DataO1[16]) );
  EDFQD1 \DataO1_reg[18]  ( .D(i1[2]), .E(n1), .CP(Clk), .Q(DataO1[18]) );
  EDFQD1 \DataO1_reg[20]  ( .D(i1[4]), .E(n1), .CP(Clk), .Q(DataO1[20]) );
  EDFQD1 \DataO1_reg[24]  ( .D(i1[0]), .E(n1), .CP(Clk), .Q(DataO1[24]) );
  EDFQD1 \DataO1_reg[26]  ( .D(i1[2]), .E(n1), .CP(Clk), .Q(DataO1[26]) );
  EDFQD1 \DataO1_reg[28]  ( .D(i1[4]), .E(n1), .CP(Clk), .Q(DataO1[28]) );
  EDFQD1 \Addr1_reg[4]  ( .D(i1[4]), .E(n1), .CP(Clk), .Q(Addr1[4]) );
  EDFQD1 \Addr1_reg[2]  ( .D(i1[2]), .E(n1), .CP(Clk), .Q(Addr1[2]) );
  EDFQD1 \Addr1_reg[0]  ( .D(i1[0]), .E(n1), .CP(Clk), .Q(Addr1[0]) );
  EDFQD1 \Addr1_reg[1]  ( .D(i1[1]), .E(n1), .CP(Clk), .Q(Addr1[1]) );
  EDFQD1 \Addr1_reg[3]  ( .D(i1[3]), .E(n1), .CP(Clk), .Q(Addr1[3]) );
  EDFQD1 \Addr5_reg[4]  ( .D(i5[4]), .E(N449), .CP(Clk), .Q(Addr5[4]) );
  EDFQD1 \Addr5_reg[2]  ( .D(i5[2]), .E(N449), .CP(Clk), .Q(Addr5[2]) );
  EDFQD1 \Addr5_reg[0]  ( .D(i5[0]), .E(N449), .CP(Clk), .Q(Addr5[0]) );
  EDFQD1 \Addr5_reg[1]  ( .D(i5[1]), .E(N449), .CP(Clk), .Q(Addr5[1]) );
  EDFQD1 \Addr5_reg[3]  ( .D(i5[3]), .E(N449), .CP(Clk), .Q(Addr5[3]) );
  EDFQD1 \Addr3_reg[4]  ( .D(i3[4]), .E(N364), .CP(Clk), .Q(Addr3[4]) );
  EDFQD1 \Addr3_reg[2]  ( .D(i3[2]), .E(N364), .CP(Clk), .Q(Addr3[2]) );
  EDFQD1 \Addr3_reg[0]  ( .D(i3[0]), .E(N364), .CP(Clk), .Q(Addr3[0]) );
  EDFQD1 \Addr3_reg[1]  ( .D(i3[1]), .E(N364), .CP(Clk), .Q(Addr3[1]) );
  EDFQD1 \Addr3_reg[3]  ( .D(i3[3]), .E(N364), .CP(Clk), .Q(Addr3[3]) );
  DFNCND1 \i2_reg[3]  ( .D(n283), .CPN(Clk), .CDN(n461), .Q(i2[3]), .QN(n237)
         );
  DFNCND1 TRes6_reg ( .D(n241), .CPN(Clk), .CDN(n4), .QN(n202) );
  DFNCND1 TDone6_reg ( .D(n284), .CPN(Clk), .CDN(n4), .QN(n239) );
  DFNCND1 TDone4_reg ( .D(n259), .CPN(Clk), .CDN(n4), .QN(n213) );
  DFNCND1 TDone2_reg ( .D(n240), .CPN(Clk), .CDN(n461), .QN(n201) );
  DFNCND1 TRes2_reg ( .D(n272), .CPN(Clk), .CDN(n461), .QN(n226) );
  EDFCNQD1 \TestNo_reg[0]  ( .D(N208), .E(N211), .CP(Clk), .CDN(n460), .Q(
        TestNo[0]) );
  DFNCND1 TRes4_reg ( .D(n260), .CPN(Clk), .CDN(n4), .QN(n214) );
  EDFCNQD1 \TestNo_reg[2]  ( .D(N212), .E(N211), .CP(Clk), .CDN(n4), .Q(
        TestNo[2]) );
  EDFCNQD1 \TestNo_reg[1]  ( .D(N210), .E(N211), .CP(Clk), .CDN(n4), .Q(
        TestNo[1]) );
  EDFCNQD1 Testingr_reg ( .D(N204), .E(N203), .CP(Clk), .CDN(n4), .Q(Testing)
         );
  BUFFD1 U3 ( .I(n71), .Z(n306) );
  NR4D0 U4 ( .A1(N280), .A2(N279), .A3(N282), .A4(N281), .ZN(n71) );
  NR2D2 U5 ( .A1(n457), .A2(n127), .ZN(n1) );
  CKBXD0 U7 ( .I(n458), .Z(n5) );
  ND3D1 U8 ( .A1(TestNo[1]), .A2(n285), .A3(n126), .ZN(n2) );
  MUX3ND0 U10 ( .I0(n440), .I1(n455), .I2(n454), .S0(State[2]), .S1(State[1]), 
        .ZN(n3) );
  CKBD0 U12 ( .CLK(n285), .C(n458) );
  INVD0 U14 ( .I(n457), .ZN(n285) );
  BUFFD0 U16 ( .I(Reset), .Z(n457) );
  BUFFD0 U17 ( .I(n460), .Z(n4) );
  BUFFD0 U18 ( .I(n461), .Z(n6) );
  BUFFD0 U19 ( .I(n6), .Z(n7) );
  BUFFD0 U20 ( .I(n7), .Z(n8) );
  BUFFD0 U21 ( .I(n8), .Z(n9) );
  BUFFD0 U22 ( .I(n9), .Z(n10) );
  BUFFD0 U23 ( .I(n10), .Z(n11) );
  BUFFD0 U24 ( .I(n11), .Z(n12) );
  BUFFD0 U25 ( .I(n12), .Z(n13) );
  BUFFD0 U26 ( .I(n13), .Z(n14) );
  BUFFD0 U27 ( .I(n14), .Z(n15) );
  BUFFD0 U28 ( .I(n15), .Z(n16) );
  BUFFD0 U29 ( .I(n16), .Z(n17) );
  BUFFD0 U30 ( .I(n17), .Z(n18) );
  BUFFD0 U31 ( .I(n18), .Z(n19) );
  BUFFD0 U32 ( .I(n19), .Z(n20) );
  BUFFD0 U33 ( .I(n20), .Z(n21) );
  BUFFD0 U34 ( .I(n21), .Z(n22) );
  BUFFD0 U35 ( .I(n22), .Z(n23) );
  BUFFD0 U36 ( .I(n23), .Z(n24) );
  BUFFD0 U37 ( .I(n24), .Z(n25) );
  BUFFD0 U38 ( .I(n25), .Z(n26) );
  BUFFD0 U39 ( .I(n26), .Z(n27) );
  BUFFD0 U40 ( .I(n27), .Z(n28) );
  BUFFD0 U41 ( .I(n28), .Z(n29) );
  BUFFD0 U42 ( .I(n29), .Z(n30) );
  BUFFD0 U43 ( .I(n30), .Z(n31) );
  BUFFD0 U44 ( .I(n31), .Z(n32) );
  BUFFD0 U45 ( .I(n32), .Z(n33) );
  BUFFD0 U46 ( .I(n33), .Z(n34) );
  BUFFD0 U48 ( .I(n4), .Z(n35) );
  CKND2D0 U49 ( .A1(n113), .A2(n114), .ZN(n74) );
  BUFFD0 U50 ( .I(n37), .Z(n36) );
  BUFFD0 U54 ( .I(n38), .Z(n37) );
  BUFFD0 U57 ( .I(n40), .Z(n38) );
  BUFFD0 U58 ( .I(n74), .Z(n39) );
  BUFFD0 U60 ( .I(n41), .Z(n40) );
  BUFFD0 U61 ( .I(n42), .Z(n41) );
  BUFFD0 U63 ( .I(n43), .Z(n42) );
  BUFFD0 U65 ( .I(n44), .Z(n43) );
  BUFFD0 U67 ( .I(n45), .Z(n44) );
  BUFFD0 U69 ( .I(n46), .Z(n45) );
  BUFFD0 U70 ( .I(n47), .Z(n46) );
  BUFFD0 U71 ( .I(n48), .Z(n47) );
  BUFFD0 U73 ( .I(n49), .Z(n48) );
  BUFFD0 U74 ( .I(n50), .Z(n49) );
  BUFFD0 U75 ( .I(n51), .Z(n50) );
  BUFFD0 U76 ( .I(n52), .Z(n51) );
  BUFFD0 U77 ( .I(n53), .Z(n52) );
  BUFFD0 U78 ( .I(n54), .Z(n53) );
  BUFFD0 U79 ( .I(n55), .Z(n54) );
  BUFFD0 U80 ( .I(n56), .Z(n55) );
  BUFFD0 U81 ( .I(n57), .Z(n56) );
  BUFFD0 U82 ( .I(n58), .Z(n57) );
  BUFFD0 U83 ( .I(n59), .Z(n58) );
  BUFFD0 U84 ( .I(n60), .Z(n59) );
  BUFFD0 U85 ( .I(n61), .Z(n60) );
  BUFFD0 U86 ( .I(n62), .Z(n61) );
  BUFFD0 U87 ( .I(n63), .Z(n62) );
  BUFFD0 U88 ( .I(n64), .Z(n63) );
  BUFFD0 U89 ( .I(n65), .Z(n64) );
  BUFFD0 U91 ( .I(n66), .Z(n65) );
  BUFFD0 U92 ( .I(n67), .Z(n66) );
  BUFFD0 U93 ( .I(n68), .Z(n67) );
  BUFFD0 U94 ( .I(n175), .Z(n68) );
  BUFFD0 U96 ( .I(n182), .Z(n175) );
  BUFFD0 U98 ( .I(n225), .Z(n182) );
  BUFFD0 U100 ( .I(n236), .Z(n225) );
  BUFFD0 U102 ( .I(n238), .Z(n236) );
  BUFFD0 U103 ( .I(n286), .Z(n238) );
  BUFFD0 U104 ( .I(n287), .Z(n286) );
  BUFFD0 U106 ( .I(n288), .Z(n287) );
  BUFFD0 U107 ( .I(n289), .Z(n288) );
  BUFFD0 U108 ( .I(n290), .Z(n289) );
  BUFFD0 U109 ( .I(n291), .Z(n290) );
  BUFFD0 U110 ( .I(n292), .Z(n291) );
  BUFFD0 U111 ( .I(n293), .Z(n292) );
  BUFFD0 U112 ( .I(n294), .Z(n293) );
  BUFFD0 U113 ( .I(n295), .Z(n294) );
  BUFFD0 U114 ( .I(n296), .Z(n295) );
  BUFFD0 U115 ( .I(n297), .Z(n296) );
  BUFFD0 U116 ( .I(n298), .Z(n297) );
  BUFFD0 U117 ( .I(n299), .Z(n298) );
  BUFFD0 U122 ( .I(n300), .Z(n299) );
  BUFFD0 U127 ( .I(n301), .Z(n300) );
  BUFFD0 U128 ( .I(n302), .Z(n301) );
  BUFFD0 U129 ( .I(n303), .Z(n302) );
  BUFFD0 U130 ( .I(n304), .Z(n303) );
  BUFFD0 U131 ( .I(n39), .Z(n304) );
  OAI21D0 U132 ( .A1(n111), .A2(n75), .B(n239), .ZN(n284) );
  OAI21D0 U133 ( .A1(n69), .A2(n70), .B(n201), .ZN(n240) );
  BUFFD0 U134 ( .I(n307), .Z(n305) );
  BUFFD0 U135 ( .I(n308), .Z(n307) );
  BUFFD0 U136 ( .I(n309), .Z(n308) );
  BUFFD0 U138 ( .I(n310), .Z(n309) );
  BUFFD0 U139 ( .I(n311), .Z(n310) );
  BUFFD0 U140 ( .I(n312), .Z(n311) );
  BUFFD0 U141 ( .I(n313), .Z(n312) );
  BUFFD0 U142 ( .I(n314), .Z(n313) );
  BUFFD0 U143 ( .I(n315), .Z(n314) );
  BUFFD0 U145 ( .I(n316), .Z(n315) );
  BUFFD0 U146 ( .I(n317), .Z(n316) );
  BUFFD0 U147 ( .I(n318), .Z(n317) );
  BUFFD0 U148 ( .I(n319), .Z(n318) );
  BUFFD0 U149 ( .I(n320), .Z(n319) );
  BUFFD0 U150 ( .I(n321), .Z(n320) );
  BUFFD0 U151 ( .I(n322), .Z(n321) );
  BUFFD0 U152 ( .I(n323), .Z(n322) );
  BUFFD0 U153 ( .I(n324), .Z(n323) );
  BUFFD0 U154 ( .I(n325), .Z(n324) );
  BUFFD0 U155 ( .I(n326), .Z(n325) );
  BUFFD0 U156 ( .I(n327), .Z(n326) );
  BUFFD0 U157 ( .I(n328), .Z(n327) );
  BUFFD0 U158 ( .I(n329), .Z(n328) );
  BUFFD0 U159 ( .I(n330), .Z(n329) );
  BUFFD0 U160 ( .I(n331), .Z(n330) );
  BUFFD0 U161 ( .I(n332), .Z(n331) );
  BUFFD0 U162 ( .I(n333), .Z(n332) );
  BUFFD0 U164 ( .I(n334), .Z(n333) );
  BUFFD0 U165 ( .I(n335), .Z(n334) );
  BUFFD0 U166 ( .I(n336), .Z(n335) );
  BUFFD0 U167 ( .I(n337), .Z(n336) );
  BUFFD0 U168 ( .I(n338), .Z(n337) );
  BUFFD0 U169 ( .I(n339), .Z(n338) );
  BUFFD0 U170 ( .I(n340), .Z(n339) );
  BUFFD0 U171 ( .I(n341), .Z(n340) );
  BUFFD0 U172 ( .I(n342), .Z(n341) );
  BUFFD0 U173 ( .I(n343), .Z(n342) );
  BUFFD0 U174 ( .I(n344), .Z(n343) );
  BUFFD0 U175 ( .I(n345), .Z(n344) );
  BUFFD0 U176 ( .I(n346), .Z(n345) );
  BUFFD0 U177 ( .I(n347), .Z(n346) );
  BUFFD0 U178 ( .I(n348), .Z(n347) );
  BUFFD0 U179 ( .I(n349), .Z(n348) );
  BUFFD0 U180 ( .I(n350), .Z(n349) );
  BUFFD0 U181 ( .I(n351), .Z(n350) );
  BUFFD0 U182 ( .I(n352), .Z(n351) );
  BUFFD0 U183 ( .I(n353), .Z(n352) );
  BUFFD0 U184 ( .I(n354), .Z(n353) );
  BUFFD0 U185 ( .I(n355), .Z(n354) );
  BUFFD0 U186 ( .I(n356), .Z(n355) );
  BUFFD0 U187 ( .I(n357), .Z(n356) );
  BUFFD0 U189 ( .I(n358), .Z(n357) );
  BUFFD0 U190 ( .I(n359), .Z(n358) );
  BUFFD0 U191 ( .I(n360), .Z(n359) );
  BUFFD0 U192 ( .I(n361), .Z(n360) );
  BUFFD0 U193 ( .I(n362), .Z(n361) );
  BUFFD0 U194 ( .I(n306), .Z(n362) );
  BUFFD0 U195 ( .I(n364), .Z(n363) );
  BUFFD0 U196 ( .I(n365), .Z(n364) );
  BUFFD0 U197 ( .I(n366), .Z(n365) );
  BUFFD0 U198 ( .I(n367), .Z(n366) );
  BUFFD0 U199 ( .I(n368), .Z(n367) );
  BUFFD0 U200 ( .I(n369), .Z(n368) );
  BUFFD0 U201 ( .I(n370), .Z(n369) );
  BUFFD0 U202 ( .I(n371), .Z(n370) );
  BUFFD0 U203 ( .I(n372), .Z(n371) );
  BUFFD0 U204 ( .I(n373), .Z(n372) );
  BUFFD0 U205 ( .I(n374), .Z(n373) );
  BUFFD0 U206 ( .I(n375), .Z(n374) );
  BUFFD0 U207 ( .I(n376), .Z(n375) );
  BUFFD0 U208 ( .I(n377), .Z(n376) );
  BUFFD0 U209 ( .I(n378), .Z(n377) );
  BUFFD0 U210 ( .I(n379), .Z(n378) );
  BUFFD0 U211 ( .I(n380), .Z(n379) );
  BUFFD0 U212 ( .I(n381), .Z(n380) );
  BUFFD0 U213 ( .I(n382), .Z(n381) );
  BUFFD0 U214 ( .I(n383), .Z(n382) );
  BUFFD0 U215 ( .I(n384), .Z(n383) );
  BUFFD0 U216 ( .I(n385), .Z(n384) );
  BUFFD0 U217 ( .I(n386), .Z(n385) );
  BUFFD0 U218 ( .I(n387), .Z(n386) );
  BUFFD0 U219 ( .I(n388), .Z(n387) );
  BUFFD0 U220 ( .I(n389), .Z(n388) );
  BUFFD0 U221 ( .I(n390), .Z(n389) );
  BUFFD0 U222 ( .I(n391), .Z(n390) );
  BUFFD0 U223 ( .I(n392), .Z(n391) );
  BUFFD0 U224 ( .I(n393), .Z(n392) );
  BUFFD0 U225 ( .I(n394), .Z(n393) );
  BUFFD0 U226 ( .I(n395), .Z(n394) );
  BUFFD0 U227 ( .I(n396), .Z(n395) );
  BUFFD0 U228 ( .I(n397), .Z(n396) );
  BUFFD0 U229 ( .I(n398), .Z(n397) );
  BUFFD0 U230 ( .I(n399), .Z(n398) );
  BUFFD0 U231 ( .I(n400), .Z(n399) );
  BUFFD0 U232 ( .I(n401), .Z(n400) );
  BUFFD0 U233 ( .I(n402), .Z(n401) );
  BUFFD0 U234 ( .I(n403), .Z(n402) );
  BUFFD0 U235 ( .I(n404), .Z(n403) );
  BUFFD0 U236 ( .I(n405), .Z(n404) );
  BUFFD0 U237 ( .I(n406), .Z(n405) );
  BUFFD0 U238 ( .I(n407), .Z(n406) );
  BUFFD0 U239 ( .I(n408), .Z(n407) );
  BUFFD0 U240 ( .I(n409), .Z(n408) );
  BUFFD0 U241 ( .I(n410), .Z(n409) );
  BUFFD0 U242 ( .I(n411), .Z(n410) );
  BUFFD0 U243 ( .I(n412), .Z(n411) );
  BUFFD0 U244 ( .I(n413), .Z(n412) );
  BUFFD0 U245 ( .I(n414), .Z(n413) );
  BUFFD0 U246 ( .I(n415), .Z(n414) );
  BUFFD0 U247 ( .I(n416), .Z(n415) );
  BUFFD0 U248 ( .I(n417), .Z(n416) );
  BUFFD0 U249 ( .I(n418), .Z(n417) );
  BUFFD0 U250 ( .I(n419), .Z(n418) );
  BUFFD0 U251 ( .I(n420), .Z(n419) );
  BUFFD0 U252 ( .I(n84), .Z(n420) );
  CKBD0 U253 ( .CLK(n456), .C(n421) );
  CKNXD16 U254 ( .I(n421), .ZN(TestOK) );
  AO211D0 U255 ( .A1(N172), .A2(n134), .B(ParityErr), .C(n174), .Z(N205) );
  NR2D0 U256 ( .A1(n158), .A2(Testing), .ZN(N204) );
  CKAN2D0 U257 ( .A1(n169), .A2(Testing), .Z(N186) );
  NR2D0 U258 ( .A1(n179), .A2(n464), .ZN(N185) );
  NR2D0 U259 ( .A1(n464), .A2(n158), .ZN(n134) );
  INVD1 U260 ( .I(n88), .ZN(n87) );
  BUFFD1 U261 ( .I(n34), .Z(n460) );
  BUFFD1 U262 ( .I(n458), .Z(n461) );
  ND2D1 U263 ( .A1(n89), .A2(n35), .ZN(n88) );
  INVD1 U264 ( .I(n77), .ZN(n76) );
  INVD1 U265 ( .I(n109), .ZN(n108) );
  BUFFD1 U266 ( .I(n285), .Z(n459) );
  INR2D1 U267 ( .A1(n307), .B1(n70), .ZN(n104) );
  ND2D1 U268 ( .A1(n78), .A2(n35), .ZN(n77) );
  ND2D1 U269 ( .A1(n105), .A2(n35), .ZN(n109) );
  INVD1 U270 ( .I(n102), .ZN(n89) );
  INVD1 U271 ( .I(n2), .ZN(DataO[31]) );
  INVD1 U272 ( .I(n134), .ZN(n138) );
  INVD1 U273 ( .I(n152), .ZN(n140) );
  INVD1 U274 ( .I(n164), .ZN(N145) );
  INVD1 U275 ( .I(n155), .ZN(N158) );
  NR2D1 U276 ( .A1(n40), .A2(n75), .ZN(n73) );
  NR2D1 U277 ( .A1(n83), .A2(n363), .ZN(n86) );
  OAI21D1 U278 ( .A1(n78), .A2(n79), .B(n80), .ZN(n252) );
  INVD1 U279 ( .I(n73), .ZN(n80) );
  OAI21D1 U280 ( .A1(n105), .A2(n106), .B(n107), .ZN(n273) );
  INVD1 U281 ( .I(n104), .ZN(n107) );
  OAI21D1 U282 ( .A1(n89), .A2(n90), .B(n91), .ZN(n271) );
  INVD1 U283 ( .I(n86), .ZN(n91) );
  ND2D1 U284 ( .A1(n124), .A2(n199), .ZN(n102) );
  ND2D1 U285 ( .A1(n105), .A2(n106), .ZN(n70) );
  ND2D1 U286 ( .A1(n78), .A2(n79), .ZN(n75) );
  ND2D1 U287 ( .A1(n89), .A2(n90), .ZN(n83) );
  INVD1 U288 ( .I(n112), .ZN(n78) );
  INVD1 U289 ( .I(n110), .ZN(n105) );
  INVD1 U290 ( .I(n154), .ZN(N165) );
  NR2D1 U291 ( .A1(n153), .A2(n138), .ZN(N212) );
  AOI222D0 U292 ( .A1(n140), .A2(n154), .B1(n143), .B2(n155), .C1(n141), .C2(
        n156), .ZN(n153) );
  NR2D1 U293 ( .A1(n161), .A2(n138), .ZN(N210) );
  AOI222D0 U294 ( .A1(n162), .A2(n163), .B1(n139), .B2(n164), .C1(n140), .C2(
        n154), .ZN(n161) );
  INVD1 U295 ( .I(n163), .ZN(N138) );
  INVD1 U296 ( .I(n156), .ZN(N151) );
  INVD1 U297 ( .I(n141), .ZN(n180) );
  INVD1 U298 ( .I(n463), .ZN(n462) );
  INVD1 U299 ( .I(N221), .ZN(n158) );
  OAI21D1 U300 ( .A1(n157), .A2(n158), .B(n146), .ZN(N211) );
  NR2D1 U301 ( .A1(n159), .A2(n160), .ZN(n157) );
  OAI21D1 U302 ( .A1(n170), .A2(n158), .B(n135), .ZN(N206) );
  NR2D1 U303 ( .A1(n132), .A2(n160), .ZN(n170) );
  NR2D1 U304 ( .A1(n174), .A2(N204), .ZN(n146) );
  OAI222D0 U305 ( .A1(TestDone[5]), .A2(n168), .B1(TestDone[1]), .B2(n171), 
        .C1(TestDone[3]), .C2(n173), .ZN(n169) );
  INVD1 U306 ( .I(n125), .ZN(N326) );
  INVD1 U307 ( .I(n123), .ZN(N411) );
  INVD1 U308 ( .I(n127), .ZN(N233) );
  NR2D1 U309 ( .A1(n457), .A2(n125), .ZN(N364) );
  NR2D1 U310 ( .A1(n457), .A2(n123), .ZN(N449) );
  INVD1 U311 ( .I(n143), .ZN(n168) );
  NR2D1 U312 ( .A1(n178), .A2(n176), .ZN(n132) );
  ND2D1 U313 ( .A1(n132), .A2(n159), .ZN(n152) );
  ND4D1 U314 ( .A1(n171), .A2(n168), .A3(n172), .A4(n173), .ZN(n160) );
  NR2D1 U315 ( .A1(n162), .A2(n141), .ZN(n172) );
  INVD1 U316 ( .I(n142), .ZN(n171) );
  INVD1 U317 ( .I(n139), .ZN(n173) );
  INVD1 U318 ( .I(n162), .ZN(n145) );
  NR2D1 U319 ( .A1(n167), .A2(n177), .ZN(N132) );
  INVD1 U320 ( .I(n131), .ZN(n167) );
  ND2D1 U321 ( .A1(TestDone[5]), .A2(n130), .ZN(n155) );
  ND2D1 U322 ( .A1(TestDone[3]), .A2(n81), .ZN(n164) );
  INVD1 U323 ( .I(n177), .ZN(TestDone[1]) );
  AN3D1 U324 ( .A1(n151), .A2(n152), .A3(n145), .Z(n147) );
  OAI21D1 U325 ( .A1(n457), .A2(n81), .B(n139), .ZN(n151) );
  IOA21D1 U326 ( .A1(N326), .A2(N324), .B(n81), .ZN(n256) );
  INVD1 U327 ( .I(Testing), .ZN(n464) );
  NR4D0 U328 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(n113) );
  NR4D0 U329 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(n114) );
  ND2D1 U330 ( .A1(n92), .A2(n93), .ZN(n84) );
  NR4D0 U331 ( .A1(n98), .A2(n99), .A3(n100), .A4(n101), .ZN(n92) );
  NR4D0 U332 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(n93) );
  ND4D1 U333 ( .A1(DataI[27]), .A2(DataI[26]), .A3(DataI[25]), .A4(DataI[24]), 
        .ZN(n98) );
  NR2D1 U334 ( .A1(n305), .A2(n70), .ZN(n103) );
  INR2D1 U335 ( .A1(n36), .B1(n75), .ZN(n72) );
  INR2D1 U336 ( .A1(n363), .B1(n83), .ZN(n85) );
  ND4D1 U337 ( .A1(DataI[1]), .A2(DataI[19]), .A3(DataI[18]), .A4(DataI[17]), 
        .ZN(n96) );
  ND4D1 U338 ( .A1(DataI[9]), .A2(DataI[8]), .A3(DataI[7]), .A4(DataI[6]), 
        .ZN(n101) );
  ND4D1 U339 ( .A1(DataI[30]), .A2(DataI[2]), .A3(DataI[29]), .A4(DataI[28]), 
        .ZN(n99) );
  ND4D1 U340 ( .A1(DataI[12]), .A2(DataI[11]), .A3(DataI[10]), .A4(DataI[0]), 
        .ZN(n94) );
  ND4D1 U341 ( .A1(DataI[16]), .A2(DataI[15]), .A3(DataI[14]), .A4(DataI[13]), 
        .ZN(n95) );
  ND4D1 U342 ( .A1(DataI[5]), .A2(DataI[4]), .A3(DataI[3]), .A4(DataI[31]), 
        .ZN(n100) );
  ND4D1 U343 ( .A1(DataI[23]), .A2(DataI[22]), .A3(DataI[21]), .A4(DataI[20]), 
        .ZN(n97) );
  INR2D1 U344 ( .A1(n305), .B1(N289), .ZN(n69) );
  NR2D1 U345 ( .A1(N460), .A2(n36), .ZN(n111) );
  OAI21D1 U346 ( .A1(n82), .A2(n83), .B(n213), .ZN(n259) );
  NR2D1 U347 ( .A1(N375), .A2(n363), .ZN(n82) );
  ND2D1 U348 ( .A1(n196), .A2(n197), .ZN(Addr[0]) );
  AOI22D0 U349 ( .A1(Addr3[0]), .A2(DataO[31]), .B1(Addr5[0]), .B2(n186), .ZN(
        n196) );
  AOI22D0 U350 ( .A1(n198), .A2(n458), .B1(Addr1[0]), .B2(n462), .ZN(n197) );
  OAI222D0 U351 ( .A1(n209), .A2(n112), .B1(n221), .B2(n102), .C1(n233), .C2(
        n110), .ZN(n198) );
  ND2D1 U352 ( .A1(n193), .A2(n194), .ZN(Addr[1]) );
  AOI22D0 U353 ( .A1(Addr3[1]), .A2(DataO[31]), .B1(Addr5[1]), .B2(n186), .ZN(
        n193) );
  AOI22D0 U354 ( .A1(n195), .A2(n458), .B1(Addr1[1]), .B2(n462), .ZN(n194) );
  OAI222D0 U355 ( .A1(n207), .A2(n112), .B1(n219), .B2(n102), .C1(n231), .C2(
        n110), .ZN(n195) );
  ND2D1 U356 ( .A1(n190), .A2(n191), .ZN(Addr[2]) );
  AOI22D0 U357 ( .A1(Addr3[2]), .A2(DataO[31]), .B1(Addr5[2]), .B2(n186), .ZN(
        n190) );
  AOI22D0 U358 ( .A1(n192), .A2(n5), .B1(Addr1[2]), .B2(n462), .ZN(n191) );
  OAI222D0 U359 ( .A1(n205), .A2(n112), .B1(n217), .B2(n102), .C1(n229), .C2(
        n110), .ZN(n192) );
  ND2D1 U360 ( .A1(n187), .A2(n188), .ZN(Addr[3]) );
  AOI22D0 U361 ( .A1(Addr3[3]), .A2(DataO[31]), .B1(Addr5[3]), .B2(n186), .ZN(
        n187) );
  AOI22D0 U362 ( .A1(n189), .A2(n458), .B1(Addr1[3]), .B2(n462), .ZN(n188) );
  OAI222D0 U363 ( .A1(n211), .A2(n112), .B1(n223), .B2(n102), .C1(n235), .C2(
        n110), .ZN(n189) );
  ND2D1 U364 ( .A1(n183), .A2(n184), .ZN(Addr[4]) );
  AOI22D0 U365 ( .A1(Addr3[4]), .A2(DataO[31]), .B1(Addr5[4]), .B2(n186), .ZN(
        n183) );
  AOI22D0 U366 ( .A1(n185), .A2(n6), .B1(Addr1[4]), .B2(n462), .ZN(n184) );
  OAI222D0 U367 ( .A1(n203), .A2(n112), .B1(n215), .B2(n102), .C1(n227), .C2(
        n110), .ZN(n185) );
  AN2D1 U368 ( .A1(TestDone[6]), .A2(n159), .Z(n447) );
  ND3D1 U369 ( .A1(TestNo[1]), .A2(n199), .A3(TestNo[2]), .ZN(n112) );
  ND3D1 U370 ( .A1(n199), .A2(n200), .A3(TestNo[1]), .ZN(n110) );
  OAI22D0 U371 ( .A1(n203), .A2(n76), .B1(n204), .B2(n77), .ZN(n242) );
  OAI22D0 U372 ( .A1(n205), .A2(n76), .B1(n206), .B2(n77), .ZN(n244) );
  OAI22D0 U373 ( .A1(n207), .A2(n76), .B1(n208), .B2(n77), .ZN(n246) );
  OAI22D0 U374 ( .A1(n209), .A2(n76), .B1(n210), .B2(n77), .ZN(n248) );
  OAI22D0 U375 ( .A1(n211), .A2(n76), .B1(n212), .B2(n77), .ZN(n250) );
  OAI22D0 U376 ( .A1(n215), .A2(n87), .B1(n216), .B2(n88), .ZN(n261) );
  OAI22D0 U377 ( .A1(n217), .A2(n87), .B1(n218), .B2(n88), .ZN(n263) );
  OAI22D0 U378 ( .A1(n219), .A2(n87), .B1(n220), .B2(n88), .ZN(n265) );
  OAI22D0 U379 ( .A1(n221), .A2(n87), .B1(n222), .B2(n88), .ZN(n267) );
  OAI22D0 U380 ( .A1(n223), .A2(n87), .B1(n224), .B2(n88), .ZN(n269) );
  OAI22D0 U381 ( .A1(n227), .A2(n108), .B1(n228), .B2(n109), .ZN(n274) );
  OAI22D0 U382 ( .A1(n229), .A2(n108), .B1(n230), .B2(n109), .ZN(n276) );
  OAI22D0 U383 ( .A1(n231), .A2(n108), .B1(n232), .B2(n109), .ZN(n278) );
  OAI22D0 U384 ( .A1(n233), .A2(n108), .B1(n234), .B2(n109), .ZN(n280) );
  OAI22D0 U385 ( .A1(n235), .A2(n108), .B1(n237), .B2(n109), .ZN(n282) );
  INVD1 U386 ( .I(TestNo[0]), .ZN(n199) );
  IND3D1 U387 ( .A1(N184), .B1(n135), .B2(n146), .ZN(N203) );
  ND2D1 U388 ( .A1(State[0]), .A2(N132), .ZN(n444) );
  INR2D1 U389 ( .A1(State[0]), .B1(N132), .ZN(n441) );
  AO22D0 U390 ( .A1(n133), .A2(ParityErr), .B1(N170), .B2(n134), .Z(N219) );
  INVD1 U391 ( .I(n135), .ZN(n133) );
  INR2D1 U392 ( .A1(State[0]), .B1(N132), .ZN(n442) );
  AOI31D0 U393 ( .A1(n147), .A2(n148), .A3(n149), .B(n138), .ZN(N216) );
  NR2D1 U394 ( .A1(n143), .A2(n142), .ZN(n149) );
  OAI21D1 U395 ( .A1(n457), .A2(n214), .B(n141), .ZN(n148) );
  ND2D1 U396 ( .A1(n202), .A2(TestDone[6]), .ZN(n154) );
  NR2D1 U397 ( .A1(n200), .A2(TestNo[1]), .ZN(n124) );
  IOA21D1 U398 ( .A1(n3), .A2(N221), .B(n146), .ZN(N217) );
  INR2D1 U399 ( .A1(State[0]), .B1(TestDone[1]), .ZN(n440) );
  AOI21D1 U400 ( .A1(n136), .A2(n137), .B(n138), .ZN(N218) );
  NR3D0 U401 ( .A1(n139), .A2(n140), .A3(n141), .ZN(n137) );
  AOI211D1 U402 ( .A1(n142), .A2(n131), .B(n143), .C(n144), .ZN(n136) );
  NR2D1 U403 ( .A1(n457), .A2(n239), .ZN(TestDone[6]) );
  NR2D1 U404 ( .A1(n457), .A2(n201), .ZN(TestDone[2]) );
  NR2D1 U405 ( .A1(n457), .A2(n213), .ZN(TestDone[4]) );
  INVD1 U406 ( .I(TestNo[2]), .ZN(n200) );
  ND2D1 U407 ( .A1(n214), .A2(TestDone[4]), .ZN(n156) );
  ND2D1 U408 ( .A1(n226), .A2(TestDone[2]), .ZN(n163) );
  NR4D0 U409 ( .A1(n128), .A2(n129), .A3(n130), .A4(n131), .ZN(N220) );
  ND4D1 U410 ( .A1(TRes3), .A2(State[0]), .A3(N221), .A4(n132), .ZN(n128) );
  IOA21D1 U411 ( .A1(DataO1[24]), .A2(n462), .B(n2), .ZN(DataO[24]) );
  IOA21D1 U412 ( .A1(DataO1[25]), .A2(n462), .B(n2), .ZN(DataO[25]) );
  IOA21D1 U413 ( .A1(DataO1[26]), .A2(n462), .B(n2), .ZN(DataO[26]) );
  IOA21D1 U414 ( .A1(DataO1[27]), .A2(n181), .B(n2), .ZN(DataO[27]) );
  IOA21D1 U415 ( .A1(DataO1[28]), .A2(n462), .B(n2), .ZN(DataO[28]) );
  NR2D1 U416 ( .A1(n199), .A2(TestNo[2]), .ZN(n126) );
  INVD1 U417 ( .I(n181), .ZN(n463) );
  INR3D0 U418 ( .A1(n126), .B1(n457), .B2(TestNo[1]), .ZN(n181) );
  AN3D1 U419 ( .A1(n124), .A2(n459), .A3(TestNo[0]), .Z(n186) );
  IOA21D1 U420 ( .A1(DataO1[0]), .A2(n462), .B(n2), .ZN(DataO[0]) );
  IOA21D1 U421 ( .A1(DataO1[1]), .A2(n462), .B(n2), .ZN(DataO[1]) );
  IOA21D1 U422 ( .A1(DataO1[2]), .A2(n181), .B(n2), .ZN(DataO[2]) );
  IOA21D1 U423 ( .A1(DataO1[3]), .A2(n181), .B(n2), .ZN(DataO[3]) );
  IOA21D1 U424 ( .A1(DataO1[4]), .A2(n181), .B(n2), .ZN(DataO[4]) );
  IOA21D1 U425 ( .A1(DataO1[8]), .A2(n181), .B(n2), .ZN(DataO[8]) );
  IOA21D1 U426 ( .A1(DataO1[9]), .A2(n181), .B(n2), .ZN(DataO[9]) );
  IOA21D1 U427 ( .A1(DataO1[10]), .A2(n462), .B(n2), .ZN(DataO[10]) );
  IOA21D1 U428 ( .A1(DataO1[11]), .A2(n462), .B(n2), .ZN(DataO[11]) );
  IOA21D1 U429 ( .A1(DataO1[12]), .A2(n462), .B(n2), .ZN(DataO[12]) );
  IOA21D1 U430 ( .A1(DataO1[16]), .A2(n462), .B(n2), .ZN(DataO[16]) );
  IOA21D1 U431 ( .A1(DataO1[17]), .A2(n462), .B(n2), .ZN(DataO[17]) );
  IOA21D1 U432 ( .A1(DataO1[18]), .A2(n462), .B(n2), .ZN(DataO[18]) );
  IOA21D1 U433 ( .A1(DataO1[19]), .A2(n462), .B(n2), .ZN(DataO[19]) );
  IOA21D1 U434 ( .A1(DataO1[20]), .A2(n181), .B(n2), .ZN(DataO[20]) );
  OAI21D0 U435 ( .A1(ParityErr), .A2(AllDoner), .B(DoSelfTest), .ZN(n135) );
  NR3D0 U436 ( .A1(AllDoner), .A2(ParityErr), .A3(n174), .ZN(N221) );
  AOI31D0 U437 ( .A1(n147), .A2(State[0]), .A3(n150), .B(n138), .ZN(N214) );
  AOI22D0 U438 ( .A1(n142), .A2(n131), .B1(n143), .B2(n130), .ZN(n150) );
  AOI21D1 U439 ( .A1(n165), .A2(n166), .B(n138), .ZN(N208) );
  AOI22D0 U440 ( .A1(n139), .A2(TRes3), .B1(n142), .B2(n167), .ZN(n166) );
  NR3D0 U441 ( .A1(State[0]), .A2(State[1]), .A3(n178), .ZN(n141) );
  NR3D0 U442 ( .A1(State[1]), .A2(State[2]), .A3(n159), .ZN(n142) );
  NR3D0 U443 ( .A1(n178), .A2(State[1]), .A3(n159), .ZN(n143) );
  NR3D0 U444 ( .A1(n176), .A2(State[2]), .A3(n159), .ZN(n139) );
  INVD1 U445 ( .I(State[0]), .ZN(n159) );
  NR3D0 U446 ( .A1(State[0]), .A2(State[2]), .A3(n176), .ZN(n162) );
  INVD1 U447 ( .I(State[2]), .ZN(n178) );
  INVD1 U448 ( .I(State[1]), .ZN(n176) );
  ND2D1 U449 ( .A1(TRes1), .A2(n460), .ZN(n131) );
  INVD1 U450 ( .I(DoSelfTest), .ZN(n174) );
  ND2D1 U451 ( .A1(TRes5), .A2(n460), .ZN(n130) );
  ND2D1 U452 ( .A1(n126), .A2(TestNo[1]), .ZN(n125) );
  INVD1 U453 ( .I(TRes3), .ZN(n81) );
  ND2D1 U454 ( .A1(n124), .A2(TestNo[0]), .ZN(n123) );
  AN2D1 U455 ( .A1(TDone3), .A2(n458), .Z(TestDone[3]) );
  AN2D1 U456 ( .A1(TDone5), .A2(n458), .Z(TestDone[5]) );
  ND2D1 U457 ( .A1(TDone1), .A2(n460), .ZN(n177) );
  IND2D1 U458 ( .A1(TestNo[1]), .B1(n126), .ZN(n127) );
  BUFFD1 U459 ( .I(DataO[31]), .Z(DataO[30]) );
  BUFFD1 U460 ( .I(DataO[31]), .Z(DataO[29]) );
  BUFFD1 U461 ( .I(DataO[31]), .Z(DataO[23]) );
  BUFFD1 U462 ( .I(DataO[31]), .Z(DataO[22]) );
  BUFFD1 U463 ( .I(DataO[31]), .Z(DataO[21]) );
  BUFFD1 U464 ( .I(DataO[31]), .Z(DataO[15]) );
  BUFFD1 U465 ( .I(DataO[31]), .Z(DataO[14]) );
  BUFFD1 U466 ( .I(DataO[31]), .Z(DataO[13]) );
  BUFFD1 U467 ( .I(DataO[31]), .Z(DataO[7]) );
  BUFFD1 U468 ( .I(DataO[31]), .Z(DataO[6]) );
  BUFFD1 U469 ( .I(DataO[31]), .Z(DataO[5]) );
  OR2D1 U470 ( .A1(N165), .A2(State[0]), .Z(n443) );
  MUX3ND0 U471 ( .I0(n444), .I1(n445), .I2(n446), .S0(State[2]), .S1(State[1]), 
        .ZN(N184) );
  OR2D1 U472 ( .A1(N165), .A2(State[0]), .Z(n448) );
  MUX3ND0 U473 ( .I0(n441), .I1(n449), .I2(n450), .S0(State[2]), .S1(State[1]), 
        .ZN(N172) );
  OR2D1 U474 ( .A1(N165), .A2(State[0]), .Z(n451) );
  MUX3ND0 U475 ( .I0(n442), .I1(n452), .I2(n453), .S0(State[2]), .S1(State[1]), 
        .ZN(N170) );
  MUX3ND0 U476 ( .I0(N138), .I1(N145), .I2(n443), .S0(State[0]), .S1(State[2]), 
        .ZN(n446) );
  MUX2ND0 U477 ( .I0(N151), .I1(N158), .S(State[0]), .ZN(n445) );
  MUX3ND0 U478 ( .I0(TestDone[2]), .I1(TestDone[3]), .I2(n447), .S0(State[0]), 
        .S1(State[2]), .ZN(n454) );
  MUX2ND0 U479 ( .I0(TestDone[4]), .I1(TestDone[5]), .S(State[0]), .ZN(n455)
         );
  MUX3ND0 U480 ( .I0(N138), .I1(N145), .I2(n448), .S0(State[0]), .S1(State[2]), 
        .ZN(n450) );
  MUX2ND0 U481 ( .I0(N151), .I1(N158), .S(State[0]), .ZN(n449) );
  MUX3ND0 U482 ( .I0(N138), .I1(N145), .I2(n451), .S0(State[0]), .S1(State[2]), 
        .ZN(n453) );
  MUX2ND0 U483 ( .I0(N151), .I1(N158), .S(State[0]), .ZN(n452) );
  CKND0 U484 ( .CLK(n519), .CN(n456) );
  AN3D0 U485 ( .A1(N227), .A2(N226), .A3(N228), .Z(n465) );
  AN3D0 U486 ( .A1(N230), .A2(N229), .A3(n465), .Z(N231) );
  IND2D0 U487 ( .A1(i2[3]), .B1(DataI[27]), .ZN(n477) );
  CKND0 U488 ( .CLK(DataI[24]), .CN(n471) );
  IOA21D0 U489 ( .A1(n471), .A2(i2[0]), .B(DataI[25]), .ZN(n469) );
  INR2D0 U490 ( .A1(i2[2]), .B1(DataI[26]), .ZN(n468) );
  INR2D0 U491 ( .A1(i2[3]), .B1(DataI[27]), .ZN(n467) );
  AO21D0 U492 ( .A1(n471), .A2(i2[0]), .B(n467), .Z(n466) );
  OAI33D0 U493 ( .A1(n469), .A2(n468), .A3(n467), .B1(n466), .B2(i2[1]), .B3(
        n468), .ZN(n476) );
  CKXOR2D0 U494 ( .A1(i2[4]), .A2(DataI[28]), .Z(n470) );
  AOI21D0 U495 ( .A1(DataI[25]), .A2(n232), .B(n470), .ZN(n475) );
  CKND0 U496 ( .CLK(DataI[26]), .CN(n472) );
  OAI22D0 U497 ( .A1(i2[2]), .A2(n472), .B1(i2[0]), .B2(n471), .ZN(n473) );
  NR4D0 U498 ( .A1(n473), .A2(DataI[29]), .A3(DataI[31]), .A4(DataI[30]), .ZN(
        n474) );
  ND4D0 U499 ( .A1(n477), .A2(n476), .A3(n475), .A4(n474), .ZN(N279) );
  IND2D0 U500 ( .A1(i2[3]), .B1(DataI[19]), .ZN(n489) );
  CKND0 U501 ( .CLK(DataI[16]), .CN(n483) );
  IOA21D0 U502 ( .A1(n483), .A2(i2[0]), .B(DataI[17]), .ZN(n481) );
  INR2D0 U503 ( .A1(i2[2]), .B1(DataI[18]), .ZN(n480) );
  INR2D0 U504 ( .A1(i2[3]), .B1(DataI[19]), .ZN(n479) );
  AO21D0 U505 ( .A1(n483), .A2(i2[0]), .B(n479), .Z(n478) );
  OAI33D0 U506 ( .A1(n481), .A2(n480), .A3(n479), .B1(n478), .B2(i2[1]), .B3(
        n480), .ZN(n488) );
  CKXOR2D0 U507 ( .A1(i2[4]), .A2(DataI[20]), .Z(n482) );
  AOI21D0 U508 ( .A1(DataI[17]), .A2(n232), .B(n482), .ZN(n487) );
  CKND0 U509 ( .CLK(DataI[18]), .CN(n484) );
  OAI22D0 U510 ( .A1(i2[2]), .A2(n484), .B1(i2[0]), .B2(n483), .ZN(n485) );
  NR4D0 U511 ( .A1(n485), .A2(DataI[21]), .A3(DataI[23]), .A4(DataI[22]), .ZN(
        n486) );
  ND4D0 U512 ( .A1(n489), .A2(n488), .A3(n487), .A4(n486), .ZN(N280) );
  IND2D0 U513 ( .A1(i2[3]), .B1(DataI[11]), .ZN(n501) );
  CKND0 U514 ( .CLK(DataI[8]), .CN(n495) );
  IOA21D0 U515 ( .A1(n495), .A2(i2[0]), .B(DataI[9]), .ZN(n493) );
  INR2D0 U516 ( .A1(i2[2]), .B1(DataI[10]), .ZN(n492) );
  INR2D0 U517 ( .A1(i2[3]), .B1(DataI[11]), .ZN(n491) );
  AO21D0 U518 ( .A1(n495), .A2(i2[0]), .B(n491), .Z(n490) );
  OAI33D0 U519 ( .A1(n493), .A2(n492), .A3(n491), .B1(n490), .B2(i2[1]), .B3(
        n492), .ZN(n500) );
  CKXOR2D0 U520 ( .A1(i2[4]), .A2(DataI[12]), .Z(n494) );
  AOI21D0 U521 ( .A1(DataI[9]), .A2(n232), .B(n494), .ZN(n499) );
  CKND0 U522 ( .CLK(DataI[10]), .CN(n496) );
  OAI22D0 U523 ( .A1(i2[2]), .A2(n496), .B1(i2[0]), .B2(n495), .ZN(n497) );
  NR4D0 U524 ( .A1(n497), .A2(DataI[13]), .A3(DataI[15]), .A4(DataI[14]), .ZN(
        n498) );
  ND4D0 U525 ( .A1(n501), .A2(n500), .A3(n499), .A4(n498), .ZN(N281) );
  IND2D0 U526 ( .A1(i2[3]), .B1(DataI[3]), .ZN(n513) );
  CKND0 U527 ( .CLK(DataI[0]), .CN(n507) );
  IOA21D0 U528 ( .A1(n507), .A2(i2[0]), .B(DataI[1]), .ZN(n505) );
  INR2D0 U529 ( .A1(i2[2]), .B1(DataI[2]), .ZN(n504) );
  INR2D0 U530 ( .A1(i2[3]), .B1(DataI[3]), .ZN(n503) );
  AO21D0 U531 ( .A1(n507), .A2(i2[0]), .B(n503), .Z(n502) );
  OAI33D0 U532 ( .A1(n505), .A2(n504), .A3(n503), .B1(n502), .B2(i2[1]), .B3(
        n504), .ZN(n512) );
  CKXOR2D0 U533 ( .A1(i2[4]), .A2(DataI[4]), .Z(n506) );
  AOI21D0 U534 ( .A1(DataI[1]), .A2(n232), .B(n506), .ZN(n511) );
  CKND0 U535 ( .CLK(DataI[2]), .CN(n508) );
  OAI22D0 U536 ( .A1(i2[2]), .A2(n508), .B1(i2[0]), .B2(n507), .ZN(n509) );
  NR4D0 U537 ( .A1(n509), .A2(DataI[5]), .A3(DataI[7]), .A4(DataI[6]), .ZN(
        n510) );
  ND4D0 U538 ( .A1(n513), .A2(n512), .A3(n511), .A4(n510), .ZN(N282) );
  AN3D0 U539 ( .A1(N285), .A2(N284), .A3(N286), .Z(n514) );
  AN3D0 U540 ( .A1(N288), .A2(N287), .A3(n514), .Z(N289) );
  AN3D0 U541 ( .A1(N320), .A2(N319), .A3(N321), .Z(n515) );
  AN3D0 U542 ( .A1(N323), .A2(N322), .A3(n515), .Z(N324) );
  AN3D0 U543 ( .A1(N371), .A2(N370), .A3(N372), .Z(n516) );
  AN3D0 U544 ( .A1(N374), .A2(N373), .A3(n516), .Z(N375) );
  AN3D0 U545 ( .A1(N405), .A2(N404), .A3(N406), .Z(n517) );
  AN3D0 U546 ( .A1(N408), .A2(N407), .A3(n517), .Z(N409) );
  AN3D0 U547 ( .A1(N456), .A2(N455), .A3(N457), .Z(n518) );
  AN3D0 U548 ( .A1(N459), .A2(N458), .A3(n518), .Z(N460) );
endmodule


module Mem_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, ClkR, 
        ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, ClockR, ClockW, Dreadyr, \Storage[31][32] ,
         \Storage[31][31] , \Storage[31][30] , \Storage[31][29] ,
         \Storage[31][28] , \Storage[31][27] , \Storage[31][26] ,
         \Storage[31][25] , \Storage[31][24] , \Storage[31][23] ,
         \Storage[31][22] , \Storage[31][21] , \Storage[31][20] ,
         \Storage[31][19] , \Storage[31][18] , \Storage[31][17] ,
         \Storage[31][16] , \Storage[31][15] , \Storage[31][14] ,
         \Storage[31][13] , \Storage[31][12] , \Storage[31][11] ,
         \Storage[31][10] , \Storage[31][9] , \Storage[31][8] ,
         \Storage[31][7] , \Storage[31][6] , \Storage[31][5] ,
         \Storage[31][4] , \Storage[31][3] , \Storage[31][2] ,
         \Storage[31][1] , \Storage[31][0] , \Storage[30][32] ,
         \Storage[30][31] , \Storage[30][30] , \Storage[30][29] ,
         \Storage[30][28] , \Storage[30][27] , \Storage[30][26] ,
         \Storage[30][25] , \Storage[30][24] , \Storage[30][23] ,
         \Storage[30][22] , \Storage[30][21] , \Storage[30][20] ,
         \Storage[30][19] , \Storage[30][18] , \Storage[30][17] ,
         \Storage[30][16] , \Storage[30][15] , \Storage[30][14] ,
         \Storage[30][13] , \Storage[30][12] , \Storage[30][11] ,
         \Storage[30][10] , \Storage[30][9] , \Storage[30][8] ,
         \Storage[30][7] , \Storage[30][6] , \Storage[30][5] ,
         \Storage[30][4] , \Storage[30][3] , \Storage[30][2] ,
         \Storage[30][1] , \Storage[30][0] , \Storage[29][32] ,
         \Storage[29][31] , \Storage[29][30] , \Storage[29][29] ,
         \Storage[29][28] , \Storage[29][27] , \Storage[29][26] ,
         \Storage[29][25] , \Storage[29][24] , \Storage[29][23] ,
         \Storage[29][22] , \Storage[29][21] , \Storage[29][20] ,
         \Storage[29][19] , \Storage[29][18] , \Storage[29][17] ,
         \Storage[29][16] , \Storage[29][15] , \Storage[29][14] ,
         \Storage[29][13] , \Storage[29][12] , \Storage[29][11] ,
         \Storage[29][10] , \Storage[29][9] , \Storage[29][8] ,
         \Storage[29][7] , \Storage[29][6] , \Storage[29][5] ,
         \Storage[29][4] , \Storage[29][3] , \Storage[29][2] ,
         \Storage[29][1] , \Storage[29][0] , \Storage[28][32] ,
         \Storage[28][31] , \Storage[28][30] , \Storage[28][29] ,
         \Storage[28][28] , \Storage[28][27] , \Storage[28][26] ,
         \Storage[28][25] , \Storage[28][24] , \Storage[28][23] ,
         \Storage[28][22] , \Storage[28][21] , \Storage[28][20] ,
         \Storage[28][19] , \Storage[28][18] , \Storage[28][17] ,
         \Storage[28][16] , \Storage[28][15] , \Storage[28][14] ,
         \Storage[28][13] , \Storage[28][12] , \Storage[28][11] ,
         \Storage[28][10] , \Storage[28][9] , \Storage[28][8] ,
         \Storage[28][7] , \Storage[28][6] , \Storage[28][5] ,
         \Storage[28][4] , \Storage[28][3] , \Storage[28][2] ,
         \Storage[28][1] , \Storage[28][0] , \Storage[27][32] ,
         \Storage[27][31] , \Storage[27][30] , \Storage[27][29] ,
         \Storage[27][28] , \Storage[27][27] , \Storage[27][26] ,
         \Storage[27][25] , \Storage[27][24] , \Storage[27][23] ,
         \Storage[27][22] , \Storage[27][21] , \Storage[27][20] ,
         \Storage[27][19] , \Storage[27][18] , \Storage[27][17] ,
         \Storage[27][16] , \Storage[27][15] , \Storage[27][14] ,
         \Storage[27][13] , \Storage[27][12] , \Storage[27][11] ,
         \Storage[27][10] , \Storage[27][9] , \Storage[27][8] ,
         \Storage[27][7] , \Storage[27][6] , \Storage[27][5] ,
         \Storage[27][4] , \Storage[27][3] , \Storage[27][2] ,
         \Storage[27][1] , \Storage[27][0] , \Storage[26][32] ,
         \Storage[26][31] , \Storage[26][30] , \Storage[26][29] ,
         \Storage[26][28] , \Storage[26][27] , \Storage[26][26] ,
         \Storage[26][25] , \Storage[26][24] , \Storage[26][23] ,
         \Storage[26][22] , \Storage[26][21] , \Storage[26][20] ,
         \Storage[26][19] , \Storage[26][18] , \Storage[26][17] ,
         \Storage[26][16] , \Storage[26][15] , \Storage[26][14] ,
         \Storage[26][13] , \Storage[26][12] , \Storage[26][11] ,
         \Storage[26][10] , \Storage[26][9] , \Storage[26][8] ,
         \Storage[26][7] , \Storage[26][6] , \Storage[26][5] ,
         \Storage[26][4] , \Storage[26][3] , \Storage[26][2] ,
         \Storage[26][1] , \Storage[26][0] , \Storage[25][32] ,
         \Storage[25][31] , \Storage[25][30] , \Storage[25][29] ,
         \Storage[25][28] , \Storage[25][27] , \Storage[25][26] ,
         \Storage[25][25] , \Storage[25][24] , \Storage[25][23] ,
         \Storage[25][22] , \Storage[25][21] , \Storage[25][20] ,
         \Storage[25][19] , \Storage[25][18] , \Storage[25][17] ,
         \Storage[25][16] , \Storage[25][15] , \Storage[25][14] ,
         \Storage[25][13] , \Storage[25][12] , \Storage[25][11] ,
         \Storage[25][10] , \Storage[25][9] , \Storage[25][8] ,
         \Storage[25][7] , \Storage[25][6] , \Storage[25][5] ,
         \Storage[25][4] , \Storage[25][3] , \Storage[25][2] ,
         \Storage[25][1] , \Storage[25][0] , \Storage[24][32] ,
         \Storage[24][31] , \Storage[24][30] , \Storage[24][29] ,
         \Storage[24][28] , \Storage[24][27] , \Storage[24][26] ,
         \Storage[24][25] , \Storage[24][24] , \Storage[24][23] ,
         \Storage[24][22] , \Storage[24][21] , \Storage[24][20] ,
         \Storage[24][19] , \Storage[24][18] , \Storage[24][17] ,
         \Storage[24][16] , \Storage[24][15] , \Storage[24][14] ,
         \Storage[24][13] , \Storage[24][12] , \Storage[24][11] ,
         \Storage[24][10] , \Storage[24][9] , \Storage[24][8] ,
         \Storage[24][7] , \Storage[24][6] , \Storage[24][5] ,
         \Storage[24][4] , \Storage[24][3] , \Storage[24][2] ,
         \Storage[24][1] , \Storage[24][0] , \Storage[23][32] ,
         \Storage[23][31] , \Storage[23][30] , \Storage[23][29] ,
         \Storage[23][28] , \Storage[23][27] , \Storage[23][26] ,
         \Storage[23][25] , \Storage[23][24] , \Storage[23][23] ,
         \Storage[23][22] , \Storage[23][21] , \Storage[23][20] ,
         \Storage[23][19] , \Storage[23][18] , \Storage[23][17] ,
         \Storage[23][16] , \Storage[23][15] , \Storage[23][14] ,
         \Storage[23][13] , \Storage[23][12] , \Storage[23][11] ,
         \Storage[23][10] , \Storage[23][9] , \Storage[23][8] ,
         \Storage[23][7] , \Storage[23][6] , \Storage[23][5] ,
         \Storage[23][4] , \Storage[23][3] , \Storage[23][2] ,
         \Storage[23][1] , \Storage[23][0] , \Storage[22][32] ,
         \Storage[22][31] , \Storage[22][30] , \Storage[22][29] ,
         \Storage[22][28] , \Storage[22][27] , \Storage[22][26] ,
         \Storage[22][25] , \Storage[22][24] , \Storage[22][23] ,
         \Storage[22][22] , \Storage[22][21] , \Storage[22][20] ,
         \Storage[22][19] , \Storage[22][18] , \Storage[22][17] ,
         \Storage[22][16] , \Storage[22][15] , \Storage[22][14] ,
         \Storage[22][13] , \Storage[22][12] , \Storage[22][11] ,
         \Storage[22][10] , \Storage[22][9] , \Storage[22][8] ,
         \Storage[22][7] , \Storage[22][6] , \Storage[22][5] ,
         \Storage[22][4] , \Storage[22][3] , \Storage[22][2] ,
         \Storage[22][1] , \Storage[22][0] , \Storage[21][32] ,
         \Storage[21][31] , \Storage[21][30] , \Storage[21][29] ,
         \Storage[21][28] , \Storage[21][27] , \Storage[21][26] ,
         \Storage[21][25] , \Storage[21][24] , \Storage[21][23] ,
         \Storage[21][22] , \Storage[21][21] , \Storage[21][20] ,
         \Storage[21][19] , \Storage[21][18] , \Storage[21][17] ,
         \Storage[21][16] , \Storage[21][15] , \Storage[21][14] ,
         \Storage[21][13] , \Storage[21][12] , \Storage[21][11] ,
         \Storage[21][10] , \Storage[21][9] , \Storage[21][8] ,
         \Storage[21][7] , \Storage[21][6] , \Storage[21][5] ,
         \Storage[21][4] , \Storage[21][3] , \Storage[21][2] ,
         \Storage[21][1] , \Storage[21][0] , \Storage[20][32] ,
         \Storage[20][31] , \Storage[20][30] , \Storage[20][29] ,
         \Storage[20][28] , \Storage[20][27] , \Storage[20][26] ,
         \Storage[20][25] , \Storage[20][24] , \Storage[20][23] ,
         \Storage[20][22] , \Storage[20][21] , \Storage[20][20] ,
         \Storage[20][19] , \Storage[20][18] , \Storage[20][17] ,
         \Storage[20][16] , \Storage[20][15] , \Storage[20][14] ,
         \Storage[20][13] , \Storage[20][12] , \Storage[20][11] ,
         \Storage[20][10] , \Storage[20][9] , \Storage[20][8] ,
         \Storage[20][7] , \Storage[20][6] , \Storage[20][5] ,
         \Storage[20][4] , \Storage[20][3] , \Storage[20][2] ,
         \Storage[20][1] , \Storage[20][0] , \Storage[19][32] ,
         \Storage[19][31] , \Storage[19][30] , \Storage[19][29] ,
         \Storage[19][28] , \Storage[19][27] , \Storage[19][26] ,
         \Storage[19][25] , \Storage[19][24] , \Storage[19][23] ,
         \Storage[19][22] , \Storage[19][21] , \Storage[19][20] ,
         \Storage[19][19] , \Storage[19][18] , \Storage[19][17] ,
         \Storage[19][16] , \Storage[19][15] , \Storage[19][14] ,
         \Storage[19][13] , \Storage[19][12] , \Storage[19][11] ,
         \Storage[19][10] , \Storage[19][9] , \Storage[19][8] ,
         \Storage[19][7] , \Storage[19][6] , \Storage[19][5] ,
         \Storage[19][4] , \Storage[19][3] , \Storage[19][2] ,
         \Storage[19][1] , \Storage[19][0] , \Storage[18][32] ,
         \Storage[18][31] , \Storage[18][30] , \Storage[18][29] ,
         \Storage[18][28] , \Storage[18][27] , \Storage[18][26] ,
         \Storage[18][25] , \Storage[18][24] , \Storage[18][23] ,
         \Storage[18][22] , \Storage[18][21] , \Storage[18][20] ,
         \Storage[18][19] , \Storage[18][18] , \Storage[18][17] ,
         \Storage[18][16] , \Storage[18][15] , \Storage[18][14] ,
         \Storage[18][13] , \Storage[18][12] , \Storage[18][11] ,
         \Storage[18][10] , \Storage[18][9] , \Storage[18][8] ,
         \Storage[18][7] , \Storage[18][6] , \Storage[18][5] ,
         \Storage[18][4] , \Storage[18][3] , \Storage[18][2] ,
         \Storage[18][1] , \Storage[18][0] , \Storage[17][32] ,
         \Storage[17][31] , \Storage[17][30] , \Storage[17][29] ,
         \Storage[17][28] , \Storage[17][27] , \Storage[17][26] ,
         \Storage[17][25] , \Storage[17][24] , \Storage[17][23] ,
         \Storage[17][22] , \Storage[17][21] , \Storage[17][20] ,
         \Storage[17][19] , \Storage[17][18] , \Storage[17][17] ,
         \Storage[17][16] , \Storage[17][15] , \Storage[17][14] ,
         \Storage[17][13] , \Storage[17][12] , \Storage[17][11] ,
         \Storage[17][10] , \Storage[17][9] , \Storage[17][8] ,
         \Storage[17][7] , \Storage[17][6] , \Storage[17][5] ,
         \Storage[17][4] , \Storage[17][3] , \Storage[17][2] ,
         \Storage[17][1] , \Storage[17][0] , \Storage[16][32] ,
         \Storage[16][31] , \Storage[16][30] , \Storage[16][29] ,
         \Storage[16][28] , \Storage[16][27] , \Storage[16][26] ,
         \Storage[16][25] , \Storage[16][24] , \Storage[16][23] ,
         \Storage[16][22] , \Storage[16][21] , \Storage[16][20] ,
         \Storage[16][19] , \Storage[16][18] , \Storage[16][17] ,
         \Storage[16][16] , \Storage[16][15] , \Storage[16][14] ,
         \Storage[16][13] , \Storage[16][12] , \Storage[16][11] ,
         \Storage[16][10] , \Storage[16][9] , \Storage[16][8] ,
         \Storage[16][7] , \Storage[16][6] , \Storage[16][5] ,
         \Storage[16][4] , \Storage[16][3] , \Storage[16][2] ,
         \Storage[16][1] , \Storage[16][0] , \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N85, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  OR2D1 U3 ( .A1(n605), .A2(Dreadyr), .Z(n107) );
  XNR4D1 U18 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n84) );
  XOR4D1 U19 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n83) );
  XOR4D1 U20 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n80) );
  XOR4D1 U21 ( .A1(n615), .A2(n613), .A3(DataI[16]), .A4(n617), .Z(n77) );
  XNR4D1 U22 ( .A1(n611), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), .ZN(n74) );
  XOR4D1 U27 ( .A1(n90), .A2(N72), .A3(n91), .A4(N75), .Z(n89) );
  XNR4D1 U28 ( .A1(N69), .A2(N68), .A3(N71), .A4(N70), .ZN(n91) );
  XNR4D1 U33 ( .A1(N51), .A2(N50), .A3(N53), .A4(N52), .ZN(n97) );
  XOR4D1 U34 ( .A1(N55), .A2(N54), .A3(N57), .A4(N56), .Z(n96) );
  XNR4D1 U35 ( .A1(N62), .A2(N61), .A3(N64), .A4(N63), .ZN(n93) );
  XNR4D1 U36 ( .A1(N80), .A2(N78), .A3(N82), .A4(N81), .ZN(n87) );
  AN2D2 U81 ( .A1(ClkW), .A2(n46), .Z(ClockW) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(DataI[10]), .E(n32), .CP(ClockW), .CDN(
        n577), .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(DataI[9]), .E(n32), .CP(ClockW), .CDN(
        n588), .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(DataI[8]), .E(n32), .CP(ClockW), .CDN(
        n596), .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(n611), .E(n32), .CP(ClockW), .CDN(n572), 
        .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(n609), .E(n32), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(n607), .E(n32), .CP(ClockW), .CDN(n577), 
        .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(DataI[4]), .E(n32), .CP(ClockW), .CDN(
        n567), .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(DataI[3]), .E(n32), .CP(ClockW), .CDN(
        n577), .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(DataI[2]), .E(n32), .CP(ClockW), .CDN(
        n582), .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(DataI[1]), .E(n32), .CP(ClockW), .CDN(
        n588), .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(DataI[0]), .E(n32), .CP(ClockW), .CDN(
        n580), .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(DataI[10]), .E(n31), .CP(ClockW), .CDN(
        n595), .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(DataI[9]), .E(n31), .CP(ClockW), .CDN(
        n592), .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(DataI[8]), .E(n31), .CP(ClockW), .CDN(
        n592), .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(n611), .E(n31), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(n609), .E(n31), .CP(ClockW), .CDN(n598), 
        .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(n607), .E(n31), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(DataI[4]), .E(n31), .CP(ClockW), .CDN(
        n576), .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(DataI[3]), .E(n31), .CP(ClockW), .CDN(
        n581), .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(DataI[2]), .E(n31), .CP(ClockW), .CDN(
        n598), .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(DataI[1]), .E(n31), .CP(ClockW), .CDN(
        n597), .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(DataI[0]), .E(n31), .CP(ClockW), .CDN(
        n576), .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(DataI[10]), .E(n30), .CP(ClockW), .CDN(
        n581), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(DataI[9]), .E(n30), .CP(ClockW), .CDN(
        n589), .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(n30), .CP(ClockW), .CDN(
        n586), .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(DataI[7]), .E(n30), .CP(ClockW), .CDN(
        n585), .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(n609), .E(n30), .CP(ClockW), .CDN(n580), 
        .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(n607), .E(n30), .CP(ClockW), .CDN(n581), 
        .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(DataI[4]), .E(n30), .CP(ClockW), .CDN(
        n582), .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(DataI[3]), .E(n30), .CP(ClockW), .CDN(
        n578), .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(DataI[2]), .E(n30), .CP(ClockW), .CDN(
        n577), .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(DataI[1]), .E(n30), .CP(ClockW), .CDN(
        n576), .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(DataI[0]), .E(n30), .CP(ClockW), .CDN(
        n579), .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(DataI[10]), .E(n29), .CP(ClockW), .CDN(
        n585), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(DataI[9]), .E(n29), .CP(ClockW), .CDN(
        n573), .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(DataI[8]), .E(n29), .CP(ClockW), .CDN(
        n596), .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(DataI[7]), .E(n29), .CP(ClockW), .CDN(
        n596), .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(n609), .E(n29), .CP(ClockW), .CDN(n596), 
        .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(n607), .E(n29), .CP(ClockW), .CDN(n596), 
        .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(DataI[4]), .E(n29), .CP(ClockW), .CDN(
        n596), .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(DataI[3]), .E(n29), .CP(ClockW), .CDN(
        n596), .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(DataI[2]), .E(n29), .CP(ClockW), .CDN(
        n596), .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(n29), .CP(ClockW), .CDN(
        n596), .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(DataI[0]), .E(n29), .CP(ClockW), .CDN(
        n571), .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(DataI[10]), .E(n28), .CP(ClockW), .CDN(
        n576), .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(DataI[9]), .E(n28), .CP(ClockW), .CDN(
        n586), .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(DataI[8]), .E(n28), .CP(ClockW), .CDN(
        n585), .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(DataI[7]), .E(n28), .CP(ClockW), .CDN(
        n584), .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(n609), .E(n28), .CP(ClockW), .CDN(n583), 
        .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(n607), .E(n28), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(DataI[4]), .E(n28), .CP(ClockW), .CDN(
        n581), .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(DataI[3]), .E(n28), .CP(ClockW), .CDN(
        n580), .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(DataI[2]), .E(n28), .CP(ClockW), .CDN(
        n579), .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(DataI[1]), .E(n28), .CP(ClockW), .CDN(
        n578), .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(DataI[0]), .E(n28), .CP(ClockW), .CDN(
        n577), .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(DataI[10]), .E(n27), .CP(ClockW), .CDN(
        n571), .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(DataI[9]), .E(n27), .CP(ClockW), .CDN(
        n568), .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(DataI[8]), .E(n27), .CP(ClockW), .CDN(
        n580), .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(n611), .E(n27), .CP(ClockW), .CDN(n588), 
        .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(n609), .E(n27), .CP(ClockW), .CDN(n587), 
        .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(n607), .E(n27), .CP(ClockW), .CDN(n571), 
        .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(DataI[4]), .E(n27), .CP(ClockW), .CDN(
        n581), .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(DataI[3]), .E(n27), .CP(ClockW), .CDN(
        n586), .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(DataI[2]), .E(n27), .CP(ClockW), .CDN(
        n588), .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(DataI[1]), .E(n27), .CP(ClockW), .CDN(
        n581), .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(DataI[0]), .E(n27), .CP(ClockW), .CDN(
        n588), .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(DataI[10]), .E(n26), .CP(ClockW), .CDN(
        n577), .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(DataI[9]), .E(n26), .CP(ClockW), .CDN(
        n565), .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(DataI[8]), .E(n26), .CP(ClockW), .CDN(
        n596), .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(DataI[7]), .E(n26), .CP(ClockW), .CDN(
        n596), .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(n609), .E(n26), .CP(ClockW), .CDN(n588), 
        .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(n607), .E(n26), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(DataI[4]), .E(n26), .CP(ClockW), .CDN(
        n568), .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(DataI[3]), .E(n26), .CP(ClockW), .CDN(
        n584), .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(DataI[2]), .E(n26), .CP(ClockW), .CDN(
        n585), .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(DataI[1]), .E(n26), .CP(ClockW), .CDN(
        n598), .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(DataI[0]), .E(n26), .CP(ClockW), .CDN(
        n597), .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(DataI[10]), .E(n25), .CP(ClockW), .CDN(
        n591), .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(DataI[9]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(DataI[8]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(DataI[7]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(n609), .E(n25), .CP(ClockW), .CDN(n602), 
        .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(n607), .E(n25), .CP(ClockW), .CDN(n602), 
        .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(DataI[4]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(DataI[3]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(DataI[2]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(DataI[1]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(DataI[0]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(DataI[10]), .E(n24), .CP(ClockW), .CDN(
        n568), .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(DataI[9]), .E(n24), .CP(ClockW), .CDN(
        n580), .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(DataI[8]), .E(n24), .CP(ClockW), .CDN(
        n592), .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(DataI[7]), .E(n24), .CP(ClockW), .CDN(
        n578), .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(n609), .E(n24), .CP(ClockW), .CDN(n595), 
        .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(n607), .E(n24), .CP(ClockW), .CDN(n569), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(DataI[4]), .E(n24), .CP(ClockW), .CDN(
        n603), .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(DataI[3]), .E(n24), .CP(ClockW), .CDN(
        n592), .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(DataI[2]), .E(n24), .CP(ClockW), .CDN(
        n577), .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(DataI[1]), .E(n24), .CP(ClockW), .CDN(
        n595), .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(DataI[0]), .E(n24), .CP(ClockW), .CDN(
        n586), .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(DataI[10]), .E(n23), .CP(ClockW), .CDN(
        n593), .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(DataI[9]), .E(n23), .CP(ClockW), .CDN(
        n597), .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(DataI[8]), .E(n23), .CP(ClockW), .CDN(
        n589), .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(DataI[7]), .E(n23), .CP(ClockW), .CDN(
        n599), .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(n609), .E(n23), .CP(ClockW), .CDN(n594), 
        .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(n607), .E(n23), .CP(ClockW), .CDN(n601), 
        .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(DataI[4]), .E(n23), .CP(ClockW), .CDN(
        n595), .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(DataI[3]), .E(n23), .CP(ClockW), .CDN(
        n599), .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(DataI[2]), .E(n23), .CP(ClockW), .CDN(
        n595), .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(DataI[1]), .E(n23), .CP(ClockW), .CDN(
        n601), .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(DataI[0]), .E(n23), .CP(ClockW), .CDN(
        n594), .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(DataI[10]), .E(n22), .CP(ClockW), .CDN(
        n589), .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(DataI[9]), .E(n22), .CP(ClockW), .CDN(
        n592), .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(DataI[8]), .E(n22), .CP(ClockW), .CDN(
        n604), .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(DataI[7]), .E(n22), .CP(ClockW), .CDN(
        n604), .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(n609), .E(n22), .CP(ClockW), .CDN(n604), 
        .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(n607), .E(n22), .CP(ClockW), .CDN(n604), 
        .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(DataI[4]), .E(n22), .CP(ClockW), .CDN(
        n603), .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(DataI[3]), .E(n22), .CP(ClockW), .CDN(
        n566), .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(DataI[2]), .E(n22), .CP(ClockW), .CDN(
        n604), .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(DataI[1]), .E(n22), .CP(ClockW), .CDN(
        n588), .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(DataI[0]), .E(n22), .CP(ClockW), .CDN(
        n604), .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(DataI[10]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(DataI[9]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(DataI[7]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n609), .E(n21), .CP(ClockW), .CDN(n561), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n607), .E(n21), .CP(ClockW), .CDN(n561), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(DataI[4]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(DataI[3]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(DataI[2]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(DataI[1]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(DataI[0]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(n20), .CP(ClockW), .CDN(
        n561), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(DataI[9]), .E(n20), .CP(ClockW), .CDN(
        n595), .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(DataI[8]), .E(n20), .CP(ClockW), .CDN(
        n594), .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(n20), .CP(ClockW), .CDN(
        n594), .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n609), .E(n20), .CP(ClockW), .CDN(n593), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n607), .E(n20), .CP(ClockW), .CDN(n598), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(DataI[4]), .E(n20), .CP(ClockW), .CDN(
        n598), .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(n20), .CP(ClockW), .CDN(
        n597), .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(DataI[2]), .E(n20), .CP(ClockW), .CDN(
        n594), .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(n20), .CP(ClockW), .CDN(
        n593), .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(DataI[0]), .E(n20), .CP(ClockW), .CDN(
        n598), .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(DataI[10]), .E(n19), .CP(ClockW), .CDN(
        n583), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(DataI[9]), .E(n19), .CP(ClockW), .CDN(
        n604), .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(DataI[8]), .E(n19), .CP(ClockW), .CDN(
        n603), .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n611), .E(n19), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n609), .E(n19), .CP(ClockW), .CDN(n600), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n607), .E(n19), .CP(ClockW), .CDN(n591), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(DataI[4]), .E(n19), .CP(ClockW), .CDN(
        n592), .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(DataI[3]), .E(n19), .CP(ClockW), .CDN(
        n604), .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(DataI[2]), .E(n19), .CP(ClockW), .CDN(
        n599), .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(DataI[1]), .E(n19), .CP(ClockW), .CDN(
        n600), .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(DataI[0]), .E(n19), .CP(ClockW), .CDN(
        n591), .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(DataI[10]), .E(n18), .CP(ClockW), .CDN(
        n589), .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(n18), .CP(ClockW), .CDN(n563), .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(DataI[8]), .E(n18), .CP(ClockW), .CDN(n601), .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n611), .E(n18), .CP(ClockW), .CDN(n601), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n609), .E(n18), .CP(ClockW), .CDN(n601), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n607), .E(n18), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(n18), .CP(ClockW), .CDN(n603), .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(DataI[3]), .E(n18), .CP(ClockW), .CDN(n576), .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(DataI[2]), .E(n18), .CP(ClockW), .CDN(n562), .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(DataI[1]), .E(n18), .CP(ClockW), .CDN(n600), .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(n18), .CP(ClockW), .CDN(n564), .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n17), .CP(ClockW), .CDN(n582), .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(n17), .CP(ClockW), .CDN(n582), .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n611), .E(n17), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n609), .E(n17), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n607), .E(n17), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n17), .CP(ClockW), .CDN(n582), .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n17), .CP(ClockW), .CDN(n582), .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n17), .CP(ClockW), .CDN(n582), .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n17), .CP(ClockW), .CDN(n582), .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n17), .CP(ClockW), .CDN(n582), .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n16), .CP(ClockW), .CDN(n579), .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(n16), .CP(ClockW), .CDN(n579), .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n611), .E(n16), .CP(ClockW), .CDN(n579), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n609), .E(n16), .CP(ClockW), .CDN(n579), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n607), .E(n16), .CP(ClockW), .CDN(n579), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n16), .CP(ClockW), .CDN(n579), .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n16), .CP(ClockW), .CDN(n579), .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n16), .CP(ClockW), .CDN(n579), .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(n16), .CP(ClockW), .CDN(n579), .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n16), .CP(ClockW), .CDN(n579), .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n15), .CP(ClockW), .CDN(n571), .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n15), .CP(ClockW), .CDN(n571), .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n611), .E(n15), .CP(ClockW), .CDN(n571), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n609), .E(n15), .CP(ClockW), .CDN(n571), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n607), .E(n15), .CP(ClockW), .CDN(n571), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n15), .CP(ClockW), .CDN(n571), .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(n15), .CP(ClockW), .CDN(n571), .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n15), .CP(ClockW), .CDN(n571), .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(n15), .CP(ClockW), .CDN(n571), .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(n15), .CP(ClockW), .CDN(n571), .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n14), .CP(ClockW), .CDN(n568), .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(n14), .CP(ClockW), .CDN(n568), .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n611), .E(n14), .CP(ClockW), .CDN(n568), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n609), .E(n14), .CP(ClockW), .CDN(n568), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n607), .E(n14), .CP(ClockW), .CDN(n568), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n14), .CP(ClockW), .CDN(n568), .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n14), .CP(ClockW), .CDN(n568), .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n14), .CP(ClockW), .CDN(n568), .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n14), .CP(ClockW), .CDN(n568), .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n14), .CP(ClockW), .CDN(n568), .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(DataI[10]), .E(n13), .CP(ClockW), .CDN(
        n592), .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(DataI[9]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(DataI[8]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(DataI[7]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(n609), .E(n13), .CP(ClockW), .CDN(n591), 
        .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(n607), .E(n13), .CP(ClockW), .CDN(n591), 
        .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(DataI[4]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(DataI[3]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(DataI[2]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(DataI[1]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(DataI[0]), .E(n13), .CP(ClockW), .CDN(
        n591), .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(DataI[10]), .E(n12), .CP(ClockW), .CDN(
        n591), .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(DataI[9]), .E(n12), .CP(ClockW), .CDN(
        n594), .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(DataI[8]), .E(n12), .CP(ClockW), .CDN(
        n595), .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(DataI[7]), .E(n12), .CP(ClockW), .CDN(
        n598), .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(n609), .E(n12), .CP(ClockW), .CDN(n597), 
        .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(n607), .E(n12), .CP(ClockW), .CDN(n593), 
        .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(DataI[4]), .E(n12), .CP(ClockW), .CDN(
        n594), .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(DataI[3]), .E(n12), .CP(ClockW), .CDN(
        n596), .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(DataI[2]), .E(n12), .CP(ClockW), .CDN(
        n595), .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(DataI[1]), .E(n12), .CP(ClockW), .CDN(
        n598), .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(DataI[0]), .E(n12), .CP(ClockW), .CDN(
        n597), .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(DataI[10]), .E(n11), .CP(ClockW), .CDN(
        n593), .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(DataI[9]), .E(n11), .CP(ClockW), .CDN(
        n584), .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(DataI[8]), .E(n11), .CP(ClockW), .CDN(
        n598), .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(DataI[7]), .E(n11), .CP(ClockW), .CDN(
        n595), .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(n609), .E(n11), .CP(ClockW), .CDN(n575), 
        .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(n607), .E(n11), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(DataI[4]), .E(n11), .CP(ClockW), .CDN(
        n602), .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(DataI[3]), .E(n11), .CP(ClockW), .CDN(
        n591), .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(DataI[2]), .E(n11), .CP(ClockW), .CDN(
        n593), .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(DataI[1]), .E(n11), .CP(ClockW), .CDN(
        n596), .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(DataI[0]), .E(n11), .CP(ClockW), .CDN(
        n574), .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(DataI[10]), .E(n10), .CP(ClockW), .CDN(
        n600), .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(DataI[9]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(DataI[8]), .E(n10), .CP(ClockW), .CDN(
        n603), .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(DataI[7]), .E(n10), .CP(ClockW), .CDN(
        n589), .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(n609), .E(n10), .CP(ClockW), .CDN(n604), 
        .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(n607), .E(n10), .CP(ClockW), .CDN(n589), 
        .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(DataI[4]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(DataI[3]), .E(n10), .CP(ClockW), .CDN(
        n603), .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(DataI[2]), .E(n10), .CP(ClockW), .CDN(
        n589), .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(DataI[1]), .E(n10), .CP(ClockW), .CDN(
        n588), .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(DataI[0]), .E(n10), .CP(ClockW), .CDN(
        n598), .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(DataI[10]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(DataI[9]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(DataI[7]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n609), .E(n9), .CP(ClockW), .CDN(n564), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n607), .E(n9), .CP(ClockW), .CDN(n564), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(DataI[4]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(DataI[3]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(DataI[2]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(DataI[1]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(DataI[0]), .E(n9), .CP(ClockW), .CDN(n564), .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(DataI[10]), .E(n8), .CP(ClockW), .CDN(
        n594), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(DataI[9]), .E(n8), .CP(ClockW), .CDN(n598), .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(DataI[8]), .E(n8), .CP(ClockW), .CDN(n597), .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n611), .E(n8), .CP(ClockW), .CDN(n600), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n609), .E(n8), .CP(ClockW), .CDN(n601), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n607), .E(n8), .CP(ClockW), .CDN(n595), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(DataI[4]), .E(n8), .CP(ClockW), .CDN(n600), .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(DataI[3]), .E(n8), .CP(ClockW), .CDN(n601), .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(DataI[2]), .E(n8), .CP(ClockW), .CDN(n594), .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(DataI[1]), .E(n8), .CP(ClockW), .CDN(n600), .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(DataI[0]), .E(n8), .CP(ClockW), .CDN(n601), .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(DataI[10]), .E(n7), .CP(ClockW), .CDN(
        n597), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(DataI[9]), .E(n7), .CP(ClockW), .CDN(n599), .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(DataI[8]), .E(n7), .CP(ClockW), .CDN(n598), .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n611), .E(n7), .CP(ClockW), .CDN(n597), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n609), .E(n7), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n607), .E(n7), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(DataI[4]), .E(n7), .CP(ClockW), .CDN(n600), .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(DataI[3]), .E(n7), .CP(ClockW), .CDN(n601), .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(DataI[2]), .E(n7), .CP(ClockW), .CDN(n563), .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(DataI[1]), .E(n7), .CP(ClockW), .CDN(n598), .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(DataI[0]), .E(n7), .CP(ClockW), .CDN(n597), .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(DataI[10]), .E(n6), .CP(ClockW), .CDN(
        n584), .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(n6), .CP(ClockW), .CDN(n108), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(DataI[8]), .E(n6), .CP(ClockW), .CDN(n603), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n611), .E(n6), .CP(ClockW), .CDN(n603), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n609), .E(n6), .CP(ClockW), .CDN(n603), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n607), .E(n6), .CP(ClockW), .CDN(n568), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(n6), .CP(ClockW), .CDN(n589), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(DataI[3]), .E(n6), .CP(ClockW), .CDN(n562), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(DataI[2]), .E(n6), .CP(ClockW), .CDN(n593), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(DataI[1]), .E(n6), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(n6), .CP(ClockW), .CDN(n601), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n611), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n609), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n607), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(n5), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n611), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n609), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n607), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(n4), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n611), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n609), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n607), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(n3), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n611), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n609), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n607), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n2), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(DataI[10]), .E(n1), .CP(ClockW), .CDN(
        n590), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(DataI[9]), .E(n1), .CP(ClockW), .CDN(n603), .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(DataI[8]), .E(n1), .CP(ClockW), .CDN(n592), .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(DataI[7]), .E(n1), .CP(ClockW), .CDN(n590), .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(n609), .E(n1), .CP(ClockW), .CDN(n590), 
        .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(n607), .E(n1), .CP(ClockW), .CDN(n590), 
        .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(DataI[4]), .E(n1), .CP(ClockW), .CDN(n590), .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(DataI[3]), .E(n1), .CP(ClockW), .CDN(n590), .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(DataI[2]), .E(n1), .CP(ClockW), .CDN(n590), .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(DataI[1]), .E(n1), .CP(ClockW), .CDN(n589), .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(DataI[0]), .E(n1), .CP(ClockW), .CDN(n590), .Q(\Storage[31][0] ) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(N85), .E(n32), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(DataI[31]), .E(n32), .CP(ClockW), .CDN(
        n586), .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(DataI[30]), .E(n32), .CP(ClockW), .CDN(
        n580), .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(DataI[29]), .E(n32), .CP(ClockW), .CDN(
        n580), .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(DataI[28]), .E(n32), .CP(ClockW), .CDN(
        n585), .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(DataI[27]), .E(n32), .CP(ClockW), .CDN(
        n584), .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(DataI[26]), .E(n32), .CP(ClockW), .CDN(
        n582), .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(DataI[25]), .E(n32), .CP(ClockW), .CDN(
        n588), .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(DataI[24]), .E(n32), .CP(ClockW), .CDN(
        n585), .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(DataI[23]), .E(n32), .CP(ClockW), .CDN(
        n577), .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(DataI[22]), .E(n32), .CP(ClockW), .CDN(
        n582), .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(DataI[21]), .E(n32), .CP(ClockW), .CDN(
        n579), .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(DataI[20]), .E(n32), .CP(ClockW), .CDN(
        n578), .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(DataI[19]), .E(n32), .CP(ClockW), .CDN(
        n581), .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(DataI[18]), .E(n32), .CP(ClockW), .CDN(
        n588), .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(DataI[17]), .E(n32), .CP(ClockW), .CDN(
        n580), .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(DataI[16]), .E(n32), .CP(ClockW), .CDN(
        n576), .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(n617), .E(n32), .CP(ClockW), .CDN(n583), 
        .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(n615), .E(n32), .CP(ClockW), .CDN(n578), 
        .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(DataI[13]), .E(n32), .CP(ClockW), .CDN(
        n578), .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(DataI[12]), .E(n32), .CP(ClockW), .CDN(
        n582), .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(DataI[11]), .E(n32), .CP(ClockW), .CDN(
        n580), .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(N85), .E(n31), .CP(ClockW), .CDN(n562), 
        .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(DataI[31]), .E(n31), .CP(ClockW), .CDN(
        n597), .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(DataI[30]), .E(n31), .CP(ClockW), .CDN(
        n584), .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(DataI[29]), .E(n31), .CP(ClockW), .CDN(
        n584), .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(DataI[28]), .E(n31), .CP(ClockW), .CDN(
        n592), .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(DataI[27]), .E(n31), .CP(ClockW), .CDN(
        n586), .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(DataI[26]), .E(n31), .CP(ClockW), .CDN(
        n585), .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(DataI[25]), .E(n31), .CP(ClockW), .CDN(
        n578), .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(DataI[24]), .E(n31), .CP(ClockW), .CDN(
        n592), .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(DataI[23]), .E(n31), .CP(ClockW), .CDN(
        n581), .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(DataI[22]), .E(n31), .CP(ClockW), .CDN(
        n595), .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(DataI[21]), .E(n31), .CP(ClockW), .CDN(
        n598), .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(DataI[20]), .E(n31), .CP(ClockW), .CDN(
        n593), .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(DataI[19]), .E(n31), .CP(ClockW), .CDN(
        n594), .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(DataI[18]), .E(n31), .CP(ClockW), .CDN(
        n596), .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(DataI[17]), .E(n31), .CP(ClockW), .CDN(
        n593), .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(DataI[16]), .E(n31), .CP(ClockW), .CDN(
        n594), .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(n617), .E(n31), .CP(ClockW), .CDN(n593), 
        .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(n615), .E(n31), .CP(ClockW), .CDN(n594), 
        .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(DataI[13]), .E(n31), .CP(ClockW), .CDN(
        n596), .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(DataI[12]), .E(n31), .CP(ClockW), .CDN(
        n593), .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(DataI[11]), .E(n31), .CP(ClockW), .CDN(
        n594), .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(N85), .E(n30), .CP(ClockW), .CDN(n590), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(DataI[31]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(DataI[29]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(DataI[28]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(DataI[27]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(DataI[24]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(DataI[23]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(DataI[22]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(n30), .CP(ClockW), .CDN(
        n588), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(DataI[20]), .E(n30), .CP(ClockW), .CDN(
        n568), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(DataI[19]), .E(n30), .CP(ClockW), .CDN(
        n584), .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(n30), .CP(ClockW), .CDN(
        n585), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(DataI[17]), .E(n30), .CP(ClockW), .CDN(
        n586), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(DataI[16]), .E(n30), .CP(ClockW), .CDN(
        n580), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(DataI[15]), .E(n30), .CP(ClockW), .CDN(
        n581), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(n30), .CP(ClockW), .CDN(
        n582), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(DataI[13]), .E(n30), .CP(ClockW), .CDN(
        n578), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(DataI[12]), .E(n30), .CP(ClockW), .CDN(
        n577), .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(n30), .CP(ClockW), .CDN(
        n576), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(n560), .E(n29), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(DataI[31]), .E(n29), .CP(ClockW), .CDN(
        n580), .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(DataI[30]), .E(n29), .CP(ClockW), .CDN(
        n581), .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(DataI[29]), .E(n29), .CP(ClockW), .CDN(
        n582), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(DataI[28]), .E(n29), .CP(ClockW), .CDN(
        n576), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(DataI[27]), .E(n29), .CP(ClockW), .CDN(
        n579), .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(DataI[26]), .E(n29), .CP(ClockW), .CDN(
        n578), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(DataI[25]), .E(n29), .CP(ClockW), .CDN(
        n577), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(DataI[24]), .E(n29), .CP(ClockW), .CDN(
        n567), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(DataI[23]), .E(n29), .CP(ClockW), .CDN(
        n584), .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(DataI[22]), .E(n29), .CP(ClockW), .CDN(
        n571), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(DataI[21]), .E(n29), .CP(ClockW), .CDN(
        n568), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(DataI[20]), .E(n29), .CP(ClockW), .CDN(
        n582), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(DataI[19]), .E(n29), .CP(ClockW), .CDN(
        n581), .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(DataI[18]), .E(n29), .CP(ClockW), .CDN(
        n576), .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(DataI[17]), .E(n29), .CP(ClockW), .CDN(
        n579), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(DataI[16]), .E(n29), .CP(ClockW), .CDN(
        n578), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(DataI[15]), .E(n29), .CP(ClockW), .CDN(
        n577), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(DataI[14]), .E(n29), .CP(ClockW), .CDN(
        n581), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(DataI[13]), .E(n29), .CP(ClockW), .CDN(
        n567), .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(DataI[12]), .E(n29), .CP(ClockW), .CDN(
        n571), .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(DataI[11]), .E(n29), .CP(ClockW), .CDN(
        n568), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(N85), .E(n28), .CP(ClockW), .CDN(n596), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(DataI[31]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(DataI[30]), .E(n28), .CP(ClockW), .CDN(
        n589), .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(DataI[29]), .E(n28), .CP(ClockW), .CDN(
        n589), .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(DataI[28]), .E(n28), .CP(ClockW), .CDN(
        n589), .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(DataI[27]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(DataI[26]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(DataI[25]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(DataI[24]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(DataI[23]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(DataI[22]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(DataI[21]), .E(n28), .CP(ClockW), .CDN(
        n562), .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(DataI[20]), .E(n28), .CP(ClockW), .CDN(
        n568), .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(DataI[19]), .E(n28), .CP(ClockW), .CDN(
        n566), .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(DataI[18]), .E(n28), .CP(ClockW), .CDN(
        n572), .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(DataI[17]), .E(n28), .CP(ClockW), .CDN(
        n571), .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(DataI[16]), .E(n28), .CP(ClockW), .CDN(
        n570), .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(DataI[15]), .E(n28), .CP(ClockW), .CDN(
        n569), .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(DataI[14]), .E(n28), .CP(ClockW), .CDN(
        n587), .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(DataI[13]), .E(n28), .CP(ClockW), .CDN(
        n586), .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(DataI[12]), .E(n28), .CP(ClockW), .CDN(
        n585), .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(DataI[11]), .E(n28), .CP(ClockW), .CDN(
        n584), .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(n560), .E(n27), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(DataI[31]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(DataI[30]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(DataI[29]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(DataI[28]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(DataI[27]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(DataI[26]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(DataI[25]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(DataI[24]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(DataI[23]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(DataI[22]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(DataI[21]), .E(n27), .CP(ClockW), .CDN(
        n567), .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(DataI[20]), .E(n27), .CP(ClockW), .CDN(
        n569), .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(DataI[19]), .E(n27), .CP(ClockW), .CDN(
        n582), .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(DataI[18]), .E(n27), .CP(ClockW), .CDN(
        n588), .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(DataI[17]), .E(n27), .CP(ClockW), .CDN(
        n571), .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(DataI[16]), .E(n27), .CP(ClockW), .CDN(
        n568), .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(n617), .E(n27), .CP(ClockW), .CDN(n588), 
        .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(n615), .E(n27), .CP(ClockW), .CDN(n584), 
        .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(DataI[13]), .E(n27), .CP(ClockW), .CDN(
        n585), .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(DataI[12]), .E(n27), .CP(ClockW), .CDN(
        n584), .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(DataI[11]), .E(n27), .CP(ClockW), .CDN(
        n587), .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(n560), .E(n26), .CP(ClockW), .CDN(n565), 
        .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(DataI[31]), .E(n26), .CP(ClockW), .CDN(
        n581), .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(DataI[30]), .E(n26), .CP(ClockW), .CDN(
        n568), .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(DataI[29]), .E(n26), .CP(ClockW), .CDN(
        n596), .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(DataI[28]), .E(n26), .CP(ClockW), .CDN(
        n588), .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(DataI[27]), .E(n26), .CP(ClockW), .CDN(
        n578), .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(DataI[26]), .E(n26), .CP(ClockW), .CDN(
        n580), .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(DataI[25]), .E(n26), .CP(ClockW), .CDN(
        n582), .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(DataI[24]), .E(n26), .CP(ClockW), .CDN(
        n576), .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(DataI[23]), .E(n26), .CP(ClockW), .CDN(
        n580), .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(DataI[22]), .E(n26), .CP(ClockW), .CDN(
        n566), .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(DataI[21]), .E(n26), .CP(ClockW), .CDN(
        n596), .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(DataI[20]), .E(n26), .CP(ClockW), .CDN(
        n567), .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(DataI[19]), .E(n26), .CP(ClockW), .CDN(
        n579), .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(DataI[18]), .E(n26), .CP(ClockW), .CDN(
        n571), .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(DataI[17]), .E(n26), .CP(ClockW), .CDN(
        n579), .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(DataI[16]), .E(n26), .CP(ClockW), .CDN(
        n572), .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(DataI[15]), .E(n26), .CP(ClockW), .CDN(
        n596), .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(DataI[14]), .E(n26), .CP(ClockW), .CDN(
        n588), .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(DataI[13]), .E(n26), .CP(ClockW), .CDN(
        n576), .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(DataI[12]), .E(n26), .CP(ClockW), .CDN(
        n571), .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(DataI[11]), .E(n26), .CP(ClockW), .CDN(
        n585), .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(N85), .E(n25), .CP(ClockW), .CDN(n591), 
        .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(DataI[31]), .E(n25), .CP(ClockW), .CDN(
        n585), .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(DataI[30]), .E(n25), .CP(ClockW), .CDN(
        n588), .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(DataI[29]), .E(n25), .CP(ClockW), .CDN(
        n575), .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(DataI[28]), .E(n25), .CP(ClockW), .CDN(
        n578), .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(DataI[27]), .E(n25), .CP(ClockW), .CDN(
        n571), .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(DataI[26]), .E(n25), .CP(ClockW), .CDN(
        n571), .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(DataI[25]), .E(n25), .CP(ClockW), .CDN(
        n568), .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(DataI[24]), .E(n25), .CP(ClockW), .CDN(
        n579), .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(DataI[23]), .E(n25), .CP(ClockW), .CDN(
        n568), .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(DataI[22]), .E(n25), .CP(ClockW), .CDN(
        n588), .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(DataI[21]), .E(n25), .CP(ClockW), .CDN(
        n596), .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(DataI[20]), .E(n25), .CP(ClockW), .CDN(
        n596), .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(DataI[19]), .E(n25), .CP(ClockW), .CDN(
        n578), .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(DataI[18]), .E(n25), .CP(ClockW), .CDN(
        n567), .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(DataI[17]), .E(n25), .CP(ClockW), .CDN(
        n602), .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(DataI[16]), .E(n25), .CP(ClockW), .CDN(
        n588), .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(DataI[15]), .E(n25), .CP(ClockW), .CDN(
        n592), .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(DataI[14]), .E(n25), .CP(ClockW), .CDN(
        n581), .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(n613), .E(n25), .CP(ClockW), .CDN(n592), 
        .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(DataI[12]), .E(n25), .CP(ClockW), .CDN(
        n586), .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(DataI[11]), .E(n25), .CP(ClockW), .CDN(
        n574), .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(n560), .E(n24), .CP(ClockW), .CDN(n602), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(DataI[31]), .E(n24), .CP(ClockW), .CDN(
        n590), .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(DataI[30]), .E(n24), .CP(ClockW), .CDN(
        n577), .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(DataI[29]), .E(n24), .CP(ClockW), .CDN(
        n595), .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(DataI[28]), .E(n24), .CP(ClockW), .CDN(
        n594), .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(DataI[27]), .E(n24), .CP(ClockW), .CDN(
        n593), .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(DataI[26]), .E(n24), .CP(ClockW), .CDN(
        n596), .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(DataI[25]), .E(n24), .CP(ClockW), .CDN(
        n570), .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(DataI[24]), .E(n24), .CP(ClockW), .CDN(
        n602), .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(DataI[23]), .E(n24), .CP(ClockW), .CDN(
        n577), .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(DataI[22]), .E(n24), .CP(ClockW), .CDN(
        n602), .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(DataI[21]), .E(n24), .CP(ClockW), .CDN(
        n571), .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(DataI[20]), .E(n24), .CP(ClockW), .CDN(
        n591), .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(DataI[19]), .E(n24), .CP(ClockW), .CDN(
        n579), .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(DataI[18]), .E(n24), .CP(ClockW), .CDN(
        n596), .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(DataI[17]), .E(n24), .CP(ClockW), .CDN(
        n602), .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(DataI[16]), .E(n24), .CP(ClockW), .CDN(
        n568), .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(DataI[15]), .E(n24), .CP(ClockW), .CDN(
        n592), .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(DataI[14]), .E(n24), .CP(ClockW), .CDN(
        n593), .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(n613), .E(n24), .CP(ClockW), .CDN(n594), 
        .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(DataI[12]), .E(n24), .CP(ClockW), .CDN(
        n595), .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(DataI[11]), .E(n24), .CP(ClockW), .CDN(
        n571), .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(N85), .E(n23), .CP(ClockW), .CDN(n584), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(DataI[31]), .E(n23), .CP(ClockW), .CDN(
        n603), .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(DataI[30]), .E(n23), .CP(ClockW), .CDN(
        n592), .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(DataI[29]), .E(n23), .CP(ClockW), .CDN(
        n592), .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(DataI[28]), .E(n23), .CP(ClockW), .CDN(
        n582), .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(DataI[27]), .E(n23), .CP(ClockW), .CDN(
        n599), .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(DataI[26]), .E(n23), .CP(ClockW), .CDN(
        n590), .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(DataI[25]), .E(n23), .CP(ClockW), .CDN(
        n604), .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(DataI[24]), .E(n23), .CP(ClockW), .CDN(
        n579), .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(DataI[23]), .E(n23), .CP(ClockW), .CDN(
        n599), .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(DataI[22]), .E(n23), .CP(ClockW), .CDN(
        n571), .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(DataI[21]), .E(n23), .CP(ClockW), .CDN(
        n604), .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(DataI[20]), .E(n23), .CP(ClockW), .CDN(
        n567), .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(DataI[19]), .E(n23), .CP(ClockW), .CDN(
        n584), .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(DataI[18]), .E(n23), .CP(ClockW), .CDN(
        n568), .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(DataI[17]), .E(n23), .CP(ClockW), .CDN(
        n585), .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(DataI[16]), .E(n23), .CP(ClockW), .CDN(
        n565), .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(DataI[15]), .E(n23), .CP(ClockW), .CDN(
        n597), .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(DataI[14]), .E(n23), .CP(ClockW), .CDN(
        n599), .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(n613), .E(n23), .CP(ClockW), .CDN(n598), 
        .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(DataI[12]), .E(n23), .CP(ClockW), .CDN(
        n594), .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(DataI[11]), .E(n23), .CP(ClockW), .CDN(
        n599), .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(n560), .E(n22), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(DataI[31]), .E(n22), .CP(ClockW), .CDN(
        n601), .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(DataI[30]), .E(n22), .CP(ClockW), .CDN(
        n600), .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(DataI[29]), .E(n22), .CP(ClockW), .CDN(
        n600), .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(DataI[28]), .E(n22), .CP(ClockW), .CDN(
        n600), .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(DataI[27]), .E(n22), .CP(ClockW), .CDN(
        n571), .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(DataI[26]), .E(n22), .CP(ClockW), .CDN(
        n604), .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(DataI[25]), .E(n22), .CP(ClockW), .CDN(
        n599), .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(DataI[24]), .E(n22), .CP(ClockW), .CDN(
        n599), .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(DataI[23]), .E(n22), .CP(ClockW), .CDN(
        n599), .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(DataI[22]), .E(n22), .CP(ClockW), .CDN(
        n579), .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(DataI[21]), .E(n22), .CP(ClockW), .CDN(
        n592), .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(DataI[20]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(DataI[19]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(DataI[18]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(DataI[17]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(DataI[16]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(DataI[15]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(DataI[14]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(DataI[13]), .E(n22), .CP(ClockW), .CDN(
        n563), .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(DataI[12]), .E(n22), .CP(ClockW), .CDN(
        n604), .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(DataI[11]), .E(n22), .CP(ClockW), .CDN(
        n604), .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N85), .E(n21), .CP(ClockW), .CDN(n564), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(n21), .CP(ClockW), .CDN(
        n564), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(DataI[29]), .E(n21), .CP(ClockW), .CDN(
        n564), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(n21), .CP(ClockW), .CDN(
        n564), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(n21), .CP(ClockW), .CDN(
        n564), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(DataI[22]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(DataI[20]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(DataI[17]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(DataI[15]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(DataI[12]), .E(n21), .CP(ClockW), .CDN(
        n562), .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(n21), .CP(ClockW), .CDN(
        n561), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n560), .E(n20), .CP(ClockW), .CDN(n561), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(DataI[31]), .E(n20), .CP(ClockW), .CDN(
        n561), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(DataI[30]), .E(n20), .CP(ClockW), .CDN(
        n591), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(n20), .CP(ClockW), .CDN(
        n561), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(DataI[28]), .E(n20), .CP(ClockW), .CDN(
        n591), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(DataI[27]), .E(n20), .CP(ClockW), .CDN(
        n561), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(DataI[26]), .E(n20), .CP(ClockW), .CDN(
        n591), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(DataI[25]), .E(n20), .CP(ClockW), .CDN(
        n561), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(DataI[24]), .E(n20), .CP(ClockW), .CDN(
        n591), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(DataI[23]), .E(n20), .CP(ClockW), .CDN(
        n561), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(DataI[22]), .E(n20), .CP(ClockW), .CDN(
        n562), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(DataI[21]), .E(n20), .CP(ClockW), .CDN(
        n591), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(n20), .CP(ClockW), .CDN(
        n108), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(DataI[19]), .E(n20), .CP(ClockW), .CDN(
        n108), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(DataI[18]), .E(n20), .CP(ClockW), .CDN(
        n108), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(n20), .CP(ClockW), .CDN(
        n108), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(DataI[16]), .E(n20), .CP(ClockW), .CDN(
        n603), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(n20), .CP(ClockW), .CDN(
        n591), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(DataI[14]), .E(n20), .CP(ClockW), .CDN(
        n604), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(DataI[13]), .E(n20), .CP(ClockW), .CDN(
        n604), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(DataI[12]), .E(n20), .CP(ClockW), .CDN(
        n563), .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(DataI[11]), .E(n20), .CP(ClockW), .CDN(
        n562), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N85), .E(n19), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(DataI[31]), .E(n19), .CP(ClockW), .CDN(
        n108), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(DataI[30]), .E(n19), .CP(ClockW), .CDN(
        n602), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(DataI[29]), .E(n19), .CP(ClockW), .CDN(
        n592), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(DataI[28]), .E(n19), .CP(ClockW), .CDN(
        n576), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(DataI[27]), .E(n19), .CP(ClockW), .CDN(
        n562), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(DataI[26]), .E(n19), .CP(ClockW), .CDN(
        n599), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(DataI[25]), .E(n19), .CP(ClockW), .CDN(
        n563), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(DataI[24]), .E(n19), .CP(ClockW), .CDN(
        n108), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(DataI[23]), .E(n19), .CP(ClockW), .CDN(
        n108), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(DataI[22]), .E(n19), .CP(ClockW), .CDN(
        n108), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(DataI[21]), .E(n19), .CP(ClockW), .CDN(
        n108), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(DataI[20]), .E(n19), .CP(ClockW), .CDN(
        n600), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(DataI[19]), .E(n19), .CP(ClockW), .CDN(
        n578), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(DataI[18]), .E(n19), .CP(ClockW), .CDN(
        n599), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(DataI[17]), .E(n19), .CP(ClockW), .CDN(
        n600), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(DataI[16]), .E(n19), .CP(ClockW), .CDN(
        n580), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n617), .E(n19), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n615), .E(n19), .CP(ClockW), .CDN(n600), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n613), .E(n19), .CP(ClockW), .CDN(n567), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(DataI[12]), .E(n19), .CP(ClockW), .CDN(
        n599), .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(DataI[11]), .E(n19), .CP(ClockW), .CDN(
        n600), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(n560), .E(n18), .CP(ClockW), .CDN(n577), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(DataI[31]), .E(n18), .CP(ClockW), .CDN(
        n108), .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(DataI[30]), .E(n18), .CP(ClockW), .CDN(
        n599), .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(DataI[29]), .E(n18), .CP(ClockW), .CDN(
        n600), .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(DataI[28]), .E(n18), .CP(ClockW), .CDN(
        n586), .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(DataI[27]), .E(n18), .CP(ClockW), .CDN(
        n590), .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(DataI[26]), .E(n18), .CP(ClockW), .CDN(
        n592), .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(DataI[25]), .E(n18), .CP(ClockW), .CDN(
        n582), .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(DataI[24]), .E(n18), .CP(ClockW), .CDN(
        n591), .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(DataI[23]), .E(n18), .CP(ClockW), .CDN(
        n593), .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(n18), .CP(ClockW), .CDN(
        n594), .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(DataI[21]), .E(n18), .CP(ClockW), .CDN(
        n576), .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(DataI[20]), .E(n18), .CP(ClockW), .CDN(
        n594), .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(DataI[19]), .E(n18), .CP(ClockW), .CDN(
        n599), .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(DataI[18]), .E(n18), .CP(ClockW), .CDN(
        n568), .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(DataI[17]), .E(n18), .CP(ClockW), .CDN(
        n593), .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(DataI[16]), .E(n18), .CP(ClockW), .CDN(
        n603), .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n617), .E(n18), .CP(ClockW), .CDN(n589), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n615), .E(n18), .CP(ClockW), .CDN(n594), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n613), .E(n18), .CP(ClockW), .CDN(n108), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(n18), .CP(ClockW), .CDN(
        n589), .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(DataI[11]), .E(n18), .CP(ClockW), .CDN(
        n591), .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N85), .E(n17), .CP(ClockW), .CDN(n585), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(n17), .CP(ClockW), .CDN(
        n584), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n617), .E(n17), .CP(ClockW), .CDN(n583), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n615), .E(n17), .CP(ClockW), .CDN(n583), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n613), .E(n17), .CP(ClockW), .CDN(n583), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n17), .CP(ClockW), .CDN(
        n583), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(n560), .E(n16), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(n16), .CP(ClockW), .CDN(
        n581), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n617), .E(n16), .CP(ClockW), .CDN(n580), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n615), .E(n16), .CP(ClockW), .CDN(n580), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n613), .E(n16), .CP(ClockW), .CDN(n580), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n16), .CP(ClockW), .CDN(
        n580), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N85), .E(n15), .CP(ClockW), .CDN(n573), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(n15), .CP(ClockW), .CDN(
        n577), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(n15), .CP(ClockW), .CDN(
        n573), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(n15), .CP(ClockW), .CDN(
        n574), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n15), .CP(ClockW), .CDN(
        n575), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n15), .CP(ClockW), .CDN(
        n586), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n15), .CP(ClockW), .CDN(
        n584), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(n15), .CP(ClockW), .CDN(
        n582), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n15), .CP(ClockW), .CDN(
        n581), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(n15), .CP(ClockW), .CDN(
        n580), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n15), .CP(ClockW), .CDN(
        n579), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n15), .CP(ClockW), .CDN(
        n578), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n617), .E(n15), .CP(ClockW), .CDN(n572), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n615), .E(n15), .CP(ClockW), .CDN(n572), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n613), .E(n15), .CP(ClockW), .CDN(n572), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n15), .CP(ClockW), .CDN(
        n572), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(n560), .E(n14), .CP(ClockW), .CDN(n571), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(n14), .CP(ClockW), .CDN(
        n570), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n617), .E(n14), .CP(ClockW), .CDN(n569), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n615), .E(n14), .CP(ClockW), .CDN(n569), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n613), .E(n14), .CP(ClockW), .CDN(n569), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n14), .CP(ClockW), .CDN(
        n569), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(n560), .E(n13), .CP(ClockW), .CDN(n580), 
        .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(DataI[31]), .E(n13), .CP(ClockW), .CDN(
        n597), .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(DataI[30]), .E(n13), .CP(ClockW), .CDN(
        n595), .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(DataI[29]), .E(n13), .CP(ClockW), .CDN(
        n593), .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(DataI[28]), .E(n13), .CP(ClockW), .CDN(
        n594), .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(DataI[27]), .E(n13), .CP(ClockW), .CDN(
        n598), .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(DataI[26]), .E(n13), .CP(ClockW), .CDN(
        n597), .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(DataI[25]), .E(n13), .CP(ClockW), .CDN(
        n596), .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(DataI[24]), .E(n13), .CP(ClockW), .CDN(
        n595), .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(DataI[23]), .E(n13), .CP(ClockW), .CDN(
        n593), .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(DataI[22]), .E(n13), .CP(ClockW), .CDN(
        n594), .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(DataI[21]), .E(n13), .CP(ClockW), .CDN(
        n598), .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(DataI[20]), .E(n13), .CP(ClockW), .CDN(
        n577), .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(DataI[19]), .E(n13), .CP(ClockW), .CDN(
        n592), .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(DataI[18]), .E(n13), .CP(ClockW), .CDN(
        n579), .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(DataI[17]), .E(n13), .CP(ClockW), .CDN(
        n603), .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(DataI[16]), .E(n13), .CP(ClockW), .CDN(
        n595), .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(DataI[15]), .E(n13), .CP(ClockW), .CDN(
        n593), .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(DataI[14]), .E(n13), .CP(ClockW), .CDN(
        n594), .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(n613), .E(n13), .CP(ClockW), .CDN(n598), 
        .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(DataI[12]), .E(n13), .CP(ClockW), .CDN(
        n597), .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(DataI[11]), .E(n13), .CP(ClockW), .CDN(
        n578), .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(N85), .E(n12), .CP(ClockW), .CDN(n578), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(DataI[31]), .E(n12), .CP(ClockW), .CDN(
        n592), .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(DataI[30]), .E(n12), .CP(ClockW), .CDN(
        n602), .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(DataI[29]), .E(n12), .CP(ClockW), .CDN(
        n595), .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(DataI[28]), .E(n12), .CP(ClockW), .CDN(
        n584), .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(DataI[27]), .E(n12), .CP(ClockW), .CDN(
        n592), .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(DataI[26]), .E(n12), .CP(ClockW), .CDN(
        n573), .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(DataI[25]), .E(n12), .CP(ClockW), .CDN(
        n595), .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(DataI[24]), .E(n12), .CP(ClockW), .CDN(
        n585), .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(DataI[23]), .E(n12), .CP(ClockW), .CDN(
        n598), .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(DataI[22]), .E(n12), .CP(ClockW), .CDN(
        n581), .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(DataI[21]), .E(n12), .CP(ClockW), .CDN(
        n579), .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(DataI[20]), .E(n12), .CP(ClockW), .CDN(
        n585), .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(DataI[19]), .E(n12), .CP(ClockW), .CDN(
        n592), .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(DataI[18]), .E(n12), .CP(ClockW), .CDN(
        n590), .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(DataI[17]), .E(n12), .CP(ClockW), .CDN(
        n570), .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(DataI[16]), .E(n12), .CP(ClockW), .CDN(
        n595), .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(DataI[15]), .E(n12), .CP(ClockW), .CDN(
        n594), .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(DataI[14]), .E(n12), .CP(ClockW), .CDN(
        n593), .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(DataI[13]), .E(n12), .CP(ClockW), .CDN(
        n597), .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(DataI[12]), .E(n12), .CP(ClockW), .CDN(
        n598), .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(DataI[11]), .E(n12), .CP(ClockW), .CDN(
        n597), .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(n560), .E(n11), .CP(ClockW), .CDN(n593), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(DataI[31]), .E(n11), .CP(ClockW), .CDN(
        n568), .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(DataI[30]), .E(n11), .CP(ClockW), .CDN(
        n591), .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(DataI[29]), .E(n11), .CP(ClockW), .CDN(
        n592), .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(DataI[28]), .E(n11), .CP(ClockW), .CDN(
        n596), .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(DataI[27]), .E(n11), .CP(ClockW), .CDN(
        n592), .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(DataI[26]), .E(n11), .CP(ClockW), .CDN(
        n580), .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(DataI[25]), .E(n11), .CP(ClockW), .CDN(
        n588), .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(DataI[24]), .E(n11), .CP(ClockW), .CDN(
        n592), .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(DataI[23]), .E(n11), .CP(ClockW), .CDN(
        n595), .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(DataI[22]), .E(n11), .CP(ClockW), .CDN(
        n562), .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(DataI[21]), .E(n11), .CP(ClockW), .CDN(
        n594), .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(DataI[20]), .E(n11), .CP(ClockW), .CDN(
        n579), .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(DataI[19]), .E(n11), .CP(ClockW), .CDN(
        n568), .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(DataI[18]), .E(n11), .CP(ClockW), .CDN(
        n592), .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(DataI[17]), .E(n11), .CP(ClockW), .CDN(
        n595), .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(DataI[16]), .E(n11), .CP(ClockW), .CDN(
        n579), .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(DataI[15]), .E(n11), .CP(ClockW), .CDN(
        n594), .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(DataI[14]), .E(n11), .CP(ClockW), .CDN(
        n581), .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(DataI[13]), .E(n11), .CP(ClockW), .CDN(
        n593), .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(DataI[12]), .E(n11), .CP(ClockW), .CDN(
        n595), .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(DataI[11]), .E(n11), .CP(ClockW), .CDN(
        n597), .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(N85), .E(n10), .CP(ClockW), .CDN(n603), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(DataI[31]), .E(n10), .CP(ClockW), .CDN(
        n603), .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(DataI[30]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(DataI[29]), .E(n10), .CP(ClockW), .CDN(
        n585), .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(DataI[28]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(DataI[27]), .E(n10), .CP(ClockW), .CDN(
        n586), .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(DataI[26]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(DataI[25]), .E(n10), .CP(ClockW), .CDN(
        n603), .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(DataI[24]), .E(n10), .CP(ClockW), .CDN(
        n571), .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(DataI[23]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(DataI[22]), .E(n10), .CP(ClockW), .CDN(
        n579), .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(DataI[21]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(DataI[20]), .E(n10), .CP(ClockW), .CDN(
        n601), .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(DataI[19]), .E(n10), .CP(ClockW), .CDN(
        n600), .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(DataI[18]), .E(n10), .CP(ClockW), .CDN(
        n601), .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(DataI[17]), .E(n10), .CP(ClockW), .CDN(
        n600), .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(DataI[16]), .E(n10), .CP(ClockW), .CDN(
        n603), .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(DataI[15]), .E(n10), .CP(ClockW), .CDN(
        n601), .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(DataI[14]), .E(n10), .CP(ClockW), .CDN(
        n600), .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(DataI[13]), .E(n10), .CP(ClockW), .CDN(
        n604), .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(DataI[12]), .E(n10), .CP(ClockW), .CDN(
        n590), .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(DataI[11]), .E(n10), .CP(ClockW), .CDN(
        n601), .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(n560), .E(n9), .CP(ClockW), .CDN(n597), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(DataI[29]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(DataI[22]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(n9), .CP(ClockW), .CDN(
        n602), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(DataI[20]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(DataI[17]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(DataI[15]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(DataI[12]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(n9), .CP(ClockW), .CDN(
        n564), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N85), .E(n8), .CP(ClockW), .CDN(n597), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(DataI[31]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(DataI[30]), .E(n8), .CP(ClockW), .CDN(
        n595), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(DataI[29]), .E(n8), .CP(ClockW), .CDN(
        n594), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(DataI[28]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(DataI[27]), .E(n8), .CP(ClockW), .CDN(
        n593), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(DataI[26]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(DataI[25]), .E(n8), .CP(ClockW), .CDN(
        n595), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(DataI[24]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(DataI[23]), .E(n8), .CP(ClockW), .CDN(
        n597), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(DataI[22]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(DataI[21]), .E(n8), .CP(ClockW), .CDN(
        n595), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(DataI[20]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(DataI[19]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(DataI[18]), .E(n8), .CP(ClockW), .CDN(
        n600), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(DataI[17]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(DataI[16]), .E(n8), .CP(ClockW), .CDN(
        n593), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n617), .E(n8), .CP(ClockW), .CDN(n600), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n615), .E(n8), .CP(ClockW), .CDN(n601), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(DataI[13]), .E(n8), .CP(ClockW), .CDN(
        n598), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(DataI[12]), .E(n8), .CP(ClockW), .CDN(
        n600), .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(DataI[11]), .E(n8), .CP(ClockW), .CDN(
        n601), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(n560), .E(n7), .CP(ClockW), .CDN(n593), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(DataI[31]), .E(n7), .CP(ClockW), .CDN(
        n598), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(DataI[30]), .E(n7), .CP(ClockW), .CDN(
        n597), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(DataI[29]), .E(n7), .CP(ClockW), .CDN(
        n598), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(DataI[28]), .E(n7), .CP(ClockW), .CDN(
        n597), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(DataI[27]), .E(n7), .CP(ClockW), .CDN(
        n600), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(DataI[26]), .E(n7), .CP(ClockW), .CDN(
        n601), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(DataI[25]), .E(n7), .CP(ClockW), .CDN(
        n598), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(DataI[24]), .E(n7), .CP(ClockW), .CDN(
        n597), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(DataI[23]), .E(n7), .CP(ClockW), .CDN(
        n598), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(DataI[22]), .E(n7), .CP(ClockW), .CDN(
        n600), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(DataI[21]), .E(n7), .CP(ClockW), .CDN(
        n601), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(DataI[20]), .E(n7), .CP(ClockW), .CDN(
        n597), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(DataI[19]), .E(n7), .CP(ClockW), .CDN(
        n582), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(DataI[18]), .E(n7), .CP(ClockW), .CDN(
        n599), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(DataI[17]), .E(n7), .CP(ClockW), .CDN(
        n595), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(DataI[16]), .E(n7), .CP(ClockW), .CDN(
        n597), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n617), .E(n7), .CP(ClockW), .CDN(n598), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n615), .E(n7), .CP(ClockW), .CDN(n600), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(DataI[13]), .E(n7), .CP(ClockW), .CDN(
        n601), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(DataI[12]), .E(n7), .CP(ClockW), .CDN(
        n599), .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(DataI[11]), .E(n7), .CP(ClockW), .CDN(
        n599), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N85), .E(n6), .CP(ClockW), .CDN(n589), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(DataI[31]), .E(n6), .CP(ClockW), .CDN(
        n593), .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(DataI[30]), .E(n6), .CP(ClockW), .CDN(
        n584), .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(DataI[29]), .E(n6), .CP(ClockW), .CDN(
        n604), .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(DataI[28]), .E(n6), .CP(ClockW), .CDN(
        n593), .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(DataI[27]), .E(n6), .CP(ClockW), .CDN(
        n563), .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(DataI[26]), .E(n6), .CP(ClockW), .CDN(
        n576), .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(DataI[25]), .E(n6), .CP(ClockW), .CDN(
        n599), .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(DataI[24]), .E(n6), .CP(ClockW), .CDN(
        n600), .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(DataI[23]), .E(n6), .CP(ClockW), .CDN(
        n585), .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(n6), .CP(ClockW), .CDN(
        n577), .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(DataI[21]), .E(n6), .CP(ClockW), .CDN(
        n589), .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(DataI[20]), .E(n6), .CP(ClockW), .CDN(
        n604), .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(DataI[19]), .E(n6), .CP(ClockW), .CDN(
        n571), .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(DataI[18]), .E(n6), .CP(ClockW), .CDN(
        n604), .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(DataI[17]), .E(n6), .CP(ClockW), .CDN(
        n589), .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(DataI[16]), .E(n6), .CP(ClockW), .CDN(
        n600), .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n617), .E(n6), .CP(ClockW), .CDN(n592), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n615), .E(n6), .CP(ClockW), .CDN(n604), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n613), .E(n6), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(n6), .CP(ClockW), .CDN(
        n589), .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(DataI[11]), .E(n6), .CP(ClockW), .CDN(
        n600), .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(n560), .E(n5), .CP(ClockW), .CDN(n108), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(n5), .CP(ClockW), .CDN(
        n587), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n617), .E(n5), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n615), .E(n5), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n613), .E(n5), .CP(ClockW), .CDN(n586), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n5), .CP(ClockW), .CDN(
        n586), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N85), .E(n4), .CP(ClockW), .CDN(n579), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(n4), .CP(ClockW), .CDN(
        n578), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n617), .E(n4), .CP(ClockW), .CDN(n577), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n615), .E(n4), .CP(ClockW), .CDN(n577), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n613), .E(n4), .CP(ClockW), .CDN(n577), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n4), .CP(ClockW), .CDN(
        n577), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(n560), .E(n3), .CP(ClockW), .CDN(n576), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n3), .CP(ClockW), .CDN(
        n575), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n617), .E(n3), .CP(ClockW), .CDN(n574), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n615), .E(n3), .CP(ClockW), .CDN(n574), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n613), .E(n3), .CP(ClockW), .CDN(n574), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n3), .CP(ClockW), .CDN(
        n574), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N85), .E(n2), .CP(ClockW), .CDN(n568), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n2), .CP(ClockW), .CDN(
        n567), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n617), .E(n2), .CP(ClockW), .CDN(n566), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n615), .E(n2), .CP(ClockW), .CDN(n566), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n613), .E(n2), .CP(ClockW), .CDN(n566), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(n2), .CP(ClockW), .CDN(
        n566), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(n560), .E(n1), .CP(ClockW), .CDN(n589), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(DataI[31]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(DataI[30]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(DataI[29]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(DataI[28]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(DataI[27]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(DataI[26]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][26] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(DataI[25]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(DataI[24]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(DataI[23]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(DataI[22]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(DataI[21]), .E(n1), .CP(ClockW), .CDN(
        n603), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(DataI[20]), .E(n1), .CP(ClockW), .CDN(
        n592), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(DataI[19]), .E(n1), .CP(ClockW), .CDN(
        n596), .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(DataI[18]), .E(n1), .CP(ClockW), .CDN(
        n578), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(DataI[17]), .E(n1), .CP(ClockW), .CDN(
        n577), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(DataI[16]), .E(n1), .CP(ClockW), .CDN(
        n591), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(DataI[15]), .E(n1), .CP(ClockW), .CDN(
        n591), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(DataI[14]), .E(n1), .CP(ClockW), .CDN(
        n590), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(n613), .E(n1), .CP(ClockW), .CDN(n590), 
        .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(DataI[12]), .E(n1), .CP(ClockW), .CDN(
        n590), .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(DataI[11]), .E(n1), .CP(ClockW), .CDN(
        n590), .Q(\Storage[31][11] ) );
  EDFCNQD1 Parityr_reg ( .D(N83), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        ParityErr) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N51), .E(Read), .CP(ClockR), .CDN(n564), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N52), .E(n605), .CP(ClockR), .CDN(n576), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N53), .E(n605), .CP(ClockR), .CDN(n576), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N54), .E(n605), .CP(ClockR), .CDN(n586), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N55), .E(n605), .CP(ClockR), .CDN(n571), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N56), .E(n605), .CP(ClockR), .CDN(n568), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N57), .E(n605), .CP(ClockR), .CDN(n579), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N58), .E(Read), .CP(ClockR), .CDN(n585), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N59), .E(Read), .CP(ClockR), .CDN(n584), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N60), .E(Read), .CP(ClockR), .CDN(n582), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N61), .E(Read), .CP(ClockR), .CDN(n581), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N62), .E(n605), .CP(ClockR), .CDN(n580), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N63), .E(n605), .CP(ClockR), .CDN(n590), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N64), .E(Read), .CP(ClockR), .CDN(n590), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N65), .E(Read), .CP(ClockR), .CDN(n590), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N66), .E(Read), .CP(ClockR), .CDN(n590), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N67), .E(Read), .CP(ClockR), .CDN(n590), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N68), .E(Read), .CP(ClockR), .CDN(n590), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N69), .E(Read), .CP(ClockR), .CDN(n590), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N70), .E(n605), .CP(ClockR), .CDN(n590), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N71), .E(n605), .CP(ClockR), .CDN(n590), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N72), .E(n605), .CP(ClockR), .CDN(n590), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N73), .E(n605), .CP(ClockR), .CDN(n590), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N74), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N75), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N76), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N77), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N78), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N79), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N80), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N81), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N82), .E(n605), .CP(ClockR), .CDN(n589), .Q(
        DataOr[0]) );
  BUFTD1 \DataO_tri[0]  ( .I(DataOr[0]), .OE(n619), .Z(DataO[0]) );
  BUFTD1 \DataO_tri[1]  ( .I(DataOr[1]), .OE(n620), .Z(DataO[1]) );
  BUFTD1 \DataO_tri[2]  ( .I(DataOr[2]), .OE(n621), .Z(DataO[2]) );
  DFCNQD1 Dreadyr_reg ( .D(n107), .CP(ClockR), .CDN(n565), .Q(Dreadyr) );
  BUFTD1 \DataO_tri[29]  ( .I(DataOr[29]), .OE(n620), .Z(DataO[29]) );
  BUFTD1 \DataO_tri[3]  ( .I(DataOr[3]), .OE(n621), .Z(DataO[3]) );
  BUFTD1 \DataO_tri[30]  ( .I(DataOr[30]), .OE(n621), .Z(DataO[30]) );
  BUFTD1 \DataO_tri[5]  ( .I(DataOr[5]), .OE(n621), .Z(DataO[5]) );
  BUFTD1 \DataO_tri[27]  ( .I(DataOr[27]), .OE(n620), .Z(DataO[27]) );
  BUFTD1 \DataO_tri[7]  ( .I(DataOr[7]), .OE(n621), .Z(DataO[7]) );
  BUFTD1 \DataO_tri[25]  ( .I(DataOr[25]), .OE(n620), .Z(DataO[25]) );
  BUFTD1 \DataO_tri[23]  ( .I(DataOr[23]), .OE(n620), .Z(DataO[23]) );
  BUFTD1 \DataO_tri[18]  ( .I(DataOr[18]), .OE(n619), .Z(DataO[18]) );
  BUFTD1 \DataO_tri[31]  ( .I(DataOr[31]), .OE(n621), .Z(DataO[31]) );
  BUFTD1 \DataO_tri[28]  ( .I(DataOr[28]), .OE(n620), .Z(DataO[28]) );
  BUFTD1 \DataO_tri[26]  ( .I(DataOr[26]), .OE(n620), .Z(DataO[26]) );
  BUFTD1 \DataO_tri[24]  ( .I(DataOr[24]), .OE(n620), .Z(DataO[24]) );
  BUFTD1 \DataO_tri[22]  ( .I(DataOr[22]), .OE(n620), .Z(DataO[22]) );
  BUFTD1 \DataO_tri[19]  ( .I(DataOr[19]), .OE(n619), .Z(DataO[19]) );
  BUFTD1 \DataO_tri[4]  ( .I(DataOr[4]), .OE(n621), .Z(DataO[4]) );
  BUFTD1 \DataO_tri[6]  ( .I(DataOr[6]), .OE(n621), .Z(DataO[6]) );
  BUFTD1 \DataO_tri[8]  ( .I(DataOr[8]), .OE(n621), .Z(DataO[8]) );
  BUFTD1 \DataO_tri[10]  ( .I(DataOr[10]), .OE(n619), .Z(DataO[10]) );
  BUFTD1 \DataO_tri[11]  ( .I(DataOr[11]), .OE(n619), .Z(DataO[11]) );
  BUFTD1 \DataO_tri[12]  ( .I(DataOr[12]), .OE(n619), .Z(DataO[12]) );
  BUFTD1 \DataO_tri[21]  ( .I(DataOr[21]), .OE(n620), .Z(DataO[21]) );
  BUFTD1 \DataO_tri[13]  ( .I(DataOr[13]), .OE(n619), .Z(DataO[13]) );
  BUFTD1 \DataO_tri[20]  ( .I(DataOr[20]), .OE(n620), .Z(DataO[20]) );
  BUFTD1 \DataO_tri[14]  ( .I(DataOr[14]), .OE(n619), .Z(DataO[14]) );
  BUFTD1 \DataO_tri[15]  ( .I(DataOr[15]), .OE(n619), .Z(DataO[15]) );
  BUFTD1 \DataO_tri[16]  ( .I(DataOr[16]), .OE(n619), .Z(DataO[16]) );
  BUFTD1 \DataO_tri[17]  ( .I(DataOr[17]), .OE(n619), .Z(DataO[17]) );
  BUFTD1 \DataO_tri[9]  ( .I(DataOr[9]), .OE(n621), .Z(DataO[9]) );
  BUFFD1 U4 ( .I(n108), .Z(n562) );
  BUFFD1 U5 ( .I(n591), .Z(n589) );
  BUFFD1 U6 ( .I(n562), .Z(n603) );
  BUFFD1 U7 ( .I(N45), .Z(n537) );
  BUFFD1 U8 ( .I(n537), .Z(n538) );
  BUFFD1 U9 ( .I(N46), .Z(n606) );
  BUFFD0 U10 ( .I(n596), .Z(n573) );
  BUFFD0 U11 ( .I(n596), .Z(n574) );
  BUFFD0 U12 ( .I(n596), .Z(n575) );
  BUFFD0 U13 ( .I(n597), .Z(n572) );
  BUFFD0 U14 ( .I(n597), .Z(n569) );
  BUFFD0 U15 ( .I(n597), .Z(n570) );
  BUFFD0 U16 ( .I(n598), .Z(n566) );
  BUFFD0 U17 ( .I(n598), .Z(n565) );
  BUFFD0 U23 ( .I(n593), .Z(n587) );
  BUFFD0 U24 ( .I(n594), .Z(n583) );
  BUFFD1 U25 ( .I(n600), .Z(n596) );
  BUFFD1 U26 ( .I(n564), .Z(n602) );
  CKND0 U29 ( .CLK(Reset), .CN(n108) );
  BUFFD0 U30 ( .I(n596), .Z(n563) );
  AN2D1 U31 ( .A1(n36), .A2(Dreadyr), .Z(Dready) );
  INVD1 U32 ( .I(n35), .ZN(n36) );
  BUFFD1 U37 ( .I(n47), .Z(n46) );
  NR2D3 U38 ( .A1(n66), .A2(n71), .ZN(n1) );
  NR2D3 U39 ( .A1(n69), .A2(n103), .ZN(n2) );
  NR2D3 U40 ( .A1(n99), .A2(n103), .ZN(n3) );
  NR2D3 U41 ( .A1(n98), .A2(n103), .ZN(n4) );
  NR2D3 U42 ( .A1(n71), .A2(n103), .ZN(n5) );
  NR2D3 U43 ( .A1(n69), .A2(n101), .ZN(n6) );
  NR2D3 U44 ( .A1(n99), .A2(n101), .ZN(n7) );
  NR2D3 U45 ( .A1(n98), .A2(n101), .ZN(n8) );
  NR2D3 U46 ( .A1(n71), .A2(n101), .ZN(n9) );
  NR2D3 U47 ( .A1(n69), .A2(n70), .ZN(n10) );
  NR2D3 U48 ( .A1(n70), .A2(n99), .ZN(n11) );
  NR2D3 U49 ( .A1(n70), .A2(n98), .ZN(n12) );
  NR2D3 U50 ( .A1(n70), .A2(n71), .ZN(n13) );
  NR2D3 U51 ( .A1(n68), .A2(n103), .ZN(n14) );
  NR2D3 U52 ( .A1(n67), .A2(n103), .ZN(n15) );
  NR2D3 U53 ( .A1(n85), .A2(n103), .ZN(n16) );
  NR2D3 U54 ( .A1(n72), .A2(n103), .ZN(n17) );
  NR2D3 U55 ( .A1(n68), .A2(n101), .ZN(n18) );
  NR2D3 U56 ( .A1(n67), .A2(n101), .ZN(n19) );
  NR2D3 U57 ( .A1(n85), .A2(n101), .ZN(n20) );
  NR2D3 U58 ( .A1(n72), .A2(n101), .ZN(n21) );
  NR2D3 U59 ( .A1(n68), .A2(n70), .ZN(n22) );
  NR2D3 U60 ( .A1(n67), .A2(n70), .ZN(n23) );
  NR2D3 U61 ( .A1(n70), .A2(n85), .ZN(n24) );
  NR2D3 U62 ( .A1(n70), .A2(n72), .ZN(n25) );
  NR2D3 U63 ( .A1(n66), .A2(n68), .ZN(n26) );
  NR2D3 U64 ( .A1(n66), .A2(n99), .ZN(n27) );
  NR2D3 U65 ( .A1(n66), .A2(n98), .ZN(n28) );
  NR2D3 U66 ( .A1(n66), .A2(n85), .ZN(n29) );
  NR2D3 U67 ( .A1(n66), .A2(n72), .ZN(n30) );
  NR2D3 U68 ( .A1(n66), .A2(n69), .ZN(n31) );
  NR2D3 U69 ( .A1(n66), .A2(n67), .ZN(n32) );
  CKBXD0 U70 ( .I(n40), .Z(n39) );
  CKBXD0 U71 ( .I(n41), .Z(n40) );
  CKBXD0 U72 ( .I(n42), .Z(n41) );
  CKNXD0 U73 ( .I(n625), .ZN(n624) );
  INVD6 U74 ( .I(n33), .ZN(n34) );
  INVD0 U75 ( .I(n37), .ZN(n33) );
  BUFFD16 U76 ( .I(n623), .Z(n37) );
  CKND1 U77 ( .CLK(n36), .CN(n623) );
  INVD2P5 U78 ( .I(n38), .ZN(n35) );
  CKBXD0 U79 ( .I(n39), .Z(n38) );
  CKBXD0 U80 ( .I(n43), .Z(n42) );
  INVD6 U82 ( .I(ChipEna), .ZN(n625) );
  BUFFD6 U83 ( .I(n44), .Z(n43) );
  CKBXD0 U84 ( .I(n45), .Z(n44) );
  BUFFD0 U85 ( .I(n46), .Z(n45) );
  CKBXD0 U86 ( .I(n48), .Z(n47) );
  BUFFD6 U87 ( .I(n49), .Z(n48) );
  CKBXD0 U88 ( .I(n50), .Z(n49) );
  BUFFD6 U89 ( .I(n51), .Z(n50) );
  CKBXD0 U90 ( .I(n52), .Z(n51) );
  BUFFD6 U91 ( .I(n53), .Z(n52) );
  CKBXD0 U92 ( .I(n54), .Z(n53) );
  BUFFD6 U93 ( .I(n55), .Z(n54) );
  CKBXD0 U94 ( .I(n624), .Z(n55) );
  INVD0 U95 ( .I(n622), .ZN(n621) );
  INVD1 U96 ( .I(N48), .ZN(n528) );
  INVD1 U97 ( .I(DataI[13]), .ZN(n614) );
  INVD1 U98 ( .I(DataI[14]), .ZN(n616) );
  INVD1 U99 ( .I(DataI[15]), .ZN(n618) );
  INVD1 U100 ( .I(DataI[5]), .ZN(n608) );
  INVD1 U101 ( .I(DataI[6]), .ZN(n610) );
  INVD1 U102 ( .I(DataI[7]), .ZN(n612) );
  BUFFD1 U103 ( .I(n592), .Z(n588) );
  BUFFD1 U104 ( .I(n598), .Z(n567) );
  BUFFD1 U105 ( .I(n598), .Z(n568) );
  BUFFD1 U106 ( .I(n597), .Z(n571) );
  BUFFD1 U107 ( .I(n595), .Z(n576) );
  BUFFD1 U108 ( .I(n595), .Z(n577) );
  BUFFD1 U109 ( .I(n595), .Z(n578) );
  BUFFD1 U110 ( .I(n595), .Z(n579) );
  BUFFD1 U111 ( .I(n594), .Z(n580) );
  BUFFD1 U112 ( .I(n594), .Z(n581) );
  BUFFD1 U113 ( .I(n594), .Z(n582) );
  BUFFD1 U114 ( .I(n593), .Z(n584) );
  BUFFD1 U115 ( .I(n593), .Z(n585) );
  BUFFD1 U116 ( .I(n593), .Z(n586) );
  BUFFD1 U117 ( .I(n562), .Z(n592) );
  BUFFD1 U118 ( .I(n591), .Z(n590) );
  BUFFD1 U119 ( .I(n599), .Z(n597) );
  BUFFD1 U120 ( .I(n600), .Z(n595) );
  BUFFD1 U121 ( .I(n601), .Z(n594) );
  BUFFD1 U122 ( .I(n601), .Z(n593) );
  BUFFD1 U123 ( .I(n599), .Z(n598) );
  BUFFD1 U124 ( .I(n555), .Z(n551) );
  BUFFD1 U125 ( .I(n554), .Z(n550) );
  BUFFD1 U126 ( .I(n555), .Z(n552) );
  BUFFD1 U127 ( .I(n549), .Z(n553) );
  BUFFD1 U128 ( .I(n549), .Z(n554) );
  BUFFD1 U129 ( .I(n549), .Z(n555) );
  BUFFD1 U130 ( .I(n548), .Z(n556) );
  BUFFD1 U131 ( .I(n548), .Z(n557) );
  BUFFD1 U132 ( .I(n548), .Z(n558) );
  BUFFD1 U133 ( .I(n538), .Z(n544) );
  BUFFD1 U134 ( .I(n538), .Z(n545) );
  BUFFD1 U135 ( .I(n539), .Z(n541) );
  BUFFD1 U136 ( .I(n539), .Z(n542) );
  BUFFD1 U137 ( .I(n540), .Z(n543) );
  BUFFD1 U138 ( .I(n561), .Z(n600) );
  BUFFD1 U139 ( .I(n561), .Z(n601) );
  BUFFD1 U140 ( .I(n561), .Z(n599) );
  BUFFD1 U141 ( .I(n604), .Z(n591) );
  BUFFD1 U142 ( .I(n563), .Z(n604) );
  INVD1 U143 ( .I(n34), .ZN(n620) );
  INVD1 U144 ( .I(n34), .ZN(n619) );
  XOR3D1 U145 ( .A1(N60), .A2(N59), .A3(n95), .Z(n94) );
  XOR3D1 U146 ( .A1(n96), .A2(N58), .A3(n97), .Z(n95) );
  XOR3D1 U147 ( .A1(N79), .A2(N74), .A3(n86), .Z(N83) );
  XOR3D1 U148 ( .A1(N73), .A2(n87), .A3(n88), .Z(n86) );
  XOR3D1 U149 ( .A1(N77), .A2(N76), .A3(n89), .Z(n88) );
  XOR3D1 U150 ( .A1(N67), .A2(N66), .A3(n92), .Z(n90) );
  XOR3D1 U151 ( .A1(N65), .A2(n93), .A3(n94), .Z(n92) );
  BUFFD1 U152 ( .I(n538), .Z(n540) );
  BUFFD1 U153 ( .I(n547), .Z(n559) );
  BUFFD1 U154 ( .I(n546), .Z(n547) );
  BUFFD1 U155 ( .I(n530), .Z(n531) );
  BUFFD1 U156 ( .I(n533), .Z(n536) );
  BUFFD1 U157 ( .I(n536), .Z(n534) );
  BUFFD1 U158 ( .I(n533), .Z(n535) );
  BUFFD1 U159 ( .I(n532), .Z(n530) );
  BUFFD1 U160 ( .I(n546), .Z(n549) );
  BUFFD1 U161 ( .I(n546), .Z(n548) );
  BUFFD1 U162 ( .I(n538), .Z(n539) );
  ND3D1 U163 ( .A1(n106), .A2(n105), .A3(n104), .ZN(n69) );
  XOR3D1 U164 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n73), .Z(N85) );
  XOR3D1 U165 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n73), .Z(n560) );
  XOR3D1 U166 ( .A1(n83), .A2(DataI[17]), .A3(n84), .Z(n82) );
  XOR3D1 U167 ( .A1(DataI[0]), .A2(n74), .A3(n75), .Z(n73) );
  XOR3D1 U168 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n76), .Z(n75) );
  XOR3D1 U169 ( .A1(n77), .A2(DataI[3]), .A3(n78), .Z(n76) );
  XOR3D1 U170 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n79), .Z(n78) );
  XOR3D1 U171 ( .A1(n80), .A2(DataI[10]), .A3(n81), .Z(n79) );
  XOR3D1 U172 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n82), .Z(n81) );
  BUFFD1 U173 ( .I(Read), .Z(n605) );
  BUFFD1 U174 ( .I(n564), .Z(n561) );
  BUFFD1 U175 ( .I(n108), .Z(n564) );
  INVD1 U176 ( .I(n36), .ZN(n622) );
  BUFFD1 U177 ( .I(N47), .Z(n532) );
  BUFFD1 U178 ( .I(N44), .Z(n546) );
  BUFFD1 U179 ( .I(n606), .Z(n533) );
  INVD1 U180 ( .I(n528), .ZN(n529) );
  ND3D1 U181 ( .A1(n100), .A2(n102), .A3(Write), .ZN(n103) );
  ND3D1 U182 ( .A1(AddrW[3]), .A2(n102), .A3(Write), .ZN(n101) );
  ND3D1 U183 ( .A1(AddrW[4]), .A2(n100), .A3(Write), .ZN(n70) );
  ND3D1 U184 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n66) );
  ND3D1 U185 ( .A1(AddrW[0]), .A2(n106), .A3(AddrW[2]), .ZN(n85) );
  ND3D1 U186 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n71) );
  ND3D1 U187 ( .A1(AddrW[1]), .A2(n105), .A3(AddrW[0]), .ZN(n99) );
  ND3D1 U188 ( .A1(AddrW[1]), .A2(n104), .A3(AddrW[2]), .ZN(n72) );
  ND3D1 U189 ( .A1(n104), .A2(n106), .A3(AddrW[2]), .ZN(n98) );
  ND3D1 U190 ( .A1(n106), .A2(n105), .A3(AddrW[0]), .ZN(n68) );
  ND3D1 U191 ( .A1(n104), .A2(n105), .A3(AddrW[1]), .ZN(n67) );
  INVD1 U192 ( .I(AddrW[2]), .ZN(n105) );
  INVD1 U193 ( .I(AddrW[0]), .ZN(n104) );
  INVD1 U194 ( .I(AddrW[1]), .ZN(n106) );
  INVD1 U195 ( .I(AddrW[4]), .ZN(n102) );
  INVD1 U196 ( .I(AddrW[3]), .ZN(n100) );
  INVD1 U197 ( .I(n612), .ZN(n611) );
  INVD1 U198 ( .I(n616), .ZN(n615) );
  INVD1 U199 ( .I(n618), .ZN(n617) );
  INVD1 U200 ( .I(n614), .ZN(n613) );
  INVD1 U201 ( .I(n608), .ZN(n607) );
  INVD1 U202 ( .I(n610), .ZN(n609) );
  MUX4ND0 U203 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n553), .S1(n540), .ZN(
        n440) );
  MUX4ND0 U204 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n554), .S1(n540), .ZN(
        n466) );
  MUX4ND0 U205 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n547), .S1(n539), .ZN(
        n492) );
  MUX4ND0 U206 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n555), .S1(n539), .ZN(
        n505) );
  MUX4D0 U207 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n559), .S1(n543), .Z(
        n428) );
  MUX4D0 U208 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n557), .S1(n540), .Z(
        n441) );
  MUX4D0 U209 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n549), .S1(n540), .Z(
        n454) );
  MUX4D0 U210 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n558), .S1(n543), .Z(
        n467) );
  MUX4D0 U211 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n550), .S1(n540), .Z(
        n432) );
  MUX4D0 U212 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n550), .S1(n540), .Z(
        n430) );
  MUX4D0 U213 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n553), .S1(n543), .Z(
        n445) );
  MUX4D0 U214 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n549), .S1(n537), .Z(
        n443) );
  MUX4D0 U215 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n549), .S1(n540), .Z(
        n458) );
  MUX4D0 U216 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n549), .S1(n540), .Z(
        n456) );
  MUX4D0 U217 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n559), .S1(n543), .Z(
        n471) );
  MUX4D0 U218 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n557), .S1(n543), .Z(
        n469) );
  MUX4D0 U219 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n559), .S1(n542), .Z(
        n484) );
  MUX4D0 U220 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n555), .S1(n543), .Z(
        n497) );
  MUX4D0 U221 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n556), .S1(n543), .Z(
        n510) );
  MUX4D0 U222 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n555), .S1(n543), .Z(
        n429) );
  MUX4D0 U223 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n558), .S1(n540), .Z(
        n442) );
  MUX4D0 U224 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n549), .S1(n540), .Z(
        n455) );
  MUX4D0 U225 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n553), .S1(n541), .Z(
        n468) );
  MUX4D0 U226 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n552), .S1(n543), .Z(
        n433) );
  MUX4D0 U227 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n556), .S1(n545), .Z(
        n431) );
  MUX4D0 U228 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n555), .S1(n540), .Z(
        n446) );
  MUX4D0 U229 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n549), .S1(n540), .Z(
        n444) );
  MUX4D0 U230 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n554), .S1(n537), .Z(
        n459) );
  MUX4D0 U231 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n553), .S1(n537), .Z(
        n457) );
  MUX4D0 U232 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n556), .S1(n543), .Z(
        n472) );
  MUX4D0 U233 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n558), .S1(n543), .Z(
        n470) );
  MUX4D0 U234 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n547), .S1(n543), .Z(
        n485) );
  MUX4D0 U235 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n551), .S1(n543), .Z(
        n498) );
  MUX4D0 U236 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n555), .S1(n543), .Z(
        n496) );
  MUX4D0 U237 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n555), .S1(n543), .Z(
        n511) );
  MUX4ND0 U238 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n554), .S1(n539), .ZN(
        n518) );
  MUX4ND0 U239 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n557), .S1(n540), .ZN(
        n427) );
  MUX4ND0 U240 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n550), .S1(n540), .ZN(
        n453) );
  MUX4ND0 U241 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n553), .S1(n539), .ZN(
        n479) );
  MUX4ND0 U242 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n548), .S1(n537), .ZN(
        n128) );
  MUX4ND0 U243 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n559), .S1(n538), .ZN(
        n141) );
  MUX4ND0 U244 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n546), .S1(n537), .ZN(
        n154) );
  MUX4ND0 U245 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n546), .S1(n538), .ZN(
        n167) );
  MUX4ND0 U246 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n548), .S1(n543), .ZN(
        n180) );
  MUX4ND0 U247 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n554), .S1(n537), .ZN(
        n193) );
  MUX4ND0 U248 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n549), .S1(n538), .ZN(
        n206) );
  MUX4ND0 U249 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n556), .S1(n537), .ZN(
        n232) );
  MUX4ND0 U250 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n548), .S1(n537), .ZN(
        n245) );
  MUX4ND0 U251 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n556), .S1(n537), .ZN(
        n258) );
  MUX4ND0 U252 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n546), .S1(n537), .ZN(
        n271) );
  MUX4ND0 U253 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n558), .S1(n537), .ZN(
        n284) );
  MUX4ND0 U254 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n558), .S1(n537), .ZN(
        n297) );
  MUX4ND0 U255 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n557), .S1(n540), .ZN(
        n310) );
  MUX4ND0 U256 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n546), .S1(n540), .ZN(
        n323) );
  MUX4ND0 U257 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n559), .S1(n540), .ZN(
        n336) );
  MUX4ND0 U258 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n556), .S1(n540), .ZN(
        n349) );
  MUX4ND0 U259 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n553), .S1(n538), .ZN(
        n219) );
  MUX4ND0 U260 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n549), .S1(n537), .ZN(
        n59) );
  MUX4ND0 U261 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n546), .S1(n537), .ZN(
        n115) );
  MUX4D0 U262 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n549), .S1(n543), .Z(
        n519) );
  MUX4D0 U263 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n553), .S1(n537), .Z(n60) );
  MUX4D0 U264 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n546), .S1(n544), .Z(
        n116) );
  MUX4D0 U265 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n556), .S1(n545), .Z(
        n129) );
  MUX4D0 U266 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n548), .S1(n545), .Z(
        n142) );
  MUX4D0 U267 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n548), .S1(n537), .Z(
        n155) );
  MUX4D0 U268 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n546), .S1(n537), .Z(
        n168) );
  MUX4D0 U269 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n546), .S1(n540), .Z(
        n181) );
  MUX4D0 U270 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n554), .S1(n545), .Z(
        n194) );
  MUX4D0 U271 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(N44), .S1(n538), .Z(n207) );
  MUX4D0 U272 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n548), .S1(n537), .Z(
        n220) );
  MUX4D0 U273 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n553), .S1(n545), .Z(
        n233) );
  MUX4D0 U274 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n553), .S1(n539), .Z(
        n246) );
  MUX4D0 U275 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n553), .S1(n544), .Z(
        n259) );
  MUX4D0 U276 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n554), .S1(n544), .Z(
        n272) );
  MUX4D0 U277 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n554), .S1(n544), .Z(
        n285) );
  MUX4D0 U278 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n555), .S1(n539), .Z(
        n298) );
  MUX4D0 U279 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n555), .S1(n539), .Z(
        n311) );
  MUX4D0 U280 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n556), .S1(n541), .Z(
        n324) );
  MUX4D0 U281 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n556), .S1(N45), .Z(
        n337) );
  MUX4D0 U282 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n557), .S1(N45), .Z(
        n350) );
  MUX4D0 U283 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n557), .S1(n541), .Z(
        n363) );
  MUX4D0 U284 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n558), .S1(n541), .Z(
        n376) );
  MUX4D0 U285 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n558), .S1(n542), .Z(
        n389) );
  MUX4D0 U286 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n559), .S1(n542), .Z(
        n402) );
  MUX4D0 U287 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n559), .S1(n543), .Z(
        n415) );
  MUX4D0 U288 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n556), .S1(n543), .Z(
        n480) );
  MUX4D0 U289 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n547), .S1(n540), .Z(
        n493) );
  MUX4D0 U290 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n546), .S1(n543), .Z(
        n506) );
  MUX4D0 U291 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n558), .S1(n544), .Z(
        n523) );
  MUX4D0 U292 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n547), .S1(n544), .Z(
        n521) );
  MUX4D0 U293 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n555), .S1(n544), .Z(n64)
         );
  MUX4D0 U294 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n557), .S1(n544), .Z(n62) );
  MUX4D0 U295 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n547), .S1(n545), .Z(n120)
         );
  MUX4D0 U296 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n550), .S1(n544), .Z(
        n118) );
  MUX4D0 U297 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(N44), .S1(n545), .Z(n133)
         );
  MUX4D0 U298 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n547), .S1(n545), .Z(
        n131) );
  MUX4D0 U299 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n548), .S1(n545), .Z(n146)
         );
  MUX4D0 U300 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n548), .S1(n545), .Z(
        n144) );
  MUX4D0 U301 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n559), .S1(n539), .Z(n159)
         );
  MUX4D0 U302 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n547), .S1(n537), .Z(
        n157) );
  MUX4D0 U303 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(N44), .S1(n537), .Z(n172)
         );
  MUX4D0 U304 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n546), .S1(n538), .Z(
        n170) );
  MUX4D0 U305 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(N44), .S1(n545), .Z(n185)
         );
  MUX4D0 U306 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(N44), .S1(n545), .Z(n183) );
  MUX4D0 U307 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n559), .S1(n545), .Z(n198)
         );
  MUX4D0 U308 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n548), .S1(n545), .Z(
        n196) );
  MUX4D0 U309 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n551), .S1(n545), .Z(n211)
         );
  MUX4D0 U310 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n546), .S1(n545), .Z(
        n209) );
  MUX4D0 U311 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n548), .S1(n545), .Z(n224)
         );
  MUX4D0 U312 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n548), .S1(n537), .Z(
        n222) );
  MUX4D0 U313 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n548), .S1(n541), .Z(
        n237) );
  MUX4D0 U314 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n547), .S1(n542), .Z(
        n235) );
  MUX4D0 U315 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n553), .S1(n539), .Z(
        n250) );
  MUX4D0 U316 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n553), .S1(n539), .Z(
        n248) );
  MUX4D0 U317 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n553), .S1(n544), .Z(
        n263) );
  MUX4D0 U318 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n553), .S1(n544), .Z(
        n261) );
  MUX4D0 U319 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n554), .S1(n542), .Z(
        n276) );
  MUX4D0 U320 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n554), .S1(n544), .Z(
        n274) );
  MUX4D0 U321 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n554), .S1(n544), .Z(
        n289) );
  MUX4D0 U322 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n554), .S1(n544), .Z(
        n287) );
  MUX4D0 U323 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n555), .S1(n542), .Z(
        n302) );
  MUX4D0 U324 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n555), .S1(n539), .Z(
        n300) );
  MUX4D0 U325 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n555), .S1(n541), .Z(
        n315) );
  MUX4D0 U326 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n555), .S1(n543), .Z(
        n313) );
  MUX4D0 U327 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n556), .S1(n544), .Z(
        n328) );
  MUX4D0 U328 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n556), .S1(n542), .Z(
        n326) );
  MUX4D0 U329 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n556), .S1(n538), .Z(
        n341) );
  MUX4D0 U330 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n556), .S1(N45), .Z(
        n339) );
  MUX4D0 U331 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n557), .S1(n541), .Z(
        n354) );
  MUX4D0 U332 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n557), .S1(N45), .Z(
        n352) );
  MUX4D0 U333 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n557), .S1(n541), .Z(
        n367) );
  MUX4D0 U334 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n557), .S1(n541), .Z(
        n365) );
  MUX4D0 U335 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n558), .S1(n542), .Z(
        n380) );
  MUX4D0 U336 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n558), .S1(n541), .Z(
        n378) );
  MUX4D0 U337 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n558), .S1(n542), .Z(
        n393) );
  MUX4D0 U338 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n558), .S1(n542), .Z(
        n391) );
  MUX4D0 U339 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n559), .S1(n542), .Z(
        n406) );
  MUX4D0 U340 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n559), .S1(n542), .Z(
        n404) );
  MUX4D0 U341 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n558), .S1(n544), .Z(
        n419) );
  MUX4D0 U342 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n559), .S1(n540), .Z(
        n417) );
  MUX4D0 U343 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n553), .S1(n540), .Z(
        n482) );
  MUX4D0 U344 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n547), .S1(n543), .Z(
        n495) );
  MUX4D0 U345 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n557), .S1(n543), .Z(
        n508) );
  MUX4D0 U346 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n549), .S1(n543), .Z(
        n520) );
  MUX4D0 U347 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n559), .S1(n544), .Z(n61) );
  MUX4D0 U348 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n557), .S1(n544), .Z(
        n117) );
  MUX4D0 U349 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n550), .S1(n545), .Z(
        n130) );
  MUX4D0 U350 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n547), .S1(n545), .Z(
        n143) );
  MUX4D0 U351 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n548), .S1(n537), .Z(
        n156) );
  MUX4D0 U352 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n546), .S1(n538), .Z(
        n169) );
  MUX4D0 U353 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(N44), .S1(n538), .Z(n182) );
  MUX4D0 U354 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n554), .S1(n545), .Z(
        n195) );
  MUX4D0 U355 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n546), .S1(N45), .Z(n208) );
  MUX4D0 U356 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n559), .S1(n545), .Z(
        n221) );
  MUX4D0 U357 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n548), .S1(n541), .Z(
        n234) );
  MUX4D0 U358 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n553), .S1(n539), .Z(
        n247) );
  MUX4D0 U359 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n553), .S1(n539), .Z(
        n260) );
  MUX4D0 U360 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n554), .S1(n544), .Z(
        n273) );
  MUX4D0 U361 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n554), .S1(n539), .Z(
        n286) );
  MUX4D0 U362 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n555), .S1(n542), .Z(
        n299) );
  MUX4D0 U363 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n555), .S1(n539), .Z(
        n312) );
  MUX4D0 U364 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n556), .S1(n542), .Z(
        n325) );
  MUX4D0 U365 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n556), .S1(N45), .Z(
        n338) );
  MUX4D0 U366 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n557), .S1(n537), .Z(
        n351) );
  MUX4D0 U367 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n557), .S1(n541), .Z(
        n364) );
  MUX4D0 U368 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n558), .S1(n541), .Z(
        n377) );
  MUX4D0 U369 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n558), .S1(n542), .Z(
        n390) );
  MUX4D0 U370 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n559), .S1(n542), .Z(
        n403) );
  MUX4D0 U371 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n559), .S1(n543), .Z(
        n416) );
  MUX4D0 U372 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n557), .S1(n543), .Z(
        n481) );
  MUX4D0 U373 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n549), .S1(n543), .Z(
        n494) );
  MUX4D0 U374 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n558), .S1(n543), .Z(
        n507) );
  MUX4D0 U375 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n549), .S1(n544), .Z(
        n524) );
  MUX4D0 U376 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n556), .S1(n544), .Z(
        n522) );
  MUX4D0 U377 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n558), .S1(n544), .Z(n65)
         );
  MUX4D0 U378 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n550), .S1(n544), .Z(n63) );
  MUX4D0 U379 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n550), .S1(n545), .Z(n121)
         );
  MUX4D0 U380 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n547), .S1(n544), .Z(
        n119) );
  MUX4D0 U381 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n547), .S1(n545), .Z(n134)
         );
  MUX4D0 U382 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n552), .S1(n545), .Z(
        n132) );
  MUX4D0 U383 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n547), .S1(n538), .Z(n147)
         );
  MUX4D0 U384 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n547), .S1(n545), .Z(
        n145) );
  MUX4D0 U385 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n548), .S1(n542), .Z(n160)
         );
  MUX4D0 U386 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n547), .S1(n541), .Z(
        n158) );
  MUX4D0 U387 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(N44), .S1(n538), .Z(n173)
         );
  MUX4D0 U388 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n546), .S1(n538), .Z(
        n171) );
  MUX4D0 U389 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(N44), .S1(n545), .Z(n186)
         );
  MUX4D0 U390 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(N44), .S1(n538), .Z(n184) );
  MUX4D0 U391 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n548), .S1(n545), .Z(n199)
         );
  MUX4D0 U392 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n548), .S1(n545), .Z(
        n197) );
  MUX4D0 U393 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n554), .S1(n545), .Z(n212)
         );
  MUX4D0 U394 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n549), .S1(n545), .Z(
        n210) );
  MUX4D0 U395 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n547), .S1(n538), .Z(n225)
         );
  MUX4D0 U396 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n547), .S1(n545), .Z(
        n223) );
  MUX4D0 U397 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n547), .S1(n542), .Z(
        n238) );
  MUX4D0 U398 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n553), .S1(N45), .Z(
        n236) );
  MUX4D0 U399 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n553), .S1(n539), .Z(
        n251) );
  MUX4D0 U400 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n553), .S1(n539), .Z(
        n249) );
  MUX4D0 U401 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n554), .S1(n544), .Z(
        n264) );
  MUX4D0 U402 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n553), .S1(n544), .Z(
        n262) );
  MUX4D0 U403 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n554), .S1(n544), .Z(
        n277) );
  MUX4D0 U404 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n554), .S1(n542), .Z(
        n275) );
  MUX4D0 U405 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n555), .S1(n541), .Z(
        n290) );
  MUX4D0 U406 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n554), .S1(n541), .Z(
        n288) );
  MUX4D0 U407 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n555), .S1(n542), .Z(
        n303) );
  MUX4D0 U408 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n555), .S1(n541), .Z(
        n301) );
  MUX4D0 U409 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n556), .S1(n544), .Z(
        n316) );
  MUX4D0 U410 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n555), .S1(n541), .Z(
        n314) );
  MUX4D0 U411 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n556), .S1(N45), .Z(n329) );
  MUX4D0 U412 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n556), .S1(N45), .Z(
        n327) );
  MUX4D0 U413 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n557), .S1(n543), .Z(
        n342) );
  MUX4D0 U414 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n556), .S1(N45), .Z(
        n340) );
  MUX4D0 U415 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n557), .S1(n541), .Z(
        n355) );
  MUX4D0 U416 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n557), .S1(n541), .Z(
        n353) );
  MUX4D0 U417 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n558), .S1(n541), .Z(
        n368) );
  MUX4D0 U418 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n557), .S1(n541), .Z(
        n366) );
  MUX4D0 U419 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n558), .S1(n542), .Z(
        n381) );
  MUX4D0 U420 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n558), .S1(n541), .Z(
        n379) );
  MUX4D0 U421 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n559), .S1(n542), .Z(
        n394) );
  MUX4D0 U422 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n558), .S1(n542), .Z(
        n392) );
  MUX4D0 U423 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n559), .S1(n540), .Z(
        n407) );
  MUX4D0 U424 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n559), .S1(n542), .Z(
        n405) );
  MUX4D0 U425 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n546), .S1(n540), .Z(
        n420) );
  MUX4D0 U426 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n559), .S1(n540), .Z(
        n418) );
  MUX4D0 U427 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n548), .S1(n543), .Z(
        n483) );
  MUX4D0 U428 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n559), .S1(n543), .Z(
        n509) );
  MUX4ND0 U429 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n549), .S1(n540), .ZN(
        n362) );
  MUX4ND0 U430 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n548), .S1(n540), .ZN(
        n375) );
  MUX4ND0 U431 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n546), .S1(n540), .ZN(
        n388) );
  MUX4ND0 U432 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n547), .S1(n540), .ZN(
        n401) );
  MUX4ND0 U433 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n557), .S1(n540), .ZN(
        n414) );
  AN2D1 U434 ( .A1(ClkR), .A2(n621), .Z(ClockR) );
  MUX3ND0 U435 ( .I0(n57), .I1(n58), .I2(n59), .S0(n539), .S1(n533), .ZN(n56)
         );
  MUX3ND0 U436 ( .I0(n109), .I1(n110), .I2(n111), .S0(n532), .S1(n529), .ZN(
        N82) );
  MUX3ND0 U437 ( .I0(n113), .I1(n114), .I2(n115), .S0(n538), .S1(n606), .ZN(
        n112) );
  MUX3ND0 U438 ( .I0(n122), .I1(n123), .I2(n124), .S0(n530), .S1(n529), .ZN(
        N81) );
  MUX3ND0 U439 ( .I0(n126), .I1(n127), .I2(n128), .S0(n539), .S1(n534), .ZN(
        n125) );
  MUX3ND0 U440 ( .I0(n135), .I1(n136), .I2(n137), .S0(n531), .S1(n529), .ZN(
        N80) );
  MUX3ND0 U441 ( .I0(n139), .I1(n140), .I2(n141), .S0(n542), .S1(n534), .ZN(
        n138) );
  MUX3ND0 U442 ( .I0(n148), .I1(n149), .I2(n150), .S0(N47), .S1(n529), .ZN(N79) );
  MUX3ND0 U443 ( .I0(n152), .I1(n153), .I2(n154), .S0(n537), .S1(n534), .ZN(
        n151) );
  MUX3ND0 U444 ( .I0(n161), .I1(n162), .I2(n163), .S0(n532), .S1(n529), .ZN(
        N78) );
  MUX3ND0 U445 ( .I0(n165), .I1(n166), .I2(n167), .S0(n544), .S1(n534), .ZN(
        n164) );
  MUX3ND0 U446 ( .I0(n174), .I1(n175), .I2(n176), .S0(n532), .S1(n529), .ZN(
        N77) );
  MUX3ND0 U447 ( .I0(n178), .I1(n179), .I2(n180), .S0(n541), .S1(n534), .ZN(
        n177) );
  MUX3ND0 U448 ( .I0(n187), .I1(n188), .I2(n189), .S0(n530), .S1(n529), .ZN(
        N76) );
  MUX3ND0 U449 ( .I0(n191), .I1(n192), .I2(n193), .S0(n542), .S1(n534), .ZN(
        n190) );
  MUX3ND0 U450 ( .I0(n200), .I1(n201), .I2(n202), .S0(n530), .S1(n529), .ZN(
        N75) );
  MUX3ND0 U451 ( .I0(n204), .I1(n205), .I2(n206), .S0(N45), .S1(n534), .ZN(
        n203) );
  MUX3ND0 U452 ( .I0(n213), .I1(n214), .I2(n215), .S0(N47), .S1(n529), .ZN(N74) );
  MUX3ND0 U453 ( .I0(n217), .I1(n218), .I2(n219), .S0(n539), .S1(n534), .ZN(
        n216) );
  MUX3ND0 U454 ( .I0(n226), .I1(n227), .I2(n228), .S0(N47), .S1(n529), .ZN(N73) );
  MUX3ND0 U455 ( .I0(n230), .I1(n231), .I2(n232), .S0(n539), .S1(n534), .ZN(
        n229) );
  MUX3ND0 U456 ( .I0(n239), .I1(n240), .I2(n241), .S0(n530), .S1(n529), .ZN(
        N72) );
  MUX3ND0 U457 ( .I0(n243), .I1(n244), .I2(n245), .S0(n539), .S1(n534), .ZN(
        n242) );
  MUX3ND0 U458 ( .I0(n252), .I1(n253), .I2(n254), .S0(n530), .S1(n529), .ZN(
        N71) );
  MUX3ND0 U459 ( .I0(n256), .I1(n257), .I2(n258), .S0(n541), .S1(n534), .ZN(
        n255) );
  MUX3ND0 U460 ( .I0(n265), .I1(n266), .I2(n267), .S0(n530), .S1(n529), .ZN(
        N70) );
  MUX3ND0 U461 ( .I0(n269), .I1(n270), .I2(n271), .S0(N45), .S1(n534), .ZN(
        n268) );
  MUX3ND0 U462 ( .I0(n278), .I1(n279), .I2(n280), .S0(n531), .S1(n529), .ZN(
        N69) );
  MUX3ND0 U463 ( .I0(n282), .I1(n283), .I2(n284), .S0(n542), .S1(n534), .ZN(
        n281) );
  MUX3ND0 U464 ( .I0(n291), .I1(n292), .I2(n293), .S0(n531), .S1(n529), .ZN(
        N68) );
  MUX3ND0 U465 ( .I0(n295), .I1(n296), .I2(n297), .S0(n541), .S1(n535), .ZN(
        n294) );
  MUX3ND0 U466 ( .I0(n304), .I1(n305), .I2(n306), .S0(n531), .S1(n529), .ZN(
        N67) );
  MUX3ND0 U467 ( .I0(n308), .I1(n309), .I2(n310), .S0(n539), .S1(n535), .ZN(
        n307) );
  MUX3ND0 U468 ( .I0(n317), .I1(n318), .I2(n319), .S0(n531), .S1(n529), .ZN(
        N66) );
  MUX3ND0 U469 ( .I0(n321), .I1(n322), .I2(n323), .S0(n537), .S1(n535), .ZN(
        n320) );
  MUX3ND0 U470 ( .I0(n330), .I1(n331), .I2(n332), .S0(n531), .S1(n529), .ZN(
        N65) );
  MUX3ND0 U471 ( .I0(n334), .I1(n335), .I2(n336), .S0(n541), .S1(n535), .ZN(
        n333) );
  MUX3ND0 U472 ( .I0(n343), .I1(n344), .I2(n345), .S0(n531), .S1(n529), .ZN(
        N64) );
  MUX3ND0 U473 ( .I0(n347), .I1(n348), .I2(n349), .S0(n542), .S1(n535), .ZN(
        n346) );
  MUX3ND0 U474 ( .I0(n356), .I1(n357), .I2(n358), .S0(n531), .S1(n529), .ZN(
        N63) );
  MUX3ND0 U475 ( .I0(n360), .I1(n361), .I2(n362), .S0(n541), .S1(n535), .ZN(
        n359) );
  MUX3ND0 U476 ( .I0(n369), .I1(n370), .I2(n371), .S0(n531), .S1(N48), .ZN(N62) );
  MUX3ND0 U477 ( .I0(n373), .I1(n374), .I2(n375), .S0(n537), .S1(n535), .ZN(
        n372) );
  MUX3ND0 U478 ( .I0(n382), .I1(n383), .I2(n384), .S0(n531), .S1(N48), .ZN(N61) );
  MUX3ND0 U479 ( .I0(n386), .I1(n387), .I2(n388), .S0(n541), .S1(n535), .ZN(
        n385) );
  MUX3ND0 U480 ( .I0(n395), .I1(n396), .I2(n397), .S0(n531), .S1(n529), .ZN(
        N60) );
  MUX3ND0 U481 ( .I0(n399), .I1(n400), .I2(n401), .S0(n539), .S1(n535), .ZN(
        n398) );
  MUX3ND0 U482 ( .I0(n408), .I1(n409), .I2(n410), .S0(n531), .S1(n529), .ZN(
        N59) );
  MUX3ND0 U483 ( .I0(n412), .I1(n413), .I2(n414), .S0(n539), .S1(n535), .ZN(
        n411) );
  MUX3ND0 U484 ( .I0(n421), .I1(n422), .I2(n423), .S0(n531), .S1(N48), .ZN(N58) );
  MUX3ND0 U485 ( .I0(n425), .I1(n426), .I2(n427), .S0(n542), .S1(n535), .ZN(
        n424) );
  MUX3ND0 U486 ( .I0(n434), .I1(n435), .I2(n436), .S0(n531), .S1(N48), .ZN(N57) );
  MUX3ND0 U487 ( .I0(n438), .I1(n439), .I2(n440), .S0(n539), .S1(n535), .ZN(
        n437) );
  MUX3ND0 U488 ( .I0(n447), .I1(n448), .I2(n449), .S0(n532), .S1(N48), .ZN(N56) );
  MUX3ND0 U489 ( .I0(n451), .I1(n452), .I2(n453), .S0(n544), .S1(n535), .ZN(
        n450) );
  MUX3ND0 U490 ( .I0(n460), .I1(n461), .I2(n462), .S0(N47), .S1(N48), .ZN(N55)
         );
  MUX3ND0 U491 ( .I0(n464), .I1(n465), .I2(n466), .S0(n541), .S1(n606), .ZN(
        n463) );
  MUX3ND0 U492 ( .I0(n473), .I1(n474), .I2(n475), .S0(N47), .S1(N48), .ZN(N54)
         );
  MUX3ND0 U493 ( .I0(n477), .I1(n478), .I2(n479), .S0(n539), .S1(n606), .ZN(
        n476) );
  MUX3ND0 U494 ( .I0(n486), .I1(n487), .I2(n488), .S0(n532), .S1(N48), .ZN(N53) );
  MUX3ND0 U495 ( .I0(n490), .I1(n491), .I2(n492), .S0(n537), .S1(n606), .ZN(
        n489) );
  MUX3ND0 U496 ( .I0(n499), .I1(n500), .I2(n501), .S0(N47), .S1(N48), .ZN(N52)
         );
  MUX3ND0 U497 ( .I0(n503), .I1(n504), .I2(n505), .S0(n542), .S1(n606), .ZN(
        n502) );
  MUX3ND0 U498 ( .I0(n512), .I1(n513), .I2(n514), .S0(N47), .S1(N48), .ZN(N51)
         );
  MUX3ND0 U499 ( .I0(n516), .I1(n517), .I2(n518), .S0(n537), .S1(n533), .ZN(
        n515) );
  MUX3ND0 U500 ( .I0(n525), .I1(n526), .I2(n527), .S0(n532), .S1(N48), .ZN(N50) );
  MUX2ND0 U501 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n550), .ZN(
        n58) );
  MUX2ND0 U502 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n550), .ZN(
        n57) );
  MUX3ND0 U503 ( .I0(n61), .I1(n60), .I2(n56), .S0(n536), .S1(n532), .ZN(n111)
         );
  MUX2ND0 U504 ( .I0(n63), .I1(n62), .S(n606), .ZN(n110) );
  MUX2ND0 U505 ( .I0(n65), .I1(n64), .S(n533), .ZN(n109) );
  MUX2ND0 U506 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n550), .ZN(
        n114) );
  MUX2ND0 U507 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n550), .ZN(
        n113) );
  MUX3ND0 U508 ( .I0(n117), .I1(n116), .I2(n112), .S0(n536), .S1(n532), .ZN(
        n124) );
  MUX2ND0 U509 ( .I0(n119), .I1(n118), .S(n533), .ZN(n123) );
  MUX2ND0 U510 ( .I0(n121), .I1(n120), .S(n535), .ZN(n122) );
  MUX2ND0 U511 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n550), .ZN(
        n127) );
  MUX2ND0 U512 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n551), .ZN(
        n126) );
  MUX3ND0 U513 ( .I0(n130), .I1(n129), .I2(n125), .S0(n536), .S1(n532), .ZN(
        n137) );
  MUX2ND0 U514 ( .I0(n132), .I1(n131), .S(n536), .ZN(n136) );
  MUX2ND0 U515 ( .I0(n134), .I1(n133), .S(n536), .ZN(n135) );
  MUX2ND0 U516 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n551), .ZN(
        n140) );
  MUX2ND0 U517 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n551), .ZN(
        n139) );
  MUX3ND0 U518 ( .I0(n143), .I1(n142), .I2(n138), .S0(n536), .S1(n531), .ZN(
        n150) );
  MUX2ND0 U519 ( .I0(n145), .I1(n144), .S(n606), .ZN(n149) );
  MUX2ND0 U520 ( .I0(n147), .I1(n146), .S(n606), .ZN(n148) );
  MUX2ND0 U521 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n551), .ZN(
        n153) );
  MUX2ND0 U522 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n551), .ZN(
        n152) );
  MUX3ND0 U523 ( .I0(n156), .I1(n155), .I2(n151), .S0(n536), .S1(n532), .ZN(
        n163) );
  MUX2ND0 U524 ( .I0(n158), .I1(n157), .S(n534), .ZN(n162) );
  MUX2ND0 U525 ( .I0(n160), .I1(n159), .S(n533), .ZN(n161) );
  MUX2ND0 U526 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n551), .ZN(
        n166) );
  MUX2ND0 U527 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n552), .ZN(
        n165) );
  MUX3ND0 U528 ( .I0(n169), .I1(n168), .I2(n164), .S0(n536), .S1(n532), .ZN(
        n176) );
  MUX2ND0 U529 ( .I0(n171), .I1(n170), .S(n533), .ZN(n175) );
  MUX2ND0 U530 ( .I0(n173), .I1(n172), .S(n535), .ZN(n174) );
  MUX2ND0 U531 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n552), .ZN(
        n179) );
  MUX2ND0 U532 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n552), .ZN(
        n178) );
  MUX3ND0 U533 ( .I0(n182), .I1(n181), .I2(n177), .S0(n536), .S1(n530), .ZN(
        n189) );
  MUX2ND0 U534 ( .I0(n184), .I1(n183), .S(n606), .ZN(n188) );
  MUX2ND0 U535 ( .I0(n186), .I1(n185), .S(n533), .ZN(n187) );
  MUX2ND0 U536 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n552), .ZN(
        n192) );
  MUX2ND0 U537 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n552), .ZN(
        n191) );
  MUX3ND0 U538 ( .I0(n195), .I1(n194), .I2(n190), .S0(n606), .S1(n530), .ZN(
        n202) );
  MUX2ND0 U539 ( .I0(n197), .I1(n196), .S(n535), .ZN(n201) );
  MUX2ND0 U540 ( .I0(n199), .I1(n198), .S(n606), .ZN(n200) );
  MUX2ND0 U541 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n547), .ZN(
        n205) );
  MUX2ND0 U542 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n552), .ZN(
        n204) );
  MUX3ND0 U543 ( .I0(n208), .I1(n207), .I2(n203), .S0(n536), .S1(n530), .ZN(
        n215) );
  MUX2ND0 U544 ( .I0(n210), .I1(n209), .S(n534), .ZN(n214) );
  MUX2ND0 U545 ( .I0(n212), .I1(n211), .S(n606), .ZN(n213) );
  MUX2ND0 U546 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n552), .ZN(
        n218) );
  MUX2ND0 U547 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n555), .ZN(
        n217) );
  MUX3ND0 U548 ( .I0(n221), .I1(n220), .I2(n216), .S0(n536), .S1(n530), .ZN(
        n228) );
  MUX2ND0 U549 ( .I0(n223), .I1(n222), .S(n533), .ZN(n227) );
  MUX2ND0 U550 ( .I0(n225), .I1(n224), .S(n535), .ZN(n226) );
  MUX2ND0 U551 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n554), 
        .ZN(n231) );
  MUX2ND0 U552 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n552), 
        .ZN(n230) );
  MUX3ND0 U553 ( .I0(n234), .I1(n233), .I2(n229), .S0(n536), .S1(n530), .ZN(
        n241) );
  MUX2ND0 U554 ( .I0(n236), .I1(n235), .S(n533), .ZN(n240) );
  MUX2ND0 U555 ( .I0(n238), .I1(n237), .S(n535), .ZN(n239) );
  MUX2ND0 U556 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n552), 
        .ZN(n244) );
  MUX2ND0 U557 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n552), 
        .ZN(n243) );
  MUX3ND0 U558 ( .I0(n247), .I1(n246), .I2(n242), .S0(n606), .S1(n530), .ZN(
        n254) );
  MUX2ND0 U559 ( .I0(n249), .I1(n248), .S(n533), .ZN(n253) );
  MUX2ND0 U560 ( .I0(n251), .I1(n250), .S(N46), .ZN(n252) );
  MUX2ND0 U561 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n552), 
        .ZN(n257) );
  MUX2ND0 U562 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n552), 
        .ZN(n256) );
  MUX3ND0 U563 ( .I0(n260), .I1(n259), .I2(n255), .S0(n533), .S1(n530), .ZN(
        n267) );
  MUX2ND0 U564 ( .I0(n262), .I1(n261), .S(n533), .ZN(n266) );
  MUX2ND0 U565 ( .I0(n264), .I1(n263), .S(N46), .ZN(n265) );
  MUX2ND0 U566 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n552), 
        .ZN(n270) );
  MUX2ND0 U567 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n552), 
        .ZN(n269) );
  MUX3ND0 U568 ( .I0(n273), .I1(n272), .I2(n268), .S0(n533), .S1(n530), .ZN(
        n280) );
  MUX2ND0 U569 ( .I0(n275), .I1(n274), .S(n535), .ZN(n279) );
  MUX2ND0 U570 ( .I0(n277), .I1(n276), .S(n533), .ZN(n278) );
  MUX2ND0 U571 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n552), 
        .ZN(n283) );
  MUX2ND0 U572 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n552), 
        .ZN(n282) );
  MUX3ND0 U573 ( .I0(n286), .I1(n285), .I2(n281), .S0(n606), .S1(n530), .ZN(
        n293) );
  MUX2ND0 U574 ( .I0(n288), .I1(n287), .S(n535), .ZN(n292) );
  MUX2ND0 U575 ( .I0(n290), .I1(n289), .S(n533), .ZN(n291) );
  MUX2ND0 U576 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n552), 
        .ZN(n296) );
  MUX2ND0 U577 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n552), 
        .ZN(n295) );
  MUX3ND0 U578 ( .I0(n299), .I1(n298), .I2(n294), .S0(n535), .S1(n530), .ZN(
        n306) );
  MUX2ND0 U579 ( .I0(n301), .I1(n300), .S(n533), .ZN(n305) );
  MUX2ND0 U580 ( .I0(n303), .I1(n302), .S(n606), .ZN(n304) );
  MUX2ND0 U581 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n552), 
        .ZN(n309) );
  MUX2ND0 U582 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n552), 
        .ZN(n308) );
  MUX3ND0 U583 ( .I0(n312), .I1(n311), .I2(n307), .S0(n536), .S1(n530), .ZN(
        n319) );
  MUX2ND0 U584 ( .I0(n314), .I1(n313), .S(n533), .ZN(n318) );
  MUX2ND0 U585 ( .I0(n316), .I1(n315), .S(N46), .ZN(n317) );
  MUX2ND0 U586 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n551), 
        .ZN(n322) );
  MUX2ND0 U587 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n552), 
        .ZN(n321) );
  MUX3ND0 U588 ( .I0(n325), .I1(n324), .I2(n320), .S0(n533), .S1(n530), .ZN(
        n332) );
  MUX2ND0 U589 ( .I0(n327), .I1(n326), .S(n536), .ZN(n331) );
  MUX2ND0 U590 ( .I0(n329), .I1(n328), .S(N46), .ZN(n330) );
  MUX2ND0 U591 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n552), 
        .ZN(n335) );
  MUX2ND0 U592 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n551), 
        .ZN(n334) );
  MUX3ND0 U593 ( .I0(n338), .I1(n337), .I2(n333), .S0(n533), .S1(n530), .ZN(
        n345) );
  MUX2ND0 U594 ( .I0(n340), .I1(n339), .S(N46), .ZN(n344) );
  MUX2ND0 U595 ( .I0(n342), .I1(n341), .S(N46), .ZN(n343) );
  MUX2ND0 U596 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n551), 
        .ZN(n348) );
  MUX2ND0 U597 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n551), 
        .ZN(n347) );
  MUX3ND0 U598 ( .I0(n351), .I1(n350), .I2(n346), .S0(N46), .S1(n532), .ZN(
        n358) );
  MUX2ND0 U599 ( .I0(n353), .I1(n352), .S(N46), .ZN(n357) );
  MUX2ND0 U600 ( .I0(n355), .I1(n354), .S(n533), .ZN(n356) );
  MUX2ND0 U601 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n551), 
        .ZN(n361) );
  MUX2ND0 U602 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n551), 
        .ZN(n360) );
  MUX3ND0 U603 ( .I0(n364), .I1(n363), .I2(n359), .S0(n533), .S1(n532), .ZN(
        n371) );
  MUX2ND0 U604 ( .I0(n366), .I1(n365), .S(N46), .ZN(n370) );
  MUX2ND0 U605 ( .I0(n368), .I1(n367), .S(n533), .ZN(n369) );
  MUX2ND0 U606 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n551), 
        .ZN(n374) );
  MUX2ND0 U607 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n551), 
        .ZN(n373) );
  MUX3ND0 U608 ( .I0(n377), .I1(n376), .I2(n372), .S0(N46), .S1(n532), .ZN(
        n384) );
  MUX2ND0 U609 ( .I0(n379), .I1(n378), .S(N46), .ZN(n383) );
  MUX2ND0 U610 ( .I0(n381), .I1(n380), .S(n606), .ZN(n382) );
  MUX2ND0 U611 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n551), 
        .ZN(n387) );
  MUX2ND0 U612 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n551), 
        .ZN(n386) );
  MUX3ND0 U613 ( .I0(n390), .I1(n389), .I2(n385), .S0(n536), .S1(n532), .ZN(
        n397) );
  MUX2ND0 U614 ( .I0(n392), .I1(n391), .S(n533), .ZN(n396) );
  MUX2ND0 U615 ( .I0(n394), .I1(n393), .S(n534), .ZN(n395) );
  MUX2ND0 U616 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n551), 
        .ZN(n400) );
  MUX2ND0 U617 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n551), 
        .ZN(n399) );
  MUX3ND0 U618 ( .I0(n403), .I1(n402), .I2(n398), .S0(n533), .S1(n532), .ZN(
        n410) );
  MUX2ND0 U619 ( .I0(n405), .I1(n404), .S(n535), .ZN(n409) );
  MUX2ND0 U620 ( .I0(n407), .I1(n406), .S(n534), .ZN(n408) );
  MUX2ND0 U621 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n551), 
        .ZN(n413) );
  MUX2ND0 U622 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n551), 
        .ZN(n412) );
  MUX3ND0 U623 ( .I0(n416), .I1(n415), .I2(n411), .S0(n533), .S1(n532), .ZN(
        n423) );
  MUX2ND0 U624 ( .I0(n418), .I1(n417), .S(n536), .ZN(n422) );
  MUX2ND0 U625 ( .I0(n420), .I1(n419), .S(n534), .ZN(n421) );
  MUX2ND0 U626 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n551), 
        .ZN(n426) );
  MUX2ND0 U627 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n551), 
        .ZN(n425) );
  MUX3ND0 U628 ( .I0(n429), .I1(n428), .I2(n424), .S0(n606), .S1(n530), .ZN(
        n436) );
  MUX2ND0 U629 ( .I0(n431), .I1(n430), .S(n535), .ZN(n435) );
  MUX2ND0 U630 ( .I0(n433), .I1(n432), .S(n534), .ZN(n434) );
  MUX2ND0 U631 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n551), 
        .ZN(n439) );
  MUX2ND0 U632 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n550), 
        .ZN(n438) );
  MUX3ND0 U633 ( .I0(n442), .I1(n441), .I2(n437), .S0(n536), .S1(n531), .ZN(
        n449) );
  MUX2ND0 U634 ( .I0(n444), .I1(n443), .S(n535), .ZN(n448) );
  MUX2ND0 U635 ( .I0(n446), .I1(n445), .S(n535), .ZN(n447) );
  MUX2ND0 U636 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n550), 
        .ZN(n452) );
  MUX2ND0 U637 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n550), 
        .ZN(n451) );
  MUX3ND0 U638 ( .I0(n455), .I1(n454), .I2(n450), .S0(n606), .S1(n532), .ZN(
        n462) );
  MUX2ND0 U639 ( .I0(n457), .I1(n456), .S(n534), .ZN(n461) );
  MUX2ND0 U640 ( .I0(n459), .I1(n458), .S(n534), .ZN(n460) );
  MUX2ND0 U641 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n550), 
        .ZN(n465) );
  MUX2ND0 U642 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n550), 
        .ZN(n464) );
  MUX3ND0 U643 ( .I0(n468), .I1(n467), .I2(n463), .S0(n536), .S1(N47), .ZN(
        n475) );
  MUX2ND0 U644 ( .I0(n470), .I1(n469), .S(n535), .ZN(n474) );
  MUX2ND0 U645 ( .I0(n472), .I1(n471), .S(n606), .ZN(n473) );
  MUX2ND0 U646 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n550), 
        .ZN(n478) );
  MUX2ND0 U647 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n550), 
        .ZN(n477) );
  MUX3ND0 U648 ( .I0(n481), .I1(n480), .I2(n476), .S0(n536), .S1(N47), .ZN(
        n488) );
  MUX2ND0 U649 ( .I0(n483), .I1(n482), .S(n534), .ZN(n487) );
  MUX2ND0 U650 ( .I0(n485), .I1(n484), .S(n606), .ZN(n486) );
  MUX2ND0 U651 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n550), 
        .ZN(n491) );
  MUX2ND0 U652 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n550), 
        .ZN(n490) );
  MUX3ND0 U653 ( .I0(n494), .I1(n493), .I2(n489), .S0(n536), .S1(N47), .ZN(
        n501) );
  MUX2ND0 U654 ( .I0(n496), .I1(n495), .S(n606), .ZN(n500) );
  MUX2ND0 U655 ( .I0(n498), .I1(n497), .S(n606), .ZN(n499) );
  MUX2ND0 U656 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n550), 
        .ZN(n504) );
  MUX2ND0 U657 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n550), 
        .ZN(n503) );
  MUX3ND0 U658 ( .I0(n507), .I1(n506), .I2(n502), .S0(n536), .S1(N47), .ZN(
        n514) );
  MUX2ND0 U659 ( .I0(n509), .I1(n508), .S(n535), .ZN(n513) );
  MUX2ND0 U660 ( .I0(n511), .I1(n510), .S(n606), .ZN(n512) );
  MUX2ND0 U661 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n550), 
        .ZN(n517) );
  MUX2ND0 U662 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n552), 
        .ZN(n516) );
  MUX3ND0 U663 ( .I0(n520), .I1(n519), .I2(n515), .S0(n536), .S1(n530), .ZN(
        n527) );
  MUX2ND0 U664 ( .I0(n522), .I1(n521), .S(n606), .ZN(n526) );
  MUX2ND0 U665 ( .I0(n524), .I1(n523), .S(n606), .ZN(n525) );
endmodule


module MemBIST_Top ( Dready, ParityErr, Testing, TestOK, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, DoSelfTest, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, DoSelfTest, Read, Write, Reset;
  output Dready, ParityErr, Testing, TestOK;
  wire   N9, n195, Dreadyw, ClkWw, Readw, ReadCmdBISTw, Writew, WriteCmdBISTw,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n161, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194;
  wire   [31:0] DataOw;
  wire   [31:0] DataIw;
  wire   [31:0] DataOBISTw;
  wire   [4:0] AddrRw;
  wire   [4:0] AddrBISTw;
  wire   [4:0] AddrWw;
  wire   [31:0] DataIBISTw;

  Mem_AWid5_DWid32 Mem_U1 ( .Dready(Dreadyw), .ParityErr(n195), .DataO(DataOw), 
        .DataI({n188, n187, n186, n185, n184, n183, n182, n181, n180, n179, 
        n178, n177, n176, n175, n174, n173, DataIw[15:13], n172, n171, n170, 
        n169, n168, DataIw[7:5], n167, n166, n165, n164, n163}), .AddrR(AddrRw), .AddrW(AddrWw), .ClkR(ClkR), .ClkW(ClkWw), .ChipEna(n189), .Read(Readw), 
        .Write(Writew), .Reset(n157) );
  BIST_AWid5_DWid32 BIST_U1 ( .DataO(DataOBISTw), .Addr(AddrBISTw), .ReadCmd(
        ReadCmdBISTw), .WriteCmd(WriteCmdBISTw), .Testing(N9), .TestOK(TestOK), 
        .DataI(DataIBISTw), .DoSelfTest(DoSelfTest), .ParityErr(n132), .Clk(
        ClkR), .Reset(n155) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOw[29]), .OE(n193), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOw[19]), .OE(n194), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOw[28]), .OE(n194), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOw[18]), .OE(n194), .Z(DataO[18]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOw[27]), .OE(n191), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOw[17]), .OE(n191), .Z(DataO[17]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOw[26]), .OE(n194), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOw[16]), .OE(n191), .Z(DataO[16]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOw[25]), .OE(n193), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOw[15]), .OE(n191), .Z(DataO[15]) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOw[31]), .OE(n193), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOw[24]), .OE(n194), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOw[14]), .OE(n191), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOw[30]), .OE(n193), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOw[23]), .OE(n192), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOw[13]), .OE(n191), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOw[9]), .OE(n191), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOw[22]), .OE(n194), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOw[12]), .OE(n191), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOw[8]), .OE(n191), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOw[21]), .OE(n191), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOw[11]), .OE(n191), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOw[7]), .OE(n194), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOw[20]), .OE(n191), .Z(DataO[20]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOw[10]), .OE(n191), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOw[6]), .OE(n194), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOw[5]), .OE(n194), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOw[4]), .OE(n191), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOw[3]), .OE(n193), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[0]  ( .I(DataOw[0]), .OE(n191), .Z(DataO[0]) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOw[1]), .OE(n191), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOw[2]), .OE(n194), .Z(DataO[2]) );
  BUFTD0 \DataIBISTw_tri[12]  ( .I(DataOw[12]), .OE(n190), .Z(DataIBISTw[12])
         );
  BUFTD0 \DataIBISTw_tri[16]  ( .I(DataOw[16]), .OE(n190), .Z(DataIBISTw[16])
         );
  BUFTD0 \DataIBISTw_tri[15]  ( .I(DataOw[15]), .OE(n190), .Z(DataIBISTw[15])
         );
  BUFTD0 \DataIBISTw_tri[24]  ( .I(DataOw[24]), .OE(n190), .Z(DataIBISTw[24])
         );
  BUFTD0 \DataIBISTw_tri[28]  ( .I(DataOw[28]), .OE(n190), .Z(DataIBISTw[28])
         );
  BUFTD0 \DataIBISTw_tri[14]  ( .I(DataOw[14]), .OE(n190), .Z(DataIBISTw[14])
         );
  BUFTD0 \DataIBISTw_tri[0]  ( .I(DataOw[0]), .OE(n190), .Z(DataIBISTw[0]) );
  BUFTD0 \DataIBISTw_tri[13]  ( .I(DataOw[13]), .OE(n190), .Z(DataIBISTw[13])
         );
  BUFTD0 \DataIBISTw_tri[29]  ( .I(DataOw[29]), .OE(n190), .Z(DataIBISTw[29])
         );
  BUFTD0 \DataIBISTw_tri[27]  ( .I(DataOw[27]), .OE(n190), .Z(DataIBISTw[27])
         );
  BUFTD0 \DataIBISTw_tri[23]  ( .I(DataOw[23]), .OE(n190), .Z(DataIBISTw[23])
         );
  BUFTD0 \DataIBISTw_tri[11]  ( .I(DataOw[11]), .OE(n190), .Z(DataIBISTw[11])
         );
  BUFTD0 \DataIBISTw_tri[22]  ( .I(DataOw[22]), .OE(n190), .Z(DataIBISTw[22])
         );
  BUFTD0 \DataIBISTw_tri[26]  ( .I(DataOw[26]), .OE(n190), .Z(DataIBISTw[26])
         );
  BUFTD0 \DataIBISTw_tri[21]  ( .I(DataOw[21]), .OE(n190), .Z(DataIBISTw[21])
         );
  BUFTD0 \DataIBISTw_tri[10]  ( .I(DataOw[10]), .OE(n190), .Z(DataIBISTw[10])
         );
  BUFTD0 \DataIBISTw_tri[20]  ( .I(DataOw[20]), .OE(n190), .Z(DataIBISTw[20])
         );
  BUFTD0 \DataIBISTw_tri[19]  ( .I(DataOw[19]), .OE(n190), .Z(DataIBISTw[19])
         );
  BUFTD0 \DataIBISTw_tri[1]  ( .I(DataOw[1]), .OE(n190), .Z(DataIBISTw[1]) );
  BUFTD0 \DataIBISTw_tri[25]  ( .I(DataOw[25]), .OE(n190), .Z(DataIBISTw[25])
         );
  BUFTD0 \DataIBISTw_tri[17]  ( .I(DataOw[17]), .OE(n190), .Z(DataIBISTw[17])
         );
  BUFTD0 \DataIBISTw_tri[18]  ( .I(DataOw[18]), .OE(n190), .Z(DataIBISTw[18])
         );
  BUFTD0 \DataIBISTw_tri[30]  ( .I(DataOw[30]), .OE(n190), .Z(DataIBISTw[30])
         );
  BUFTD0 \DataIBISTw_tri[4]  ( .I(DataOw[4]), .OE(n190), .Z(DataIBISTw[4]) );
  BUFTD0 \DataIBISTw_tri[5]  ( .I(DataOw[5]), .OE(n190), .Z(DataIBISTw[5]) );
  BUFTD0 \DataIBISTw_tri[8]  ( .I(DataOw[8]), .OE(n190), .Z(DataIBISTw[8]) );
  BUFTD0 \DataIBISTw_tri[31]  ( .I(DataOw[31]), .OE(n190), .Z(DataIBISTw[31])
         );
  BUFTD0 \DataIBISTw_tri[6]  ( .I(DataOw[6]), .OE(n190), .Z(DataIBISTw[6]) );
  BUFTD0 \DataIBISTw_tri[9]  ( .I(DataOw[9]), .OE(n190), .Z(DataIBISTw[9]) );
  BUFTD0 \DataIBISTw_tri[7]  ( .I(DataOw[7]), .OE(n190), .Z(DataIBISTw[7]) );
  BUFTD0 \DataIBISTw_tri[2]  ( .I(DataOw[2]), .OE(n190), .Z(DataIBISTw[2]) );
  BUFTD0 \DataIBISTw_tri[3]  ( .I(DataOw[3]), .OE(n190), .Z(DataIBISTw[3]) );
  CKNXD12 U49 ( .I(Reset), .ZN(n156) );
  INVD1 U50 ( .I(n131), .ZN(n132) );
  BUFFD1 U51 ( .I(n194), .Z(n192) );
  CKNXD16 U52 ( .I(n131), .ZN(ParityErr) );
  CKND0 U53 ( .CLK(n195), .CN(n131) );
  BUFFD0 U54 ( .I(Reset), .Z(n133) );
  BUFFD0 U55 ( .I(n133), .Z(n134) );
  BUFFD0 U56 ( .I(n134), .Z(n135) );
  BUFFD0 U57 ( .I(n135), .Z(n136) );
  BUFFD0 U58 ( .I(n136), .Z(n137) );
  BUFFD0 U59 ( .I(n137), .Z(n138) );
  BUFFD0 U60 ( .I(n138), .Z(n139) );
  BUFFD0 U61 ( .I(n139), .Z(n140) );
  BUFFD0 U62 ( .I(n140), .Z(n141) );
  BUFFD0 U63 ( .I(n141), .Z(n142) );
  BUFFD0 U64 ( .I(n142), .Z(n143) );
  BUFFD0 U65 ( .I(n143), .Z(n144) );
  BUFFD0 U66 ( .I(n144), .Z(n145) );
  BUFFD0 U67 ( .I(n145), .Z(n146) );
  BUFFD0 U68 ( .I(n146), .Z(n147) );
  BUFFD0 U69 ( .I(n147), .Z(n148) );
  BUFFD0 U70 ( .I(n148), .Z(n149) );
  BUFFD0 U71 ( .I(n149), .Z(n150) );
  BUFFD0 U72 ( .I(n150), .Z(n151) );
  BUFFD0 U73 ( .I(n151), .Z(n152) );
  BUFFD0 U74 ( .I(n152), .Z(n153) );
  BUFFD0 U75 ( .I(n153), .Z(n154) );
  BUFFD0 U76 ( .I(n154), .Z(n155) );
  INVD0 U77 ( .I(n156), .ZN(n157) );
  CKNXD0 U78 ( .I(n158), .ZN(n159) );
  CKBD1 U79 ( .CLK(n159), .C(n189) );
  INVD8 U80 ( .I(ChipEna), .ZN(n158) );
  CKNXD16 U81 ( .I(n192), .ZN(Testing) );
  CKND2D0 U82 ( .A1(Dreadyw), .A2(n194), .ZN(n161) );
  INVD1 U83 ( .I(N9), .ZN(n194) );
  CKND16 U84 ( .CLK(n161), .CN(Dready) );
  INVD3 U85 ( .I(n194), .ZN(n190) );
  BUFFD1 U86 ( .I(n193), .Z(n191) );
  BUFFD1 U87 ( .I(n194), .Z(n193) );
  AO22D0 U88 ( .A1(n190), .A2(AddrBISTw[0]), .B1(AddrR[0]), .B2(n192), .Z(
        AddrRw[0]) );
  AO22D0 U89 ( .A1(n190), .A2(AddrBISTw[1]), .B1(AddrR[1]), .B2(n193), .Z(
        AddrRw[1]) );
  AO22D0 U90 ( .A1(n190), .A2(AddrBISTw[4]), .B1(AddrR[4]), .B2(n193), .Z(
        AddrRw[4]) );
  AO22D0 U91 ( .A1(n190), .A2(AddrBISTw[2]), .B1(AddrR[2]), .B2(n193), .Z(
        AddrRw[2]) );
  AO22D0 U92 ( .A1(n190), .A2(AddrBISTw[3]), .B1(AddrR[3]), .B2(n193), .Z(
        AddrRw[3]) );
  AO22D0 U93 ( .A1(n190), .A2(AddrBISTw[2]), .B1(AddrW[2]), .B2(n193), .Z(
        AddrWw[2]) );
  AO22D0 U94 ( .A1(n190), .A2(AddrBISTw[0]), .B1(AddrW[0]), .B2(n193), .Z(
        AddrWw[0]) );
  AO22D0 U95 ( .A1(n190), .A2(AddrBISTw[1]), .B1(AddrW[1]), .B2(n193), .Z(
        AddrWw[1]) );
  AO22D0 U96 ( .A1(n190), .A2(AddrBISTw[3]), .B1(AddrW[3]), .B2(n193), .Z(
        AddrWw[3]) );
  AO22D0 U97 ( .A1(n190), .A2(AddrBISTw[4]), .B1(AddrW[4]), .B2(n193), .Z(
        AddrWw[4]) );
  BUFFD1 U98 ( .I(DataIw[24]), .Z(n181) );
  AO22D0 U99 ( .A1(DataOBISTw[24]), .A2(n190), .B1(DataI[24]), .B2(n193), .Z(
        DataIw[24]) );
  BUFFD1 U100 ( .I(DataIw[25]), .Z(n182) );
  AO22D0 U101 ( .A1(DataOBISTw[25]), .A2(n190), .B1(DataI[25]), .B2(n192), .Z(
        DataIw[25]) );
  BUFFD1 U102 ( .I(DataIw[26]), .Z(n183) );
  AO22D0 U103 ( .A1(DataOBISTw[26]), .A2(n190), .B1(DataI[26]), .B2(n192), .Z(
        DataIw[26]) );
  BUFFD1 U104 ( .I(DataIw[27]), .Z(n184) );
  AO22D0 U105 ( .A1(DataOBISTw[27]), .A2(n190), .B1(DataI[27]), .B2(n192), .Z(
        DataIw[27]) );
  BUFFD1 U106 ( .I(DataIw[28]), .Z(n185) );
  AO22D0 U107 ( .A1(DataOBISTw[28]), .A2(n190), .B1(DataI[28]), .B2(n192), .Z(
        DataIw[28]) );
  BUFFD1 U108 ( .I(DataIw[29]), .Z(n186) );
  AO22D0 U109 ( .A1(DataOBISTw[29]), .A2(n190), .B1(DataI[29]), .B2(n192), .Z(
        DataIw[29]) );
  BUFFD1 U110 ( .I(DataIw[30]), .Z(n187) );
  AO22D0 U111 ( .A1(DataOBISTw[30]), .A2(n190), .B1(DataI[30]), .B2(n192), .Z(
        DataIw[30]) );
  BUFFD1 U112 ( .I(DataIw[31]), .Z(n188) );
  AO22D0 U113 ( .A1(DataOBISTw[31]), .A2(n190), .B1(DataI[31]), .B2(n192), .Z(
        DataIw[31]) );
  AO22D0 U114 ( .A1(WriteCmdBISTw), .A2(n190), .B1(Write), .B2(n192), .Z(
        Writew) );
  AO22D0 U115 ( .A1(ReadCmdBISTw), .A2(n190), .B1(Read), .B2(n193), .Z(Readw)
         );
  BUFFD1 U116 ( .I(DataIw[0]), .Z(n163) );
  AO22D0 U117 ( .A1(DataOBISTw[0]), .A2(n190), .B1(DataI[0]), .B2(n193), .Z(
        DataIw[0]) );
  BUFFD1 U118 ( .I(DataIw[1]), .Z(n164) );
  AO22D0 U119 ( .A1(DataOBISTw[1]), .A2(n190), .B1(DataI[1]), .B2(n192), .Z(
        DataIw[1]) );
  BUFFD1 U120 ( .I(DataIw[2]), .Z(n165) );
  AO22D0 U121 ( .A1(DataOBISTw[2]), .A2(n190), .B1(DataI[2]), .B2(n192), .Z(
        DataIw[2]) );
  BUFFD1 U122 ( .I(DataIw[3]), .Z(n166) );
  AO22D0 U123 ( .A1(DataOBISTw[3]), .A2(n190), .B1(DataI[3]), .B2(n193), .Z(
        DataIw[3]) );
  BUFFD1 U124 ( .I(DataIw[4]), .Z(n167) );
  AO22D0 U125 ( .A1(DataOBISTw[4]), .A2(n190), .B1(DataI[4]), .B2(n193), .Z(
        DataIw[4]) );
  AO22D0 U126 ( .A1(DataOBISTw[5]), .A2(n190), .B1(DataI[5]), .B2(n193), .Z(
        DataIw[5]) );
  AO22D0 U127 ( .A1(DataOBISTw[6]), .A2(n190), .B1(DataI[6]), .B2(n193), .Z(
        DataIw[6]) );
  AO22D0 U128 ( .A1(DataOBISTw[7]), .A2(n190), .B1(DataI[7]), .B2(n193), .Z(
        DataIw[7]) );
  BUFFD1 U129 ( .I(DataIw[8]), .Z(n168) );
  AO22D0 U130 ( .A1(DataOBISTw[8]), .A2(n190), .B1(DataI[8]), .B2(n193), .Z(
        DataIw[8]) );
  BUFFD1 U131 ( .I(DataIw[9]), .Z(n169) );
  AO22D0 U132 ( .A1(DataOBISTw[9]), .A2(n190), .B1(DataI[9]), .B2(n193), .Z(
        DataIw[9]) );
  BUFFD1 U133 ( .I(DataIw[10]), .Z(n170) );
  AO22D0 U134 ( .A1(DataOBISTw[10]), .A2(n190), .B1(DataI[10]), .B2(n193), .Z(
        DataIw[10]) );
  BUFFD1 U135 ( .I(DataIw[11]), .Z(n171) );
  AO22D0 U136 ( .A1(DataOBISTw[11]), .A2(n190), .B1(DataI[11]), .B2(n193), .Z(
        DataIw[11]) );
  BUFFD1 U137 ( .I(DataIw[12]), .Z(n172) );
  AO22D0 U138 ( .A1(DataOBISTw[12]), .A2(n190), .B1(DataI[12]), .B2(n193), .Z(
        DataIw[12]) );
  AO22D0 U139 ( .A1(DataOBISTw[13]), .A2(n190), .B1(DataI[13]), .B2(n193), .Z(
        DataIw[13]) );
  AO22D0 U140 ( .A1(DataOBISTw[14]), .A2(n190), .B1(DataI[14]), .B2(n193), .Z(
        DataIw[14]) );
  AO22D0 U141 ( .A1(DataOBISTw[15]), .A2(n190), .B1(DataI[15]), .B2(n193), .Z(
        DataIw[15]) );
  BUFFD1 U142 ( .I(DataIw[16]), .Z(n173) );
  AO22D0 U143 ( .A1(DataOBISTw[16]), .A2(n190), .B1(DataI[16]), .B2(n192), .Z(
        DataIw[16]) );
  BUFFD1 U144 ( .I(DataIw[17]), .Z(n174) );
  AO22D0 U145 ( .A1(DataOBISTw[17]), .A2(n190), .B1(DataI[17]), .B2(n192), .Z(
        DataIw[17]) );
  BUFFD1 U146 ( .I(DataIw[18]), .Z(n175) );
  AO22D0 U147 ( .A1(DataOBISTw[18]), .A2(n190), .B1(DataI[18]), .B2(n192), .Z(
        DataIw[18]) );
  BUFFD1 U148 ( .I(DataIw[19]), .Z(n176) );
  AO22D0 U149 ( .A1(DataOBISTw[19]), .A2(n190), .B1(DataI[19]), .B2(n192), .Z(
        DataIw[19]) );
  BUFFD1 U150 ( .I(DataIw[20]), .Z(n177) );
  AO22D0 U151 ( .A1(DataOBISTw[20]), .A2(n190), .B1(DataI[20]), .B2(n192), .Z(
        DataIw[20]) );
  BUFFD1 U152 ( .I(DataIw[21]), .Z(n178) );
  AO22D0 U153 ( .A1(DataOBISTw[21]), .A2(n190), .B1(DataI[21]), .B2(n192), .Z(
        DataIw[21]) );
  BUFFD1 U154 ( .I(DataIw[22]), .Z(n179) );
  AO22D0 U155 ( .A1(DataOBISTw[22]), .A2(n190), .B1(DataI[22]), .B2(n192), .Z(
        DataIw[22]) );
  BUFFD1 U156 ( .I(DataIw[23]), .Z(n180) );
  AO22D0 U157 ( .A1(DataOBISTw[23]), .A2(n190), .B1(DataI[23]), .B2(n192), .Z(
        DataIw[23]) );
  AO22D0 U158 ( .A1(ClkW), .A2(n192), .B1(ClkR), .B2(n190), .Z(ClkWw) );
endmodule

