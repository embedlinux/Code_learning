//----------------------------------------------------------------------------------
// Design Unit : Byte input FF received CRC
// Version : v1.0 2007/05/26
//----------------------------------------------------------------------------------
module ff_rcv_fcs_8b(clk,rst,en,d,fok);
input clk;
input rst;
input en;
input[7:0] d;
output fok;
//----------------------------------------------------------------------------------
//----------------------------------------------------------------------------------
reg[15:0] q;
wire[15:0] qf;
wire[15:0] qi;
wire fok;
//----------------------------------------------------------------------------------
//----------------------------------------------------------------------------------
always @(posedge clk or posedge rst)
begin
    if(rst == 1'b1)
        q <= 16'hffff;
    else if(en == 1'b1)
        q <= qi;
end
//----------------------------------------------------------------------------------
//----------------------------------------------------------------------------------
assign qf[0]  = q[8] ^ q[12] ^ q[13] ^ q[14];
assign qf[1]  = q[8] ^ q[9]  ^ q[12] ^ q[15];
assign qf[2]  = q[8] ^ q[9] ^ q[10] ^ q[12] ^ q[14];
assign qf[3]  = q[8] ^ q[9] ^ q[10] ^ q[11] ^ q[12] ^ q[14] ^ q[15];
assign qf[4]  = q[8] ^ q[9] ^ q[10] ^ q[11] ^ q[14] ^ q[15];
assign qf[5]  = q[9] ^ q[10] ^ q[11] ^ q[12];
assign qf[6]  = q[8] ^ q[11] ^ q[15];
assign qf[7]  = q[8] ^ q[9] ^ q[13] ^ q[14];
assign qf[8]  = q[0] ^ q[8] ^ q[9] ^ q[10] ^ q[12] ^ q[13] ^ q[15];
assign qf[9]  = q[1] ^ q[9] ^ q[10] ^ q[11] ^ q[13] ^ q[14];
assign qf[10] = q[2] ^ q[8] ^ q[10] ^ q[11] ^ q[13] ^ q[15];
assign qf[11] = q[3] ^ q[8] ^ q[9] ^ q[11] ^ q[13];
assign qf[12] = q[4] ^ q[8] ^ q[9] ^ q[10] ^ q[13];
assign qf[13] = q[5] ^ q[9] ^ q[10] ^ q[11] ^ q[14];
assign qf[14] = q[6] ^ q[10] ^ q[11] ^ q[12] ^ q[15];
assign qf[15] = q[7] ^ q[11] ^ q[12] ^ q[13];
//----------------------------------------------------------------------------------
//----------------------------------------------------------------------------------
assign qi[0]  = (d[0] ^ d[4] ^ d[5] ^ d[6]) ^ qf[0]; 
assign qi[1]  = (d[0] ^ d[1] ^ d[4] ^ d[7]) ^ qf[1]; 
assign qi[2]  = (d[0] ^ d[1] ^ d[2] ^ d[4] ^ d[6]) ^ qf[2];
assign qi[3]  = (d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[4] ^ d[6] ^ d[7]) ^ qf[3];
assign qi[4]  = (d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[6] ^ d[7]) ^ qf[4];
assign qi[5]  = (d[1] ^ d[2] ^ d[3] ^ d[4] ^ d[7]) ^ qf[5];
assign qi[6]  = (d[0] ^ d[3] ^ d[7]) ^ qf[6];
assign qi[7]  = (d[0] ^ d[1] ^ d[5] ^ d[6]) ^ qf[7];
assign qi[8]  = (d[0] ^ d[1] ^ d[2] ^ d[4] ^ d[5] ^ d[7]) ^ qf[8];
assign qi[9]  = (d[1] ^ d[2] ^ d[3] ^ d[5] ^ d[6]) ^ qf[9];
assign qi[10] = (d[0] ^ d[2] ^ d[3] ^ d[5] ^ d[7]) ^ qf[10];
assign qi[11] = (d[0] ^ d[1] ^ d[3] ^ d[5]) ^ qf[11];
assign qi[12] = (d[0] ^ d[1] ^ d[2] ^ d[5]) ^ qf[12];
assign qi[13] = (d[1] ^ d[2] ^ d[3] ^ d[6]) ^ qf[13];
assign qi[14] = (d[2] ^ d[3] ^ d[4] ^ d[7]) ^ qf[14];
assign qi[15] = (d[3] ^ d[4] ^ d[5]) ^ qf[15];
//-----------------------------------------------------------------------------------
assign fok = !q[0] & !q[1] & q[2] & !q[3] & q[4] & !q[5] & !q[6] & q[7] 
             & q[8] & q[9] & !q[10] & !q[11] & !q[12] & q[13] & q[14] & q[15];
//-----------------------------------------------------------------------------------
endmodule