//----------------------------------------------------------------------------------------------------------
// Design Unit : Byte input FF received CRC
// Version : v0.1 2007/05/20
//----------------------------------------------------------------------------------------------------------
module ff_rcv_fcs(clk,rst,en,d,fok);
input clk;
input rst;
input en;
input[7:0] d;
output fok;
//-----------------------------------------------------------------------------------------------------------
//-----------------------------------------------------------------------------------------------------------
reg[15:0] q;
wire[15:0] qi;
wire fok;
//-----------------------------------------------------------------------------------------------------------
//-----------------------------------------------------------------------------------------------------------
always @(posedge clk or posedge rst)
begin
    if(rst == 1'b1)
        q <= 16'hffff;
    else if(en == 1'b1)
        q <= qi;
end
//------------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------------
assign qi[0]  = (d[0] ^ d[4] ^ d[5] ^ d[6]) ^ (q[8] ^ q[12] ^ q[13] ^ q[14]); 
assign qi[1]  = (d[0] ^ d[1] ^ d[4] ^ d[7]) ^ (q[8] ^ q[9]  ^ q[12] ^ q[15]); 
assign qi[2]  = (d[0] ^ d[1] ^ d[2] ^ d[4] ^ d[6]) ^ (q[8] ^ q[9] ^ q[10] ^ q[12] ^ q[14]);
assign qi[3]  = (d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[4] ^ d[6] ^ d[7]) ^ (q[8] ^ q[9] ^ q[10] ^ q[11] ^ q[12] ^ q[14] ^ q[15]);
assign qi[4]  = (d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[6] ^ d[7]) ^ (q[8] ^ q[9] ^ q[10] ^ q[11] ^ q[14] ^ q[15]);
assign qi[5]  = (d[1] ^ d[2] ^ d[3] ^ d[4] ^ d[7]) ^ (q[9] ^ q[10] ^ q[11] ^ q[12]);
assign qi[6]  = (d[0] ^ d[3] ^ d[7]) ^ (q[8] ^ q[11] ^ q[15]);
assign qi[7]  = (d[0] ^ d[1] ^ d[5] ^ d[6]) ^ (q[8] ^ q[9] ^ q[13] ^ q[14]);
assign qi[8]  = (d[0] ^ d[1] ^ d[2] ^ d[4] ^ d[5] ^ d[7]) ^ (q[0] ^ q[8] ^ q[9] ^ q[10] ^ q[12] ^ q[13] ^ q[15]);
assign qi[9]  = (d[1] ^ d[2] ^ d[3] ^ d[5] ^ d[6]) ^ (q[1] ^ q[9] ^ q[10] ^ q[11] ^ q[13] ^ q[14]);
assign qi[10] = (d[0] ^ d[2] ^ d[3] ^ d[5] ^ d[7]) ^ (q[2] ^ q[8] ^ q[10] ^ q[11] ^ q[13] ^ q[15]);
assign qi[11] = (d[0] ^ d[1] ^ d[3] ^ d[5]) ^ (q[3] ^ q[8] ^ q[9] ^ q[11] ^ q[13]);
assign qi[12] = (d[0] ^ d[1] ^ d[2] ^ d[5]) ^ (q[4] ^ q[8] ^ q[9] ^ q[10] ^ q[13]);
assign qi[13] = (d[1] ^ d[2] ^ d[3] ^ d[6]) ^ (q[5] ^ q[9] ^ q[10] ^ q[11] ^ q[14]);
assign qi[14] = (d[2] ^ d[3] ^ d[4] ^ d[7]) ^ (q[6] ^ q[10] ^ q[11] ^ q[12] ^ q[15]);
assign qi[15] = (d[3] ^ d[4] ^ d[5]) ^ (q[7] ^ q[11] ^ q[12] ^ q[13]);
//-----------------------------------------------------------------------------------------------------------
assign fok = !q[0] & !q[1] & q[2] & !q[3] & q[4] & !q[5] & !q[6] & q[7] 
             & q[8] & q[9] & !q[10] & !q[11] & !q[12] & q[13] & q[14] & q[15];
//------------------------------------------------------------------------------------------------------------
endmodule