library verilog;
use verilog.vl_types.all;
entity adc128s022_tb is
end adc128s022_tb;
