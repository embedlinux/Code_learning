
`ifndef RKV_I2C_VIRTUAL_SEQUENCES_SVH
`define RKV_I2C_VIRTUAL_SEQUENCES_SVH

`include "rkv_i2c_base_virtual_sequence.sv" 
`include "rkv_i2c_quick_reg_access_virt_seq.sv" 
`include "rkv_i2c_directed_tx_virt_seq.sv" 
`include "rkv_i2c_directed_rx_virt_seq.sv" 

`endif // RKV_I2C_VIRTUAL_SEQUENCES_SVH

