library verilog;
use verilog.vl_types.all;
entity decoder3_8_tb is
end decoder3_8_tb;
