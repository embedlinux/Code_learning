`ifndef __MY_SEQUENCER__SV__
`define __MY_SEQUENCER__SV__

typedef uvm_sequencer #(my_transaction) my_sequencer;

`endif // __MY_SEQUENCER__SV__