
module FullDup ( OutParDataA, OutParDataB, InParDataA, InParDataB, InParValidA, 
        InParValidB, ClockA, ClockB, Reset );
  output [31:0] OutParDataA;
  output [31:0] OutParDataB;
  input [31:0] InParDataA;
  input [31:0] InParDataB;
  input InParValidA, InParValidB, ClockA, ClockB, Reset;
  wire   \*Logic1* , SerLine1, SerLine2, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061;

  SerDes_DWid32_RxLogDepth4_TxLogDepth3 SerDes_U1 ( .ParOutRxClk(OutParDataB), 
        .SerLineXfer(SerLine1), .ParDataIn({n825, n845, n865, n885, n905, n925, 
        n945, n967, n771, n769, n989, n1011, n1033, n1055, n767, n781, n779, 
        n775, n777, n785, n783, n773, n793, n791, n789, n795, n799, n797, n787, 
        n805, n803, n801}), .InParClk(n1061), .InParValid(n1059), .OutParClk(
        n1060), .RxRequest(\*Logic1* ), .TxRequest(n1059), .Reset(n21) );
  SerDes_DWid32_RxLogDepth3_TxLogDepth4 SerDes_U2 ( .ParOutRxClk(OutParDataA), 
        .SerLineXfer(SerLine2), .ParDataIn({n41, n61, n81, n693, n717, n737, 
        n761, n101, n121, n141, n161, n181, n203, n223, n243, n265, n287, n309, 
        n331, n353, n375, n397, n419, n441, n463, n485, n509, n533, n555, n579, 
        n603, n627}), .InParClk(n1060), .InParValid(n1057), .OutParClk(n1061), 
        .RxRequest(\*Logic1* ), .TxRequest(n1057), .Reset(n21) );
  INVD0 U2 ( .I(n1), .ZN(n2) );
  CKNXD16 U3 ( .I(InParDataB[12]), .ZN(n1) );
  INVD0 U4 ( .I(n3), .ZN(n4) );
  CKNXD16 U5 ( .I(InParDataB[9]), .ZN(n3) );
  INVD0 U6 ( .I(n5), .ZN(n6) );
  CKNXD16 U7 ( .I(InParDataB[6]), .ZN(n5) );
  INVD1 U8 ( .I(n2), .ZN(n332) );
  INVD1 U9 ( .I(n4), .ZN(n398) );
  INVD1 U10 ( .I(n6), .ZN(n464) );
  INVD1 U11 ( .I(n335), .ZN(n336) );
  INVD1 U12 ( .I(n333), .ZN(n334) );
  INVD1 U13 ( .I(n401), .ZN(n402) );
  INVD1 U14 ( .I(n399), .ZN(n400) );
  INVD1 U15 ( .I(n467), .ZN(n468) );
  INVD1 U16 ( .I(n465), .ZN(n466) );
  INVD1 U17 ( .I(n339), .ZN(n340) );
  INVD1 U18 ( .I(n337), .ZN(n338) );
  INVD1 U19 ( .I(n405), .ZN(n406) );
  INVD1 U20 ( .I(n403), .ZN(n404) );
  INVD1 U21 ( .I(n471), .ZN(n472) );
  INVD1 U22 ( .I(n469), .ZN(n470) );
  INVD1 U23 ( .I(n343), .ZN(n344) );
  INVD1 U24 ( .I(n341), .ZN(n342) );
  INVD1 U25 ( .I(n409), .ZN(n410) );
  INVD1 U26 ( .I(n407), .ZN(n408) );
  INVD1 U27 ( .I(n475), .ZN(n476) );
  INVD1 U28 ( .I(n473), .ZN(n474) );
  INVD1 U29 ( .I(n347), .ZN(n348) );
  INVD1 U30 ( .I(n345), .ZN(n346) );
  INVD1 U31 ( .I(n413), .ZN(n414) );
  INVD1 U32 ( .I(n411), .ZN(n412) );
  INVD1 U33 ( .I(n479), .ZN(n480) );
  INVD1 U34 ( .I(n477), .ZN(n478) );
  INVD1 U35 ( .I(n351), .ZN(n352) );
  INVD1 U36 ( .I(n349), .ZN(n350) );
  INVD1 U37 ( .I(n417), .ZN(n418) );
  INVD1 U38 ( .I(n415), .ZN(n416) );
  INVD1 U39 ( .I(n483), .ZN(n484) );
  INVD1 U40 ( .I(n481), .ZN(n482) );
  BUFFD0 U41 ( .I(Reset), .Z(n7) );
  BUFFD0 U42 ( .I(n7), .Z(n8) );
  BUFFD0 U43 ( .I(n8), .Z(n9) );
  BUFFD0 U44 ( .I(n9), .Z(n10) );
  BUFFD0 U45 ( .I(n10), .Z(n11) );
  BUFFD0 U46 ( .I(n11), .Z(n12) );
  BUFFD0 U47 ( .I(n12), .Z(n13) );
  BUFFD0 U48 ( .I(n13), .Z(n14) );
  BUFFD0 U49 ( .I(n14), .Z(n15) );
  BUFFD0 U50 ( .I(n15), .Z(n16) );
  BUFFD0 U51 ( .I(n16), .Z(n17) );
  BUFFD0 U52 ( .I(n17), .Z(n18) );
  BUFFD0 U53 ( .I(n18), .Z(n19) );
  BUFFD0 U54 ( .I(n19), .Z(n20) );
  BUFFD0 U55 ( .I(n20), .Z(n21) );
  INVD16 U56 ( .I(n629), .ZN(n630) );
  INVD16 U57 ( .I(n651), .ZN(n652) );
  INVD0 U58 ( .I(n142), .ZN(n143) );
  INVD0 U59 ( .I(n122), .ZN(n123) );
  INVD0 U60 ( .I(n204), .ZN(n205) );
  INVD0 U61 ( .I(n22), .ZN(n23) );
  CKNXD16 U62 ( .I(InParDataB[31]), .ZN(n22) );
  CKNXD0 U63 ( .I(n24), .ZN(n25) );
  CKNXD16 U64 ( .I(n23), .ZN(n24) );
  CKNXD0 U65 ( .I(n26), .ZN(n27) );
  CKNXD16 U66 ( .I(n25), .ZN(n26) );
  CKNXD0 U67 ( .I(n28), .ZN(n29) );
  CKNXD16 U68 ( .I(n27), .ZN(n28) );
  CKNXD0 U69 ( .I(n30), .ZN(n31) );
  CKNXD16 U70 ( .I(n29), .ZN(n30) );
  CKNXD0 U71 ( .I(n32), .ZN(n33) );
  CKNXD16 U72 ( .I(n31), .ZN(n32) );
  CKNXD0 U73 ( .I(n34), .ZN(n35) );
  CKNXD16 U74 ( .I(n33), .ZN(n34) );
  CKNXD0 U75 ( .I(n40), .ZN(n41) );
  INVD0 U76 ( .I(n36), .ZN(n37) );
  CKNXD16 U77 ( .I(n35), .ZN(n36) );
  CKNXD0 U78 ( .I(n38), .ZN(n39) );
  CKNXD16 U79 ( .I(n37), .ZN(n38) );
  CKNXD16 U80 ( .I(n39), .ZN(n40) );
  CKNXD0 U81 ( .I(n56), .ZN(n57) );
  CKNXD0 U82 ( .I(n42), .ZN(n43) );
  CKNXD16 U83 ( .I(InParDataB[30]), .ZN(n42) );
  CKNXD0 U84 ( .I(n44), .ZN(n45) );
  CKNXD16 U85 ( .I(n43), .ZN(n44) );
  CKNXD0 U86 ( .I(n46), .ZN(n47) );
  CKNXD16 U87 ( .I(n45), .ZN(n46) );
  CKNXD0 U88 ( .I(n48), .ZN(n49) );
  CKNXD16 U89 ( .I(n47), .ZN(n48) );
  CKNXD0 U90 ( .I(n50), .ZN(n51) );
  CKNXD16 U91 ( .I(n49), .ZN(n50) );
  CKNXD0 U92 ( .I(n52), .ZN(n53) );
  CKNXD16 U93 ( .I(n51), .ZN(n52) );
  CKNXD0 U94 ( .I(n54), .ZN(n55) );
  CKNXD16 U95 ( .I(n53), .ZN(n54) );
  CKNXD0 U96 ( .I(n60), .ZN(n61) );
  CKNXD16 U97 ( .I(n55), .ZN(n56) );
  CKNXD0 U98 ( .I(n58), .ZN(n59) );
  CKNXD16 U99 ( .I(n57), .ZN(n58) );
  CKNXD16 U100 ( .I(n59), .ZN(n60) );
  CKNXD0 U101 ( .I(n76), .ZN(n77) );
  CKNXD0 U102 ( .I(n62), .ZN(n63) );
  CKNXD16 U103 ( .I(InParDataB[29]), .ZN(n62) );
  CKNXD0 U104 ( .I(n64), .ZN(n65) );
  CKNXD16 U105 ( .I(n63), .ZN(n64) );
  CKNXD0 U106 ( .I(n66), .ZN(n67) );
  CKNXD16 U107 ( .I(n65), .ZN(n66) );
  CKNXD0 U108 ( .I(n68), .ZN(n69) );
  CKNXD16 U109 ( .I(n67), .ZN(n68) );
  CKNXD0 U110 ( .I(n70), .ZN(n71) );
  CKNXD16 U111 ( .I(n69), .ZN(n70) );
  CKNXD0 U112 ( .I(n72), .ZN(n73) );
  CKNXD16 U113 ( .I(n71), .ZN(n72) );
  CKNXD0 U114 ( .I(n74), .ZN(n75) );
  CKNXD16 U115 ( .I(n73), .ZN(n74) );
  CKNXD0 U116 ( .I(n80), .ZN(n81) );
  CKNXD16 U117 ( .I(n75), .ZN(n76) );
  CKNXD0 U118 ( .I(n78), .ZN(n79) );
  CKNXD16 U119 ( .I(n77), .ZN(n78) );
  CKNXD16 U120 ( .I(n79), .ZN(n80) );
  INVD0 U121 ( .I(n82), .ZN(n83) );
  CKNXD16 U122 ( .I(InParDataB[24]), .ZN(n82) );
  CKNXD0 U123 ( .I(n84), .ZN(n85) );
  CKNXD16 U124 ( .I(n83), .ZN(n84) );
  CKNXD0 U125 ( .I(n86), .ZN(n87) );
  CKNXD16 U126 ( .I(n85), .ZN(n86) );
  CKNXD0 U127 ( .I(n88), .ZN(n89) );
  CKNXD16 U128 ( .I(n87), .ZN(n88) );
  CKNXD0 U129 ( .I(n90), .ZN(n91) );
  CKNXD16 U130 ( .I(n89), .ZN(n90) );
  CKNXD0 U131 ( .I(n92), .ZN(n93) );
  CKNXD16 U132 ( .I(n91), .ZN(n92) );
  CKNXD0 U133 ( .I(n94), .ZN(n95) );
  CKNXD16 U134 ( .I(n93), .ZN(n94) );
  CKNXD0 U135 ( .I(n100), .ZN(n101) );
  INVD0 U136 ( .I(n96), .ZN(n97) );
  CKNXD16 U137 ( .I(n95), .ZN(n96) );
  CKNXD0 U138 ( .I(n98), .ZN(n99) );
  CKNXD16 U139 ( .I(n97), .ZN(n98) );
  CKNXD16 U140 ( .I(n99), .ZN(n100) );
  INVD0 U141 ( .I(n102), .ZN(n103) );
  CKNXD16 U142 ( .I(InParDataB[23]), .ZN(n102) );
  CKNXD0 U143 ( .I(n104), .ZN(n105) );
  CKNXD16 U144 ( .I(n103), .ZN(n104) );
  CKNXD0 U145 ( .I(n106), .ZN(n107) );
  CKNXD16 U146 ( .I(n105), .ZN(n106) );
  CKNXD0 U147 ( .I(n108), .ZN(n109) );
  CKNXD16 U148 ( .I(n107), .ZN(n108) );
  CKNXD0 U149 ( .I(n110), .ZN(n111) );
  CKNXD16 U150 ( .I(n109), .ZN(n110) );
  CKNXD0 U151 ( .I(n112), .ZN(n113) );
  CKNXD16 U152 ( .I(n111), .ZN(n112) );
  CKNXD0 U153 ( .I(n114), .ZN(n115) );
  CKNXD16 U154 ( .I(n113), .ZN(n114) );
  CKNXD0 U155 ( .I(n120), .ZN(n121) );
  INVD0 U156 ( .I(n116), .ZN(n117) );
  CKNXD16 U157 ( .I(n115), .ZN(n116) );
  CKNXD0 U158 ( .I(n118), .ZN(n119) );
  CKNXD16 U159 ( .I(n117), .ZN(n118) );
  CKNXD16 U160 ( .I(n119), .ZN(n120) );
  CKNXD0 U161 ( .I(n136), .ZN(n137) );
  CKNXD16 U162 ( .I(InParDataB[22]), .ZN(n122) );
  CKNXD0 U163 ( .I(n124), .ZN(n125) );
  CKNXD16 U164 ( .I(n123), .ZN(n124) );
  CKNXD0 U165 ( .I(n126), .ZN(n127) );
  CKNXD16 U166 ( .I(n125), .ZN(n126) );
  CKNXD0 U167 ( .I(n128), .ZN(n129) );
  CKNXD16 U168 ( .I(n127), .ZN(n128) );
  CKNXD0 U169 ( .I(n130), .ZN(n131) );
  CKNXD16 U170 ( .I(n129), .ZN(n130) );
  CKNXD0 U171 ( .I(n132), .ZN(n133) );
  CKNXD16 U172 ( .I(n131), .ZN(n132) );
  CKNXD0 U173 ( .I(n134), .ZN(n135) );
  CKNXD16 U174 ( .I(n133), .ZN(n134) );
  CKNXD0 U175 ( .I(n140), .ZN(n141) );
  CKNXD16 U176 ( .I(n135), .ZN(n136) );
  CKNXD0 U177 ( .I(n138), .ZN(n139) );
  CKNXD16 U178 ( .I(n137), .ZN(n138) );
  CKNXD16 U179 ( .I(n139), .ZN(n140) );
  CKNXD0 U180 ( .I(n156), .ZN(n157) );
  CKNXD16 U181 ( .I(InParDataB[21]), .ZN(n142) );
  CKNXD0 U182 ( .I(n144), .ZN(n145) );
  CKNXD16 U183 ( .I(n143), .ZN(n144) );
  CKNXD0 U184 ( .I(n146), .ZN(n147) );
  CKNXD16 U185 ( .I(n145), .ZN(n146) );
  CKNXD0 U186 ( .I(n148), .ZN(n149) );
  CKNXD16 U187 ( .I(n147), .ZN(n148) );
  CKNXD0 U188 ( .I(n150), .ZN(n151) );
  CKNXD16 U189 ( .I(n149), .ZN(n150) );
  CKNXD0 U190 ( .I(n152), .ZN(n153) );
  CKNXD16 U191 ( .I(n151), .ZN(n152) );
  CKNXD0 U192 ( .I(n154), .ZN(n155) );
  CKNXD16 U193 ( .I(n153), .ZN(n154) );
  CKNXD0 U194 ( .I(n160), .ZN(n161) );
  CKNXD16 U195 ( .I(n155), .ZN(n156) );
  CKNXD0 U196 ( .I(n158), .ZN(n159) );
  CKNXD16 U197 ( .I(n157), .ZN(n158) );
  CKNXD16 U198 ( .I(n159), .ZN(n160) );
  INVD0 U199 ( .I(n162), .ZN(n163) );
  CKNXD16 U200 ( .I(InParDataB[20]), .ZN(n162) );
  CKNXD0 U201 ( .I(n164), .ZN(n165) );
  CKNXD16 U202 ( .I(n163), .ZN(n164) );
  CKNXD0 U203 ( .I(n166), .ZN(n167) );
  CKNXD16 U204 ( .I(n165), .ZN(n166) );
  CKNXD0 U205 ( .I(n168), .ZN(n169) );
  CKNXD16 U206 ( .I(n167), .ZN(n168) );
  CKNXD0 U207 ( .I(n170), .ZN(n171) );
  CKNXD16 U208 ( .I(n169), .ZN(n170) );
  CKNXD0 U209 ( .I(n172), .ZN(n173) );
  CKNXD16 U210 ( .I(n171), .ZN(n172) );
  CKNXD0 U211 ( .I(n174), .ZN(n175) );
  CKNXD16 U212 ( .I(n173), .ZN(n174) );
  CKNXD0 U213 ( .I(n180), .ZN(n181) );
  INVD0 U214 ( .I(n176), .ZN(n177) );
  CKNXD16 U215 ( .I(n175), .ZN(n176) );
  CKNXD0 U216 ( .I(n178), .ZN(n179) );
  CKNXD16 U217 ( .I(n177), .ZN(n178) );
  CKNXD16 U218 ( .I(n179), .ZN(n180) );
  CKNXD0 U219 ( .I(n182), .ZN(n183) );
  CKNXD16 U220 ( .I(InParDataB[19]), .ZN(n182) );
  INVD0 U221 ( .I(n184), .ZN(n185) );
  CKNXD16 U222 ( .I(n183), .ZN(n184) );
  CKNXD0 U223 ( .I(n186), .ZN(n187) );
  CKNXD16 U224 ( .I(n185), .ZN(n186) );
  CKNXD0 U225 ( .I(n188), .ZN(n189) );
  CKNXD16 U226 ( .I(n187), .ZN(n188) );
  CKNXD0 U227 ( .I(n190), .ZN(n191) );
  CKNXD16 U228 ( .I(n189), .ZN(n190) );
  CKNXD0 U229 ( .I(n192), .ZN(n193) );
  CKNXD16 U230 ( .I(n191), .ZN(n192) );
  CKNXD0 U231 ( .I(n194), .ZN(n195) );
  CKNXD16 U232 ( .I(n193), .ZN(n194) );
  CKNXD0 U233 ( .I(n196), .ZN(n197) );
  CKNXD16 U234 ( .I(n195), .ZN(n196) );
  CKNXD0 U235 ( .I(n202), .ZN(n203) );
  INVD0 U236 ( .I(n198), .ZN(n199) );
  CKNXD16 U237 ( .I(n197), .ZN(n198) );
  CKNXD0 U238 ( .I(n200), .ZN(n201) );
  CKNXD16 U239 ( .I(n199), .ZN(n200) );
  CKNXD16 U240 ( .I(n201), .ZN(n202) );
  CKNXD0 U241 ( .I(n218), .ZN(n219) );
  CKNXD16 U242 ( .I(InParDataB[18]), .ZN(n204) );
  CKNXD0 U243 ( .I(n206), .ZN(n207) );
  CKNXD16 U244 ( .I(n205), .ZN(n206) );
  CKNXD0 U245 ( .I(n208), .ZN(n209) );
  CKNXD16 U246 ( .I(n207), .ZN(n208) );
  CKNXD0 U247 ( .I(n210), .ZN(n211) );
  CKNXD16 U248 ( .I(n209), .ZN(n210) );
  CKNXD0 U249 ( .I(n212), .ZN(n213) );
  CKNXD16 U250 ( .I(n211), .ZN(n212) );
  CKNXD0 U251 ( .I(n214), .ZN(n215) );
  CKNXD16 U252 ( .I(n213), .ZN(n214) );
  CKNXD0 U253 ( .I(n216), .ZN(n217) );
  CKNXD16 U254 ( .I(n215), .ZN(n216) );
  CKNXD0 U255 ( .I(n222), .ZN(n223) );
  CKNXD16 U256 ( .I(n217), .ZN(n218) );
  CKNXD0 U257 ( .I(n220), .ZN(n221) );
  CKNXD16 U258 ( .I(n219), .ZN(n220) );
  CKNXD16 U259 ( .I(n221), .ZN(n222) );
  CKNXD0 U260 ( .I(n238), .ZN(n239) );
  CKNXD0 U261 ( .I(n224), .ZN(n225) );
  CKNXD16 U262 ( .I(InParDataB[17]), .ZN(n224) );
  CKNXD0 U263 ( .I(n226), .ZN(n227) );
  CKNXD16 U264 ( .I(n225), .ZN(n226) );
  CKNXD0 U265 ( .I(n228), .ZN(n229) );
  CKNXD16 U266 ( .I(n227), .ZN(n228) );
  CKNXD0 U267 ( .I(n230), .ZN(n231) );
  CKNXD16 U268 ( .I(n229), .ZN(n230) );
  CKNXD0 U269 ( .I(n232), .ZN(n233) );
  CKNXD16 U270 ( .I(n231), .ZN(n232) );
  CKNXD0 U271 ( .I(n234), .ZN(n235) );
  CKNXD16 U272 ( .I(n233), .ZN(n234) );
  CKNXD0 U273 ( .I(n236), .ZN(n237) );
  CKNXD16 U274 ( .I(n235), .ZN(n236) );
  CKNXD0 U275 ( .I(n242), .ZN(n243) );
  CKNXD16 U276 ( .I(n237), .ZN(n238) );
  CKNXD0 U277 ( .I(n240), .ZN(n241) );
  CKNXD16 U278 ( .I(n239), .ZN(n240) );
  CKNXD16 U279 ( .I(n241), .ZN(n242) );
  CKNXD0 U280 ( .I(n244), .ZN(n245) );
  CKNXD16 U281 ( .I(InParDataB[16]), .ZN(n244) );
  INVD0 U282 ( .I(n246), .ZN(n247) );
  CKNXD16 U283 ( .I(n245), .ZN(n246) );
  CKNXD0 U284 ( .I(n248), .ZN(n249) );
  CKNXD16 U285 ( .I(n247), .ZN(n248) );
  CKNXD0 U286 ( .I(n250), .ZN(n251) );
  CKNXD16 U287 ( .I(n249), .ZN(n250) );
  CKNXD0 U288 ( .I(n252), .ZN(n253) );
  CKNXD16 U289 ( .I(n251), .ZN(n252) );
  CKNXD0 U290 ( .I(n254), .ZN(n255) );
  CKNXD16 U291 ( .I(n253), .ZN(n254) );
  CKNXD0 U292 ( .I(n256), .ZN(n257) );
  CKNXD16 U293 ( .I(n255), .ZN(n256) );
  CKNXD0 U294 ( .I(n258), .ZN(n259) );
  CKNXD16 U295 ( .I(n257), .ZN(n258) );
  CKNXD0 U296 ( .I(n264), .ZN(n265) );
  INVD0 U297 ( .I(n260), .ZN(n261) );
  CKNXD16 U298 ( .I(n259), .ZN(n260) );
  CKNXD0 U299 ( .I(n262), .ZN(n263) );
  CKNXD16 U300 ( .I(n261), .ZN(n262) );
  CKNXD16 U301 ( .I(n263), .ZN(n264) );
  CKNXD0 U302 ( .I(n268), .ZN(n269) );
  INVD0 U303 ( .I(n266), .ZN(n267) );
  CKNXD16 U304 ( .I(InParDataB[15]), .ZN(n266) );
  CKNXD16 U305 ( .I(n267), .ZN(n268) );
  CKNXD0 U306 ( .I(n270), .ZN(n271) );
  CKNXD16 U307 ( .I(n269), .ZN(n270) );
  CKNXD0 U308 ( .I(n272), .ZN(n273) );
  CKNXD16 U309 ( .I(n271), .ZN(n272) );
  CKNXD0 U310 ( .I(n274), .ZN(n275) );
  CKNXD16 U311 ( .I(n273), .ZN(n274) );
  CKNXD0 U312 ( .I(n276), .ZN(n277) );
  CKNXD16 U313 ( .I(n275), .ZN(n276) );
  CKNXD0 U314 ( .I(n278), .ZN(n279) );
  CKNXD16 U315 ( .I(n277), .ZN(n278) );
  CKNXD0 U316 ( .I(n280), .ZN(n281) );
  CKNXD16 U317 ( .I(n279), .ZN(n280) );
  CKNXD0 U318 ( .I(n286), .ZN(n287) );
  INVD0 U319 ( .I(n282), .ZN(n283) );
  CKNXD16 U320 ( .I(n281), .ZN(n282) );
  CKNXD0 U321 ( .I(n284), .ZN(n285) );
  CKNXD16 U322 ( .I(n283), .ZN(n284) );
  CKNXD16 U323 ( .I(n285), .ZN(n286) );
  CKNXD0 U324 ( .I(n290), .ZN(n291) );
  INVD0 U325 ( .I(n288), .ZN(n289) );
  CKNXD16 U326 ( .I(InParDataB[14]), .ZN(n288) );
  CKNXD16 U327 ( .I(n289), .ZN(n290) );
  CKNXD0 U328 ( .I(n292), .ZN(n293) );
  CKNXD16 U329 ( .I(n291), .ZN(n292) );
  CKNXD0 U330 ( .I(n294), .ZN(n295) );
  CKNXD16 U331 ( .I(n293), .ZN(n294) );
  CKNXD0 U332 ( .I(n296), .ZN(n297) );
  CKNXD16 U333 ( .I(n295), .ZN(n296) );
  CKNXD0 U334 ( .I(n298), .ZN(n299) );
  CKNXD16 U335 ( .I(n297), .ZN(n298) );
  CKNXD0 U336 ( .I(n300), .ZN(n301) );
  CKNXD16 U337 ( .I(n299), .ZN(n300) );
  CKNXD0 U338 ( .I(n302), .ZN(n303) );
  CKNXD16 U339 ( .I(n301), .ZN(n302) );
  CKNXD0 U340 ( .I(n308), .ZN(n309) );
  INVD0 U341 ( .I(n304), .ZN(n305) );
  CKNXD16 U342 ( .I(n303), .ZN(n304) );
  CKNXD0 U343 ( .I(n306), .ZN(n307) );
  CKNXD16 U344 ( .I(n305), .ZN(n306) );
  CKNXD16 U345 ( .I(n307), .ZN(n308) );
  CKNXD0 U346 ( .I(n310), .ZN(n311) );
  CKNXD16 U347 ( .I(InParDataB[13]), .ZN(n310) );
  INVD0 U348 ( .I(n312), .ZN(n313) );
  CKNXD16 U349 ( .I(n311), .ZN(n312) );
  CKNXD0 U350 ( .I(n314), .ZN(n315) );
  CKNXD16 U351 ( .I(n313), .ZN(n314) );
  CKNXD0 U352 ( .I(n316), .ZN(n317) );
  CKNXD16 U353 ( .I(n315), .ZN(n316) );
  CKNXD0 U354 ( .I(n318), .ZN(n319) );
  CKNXD16 U355 ( .I(n317), .ZN(n318) );
  CKNXD0 U356 ( .I(n320), .ZN(n321) );
  CKNXD16 U357 ( .I(n319), .ZN(n320) );
  CKNXD0 U358 ( .I(n322), .ZN(n323) );
  CKNXD16 U359 ( .I(n321), .ZN(n322) );
  CKNXD0 U360 ( .I(n324), .ZN(n325) );
  CKNXD16 U361 ( .I(n323), .ZN(n324) );
  CKNXD0 U362 ( .I(n330), .ZN(n331) );
  INVD0 U363 ( .I(n326), .ZN(n327) );
  CKNXD16 U364 ( .I(n325), .ZN(n326) );
  CKNXD0 U365 ( .I(n328), .ZN(n329) );
  CKNXD16 U366 ( .I(n327), .ZN(n328) );
  CKNXD16 U367 ( .I(n329), .ZN(n330) );
  CKNXD0 U368 ( .I(n332), .ZN(n333) );
  INVD0 U369 ( .I(n334), .ZN(n335) );
  CKNXD0 U370 ( .I(n336), .ZN(n337) );
  CKNXD0 U371 ( .I(n338), .ZN(n339) );
  CKNXD0 U372 ( .I(n340), .ZN(n341) );
  CKNXD0 U373 ( .I(n342), .ZN(n343) );
  CKNXD0 U374 ( .I(n344), .ZN(n345) );
  CKNXD0 U375 ( .I(n346), .ZN(n347) );
  CKNXD0 U376 ( .I(n352), .ZN(n353) );
  INVD0 U377 ( .I(n348), .ZN(n349) );
  CKNXD0 U378 ( .I(n350), .ZN(n351) );
  CKNXD0 U379 ( .I(n356), .ZN(n357) );
  INVD0 U380 ( .I(n354), .ZN(n355) );
  CKNXD16 U381 ( .I(InParDataB[11]), .ZN(n354) );
  CKNXD16 U382 ( .I(n355), .ZN(n356) );
  CKNXD0 U383 ( .I(n358), .ZN(n359) );
  CKNXD16 U384 ( .I(n357), .ZN(n358) );
  CKNXD0 U385 ( .I(n360), .ZN(n361) );
  CKNXD16 U386 ( .I(n359), .ZN(n360) );
  CKNXD0 U387 ( .I(n362), .ZN(n363) );
  CKNXD16 U388 ( .I(n361), .ZN(n362) );
  CKNXD0 U389 ( .I(n364), .ZN(n365) );
  CKNXD16 U390 ( .I(n363), .ZN(n364) );
  CKNXD0 U391 ( .I(n366), .ZN(n367) );
  CKNXD16 U392 ( .I(n365), .ZN(n366) );
  CKNXD0 U393 ( .I(n368), .ZN(n369) );
  CKNXD16 U394 ( .I(n367), .ZN(n368) );
  CKNXD0 U395 ( .I(n374), .ZN(n375) );
  INVD0 U396 ( .I(n370), .ZN(n371) );
  CKNXD16 U397 ( .I(n369), .ZN(n370) );
  CKNXD0 U398 ( .I(n372), .ZN(n373) );
  CKNXD16 U399 ( .I(n371), .ZN(n372) );
  CKNXD16 U400 ( .I(n373), .ZN(n374) );
  CKNXD0 U401 ( .I(n378), .ZN(n379) );
  INVD0 U402 ( .I(n376), .ZN(n377) );
  CKNXD16 U403 ( .I(InParDataB[10]), .ZN(n376) );
  CKNXD16 U404 ( .I(n377), .ZN(n378) );
  CKNXD0 U405 ( .I(n380), .ZN(n381) );
  CKNXD16 U406 ( .I(n379), .ZN(n380) );
  CKNXD0 U407 ( .I(n382), .ZN(n383) );
  CKNXD16 U408 ( .I(n381), .ZN(n382) );
  CKNXD0 U409 ( .I(n384), .ZN(n385) );
  CKNXD16 U410 ( .I(n383), .ZN(n384) );
  CKNXD0 U411 ( .I(n386), .ZN(n387) );
  CKNXD16 U412 ( .I(n385), .ZN(n386) );
  CKNXD0 U413 ( .I(n388), .ZN(n389) );
  CKNXD16 U414 ( .I(n387), .ZN(n388) );
  CKNXD0 U415 ( .I(n390), .ZN(n391) );
  CKNXD16 U416 ( .I(n389), .ZN(n390) );
  CKNXD0 U417 ( .I(n396), .ZN(n397) );
  INVD0 U418 ( .I(n392), .ZN(n393) );
  CKNXD16 U419 ( .I(n391), .ZN(n392) );
  CKNXD0 U420 ( .I(n394), .ZN(n395) );
  CKNXD16 U421 ( .I(n393), .ZN(n394) );
  CKNXD16 U422 ( .I(n395), .ZN(n396) );
  CKNXD0 U423 ( .I(n398), .ZN(n399) );
  INVD0 U424 ( .I(n400), .ZN(n401) );
  CKNXD0 U425 ( .I(n402), .ZN(n403) );
  CKNXD0 U426 ( .I(n404), .ZN(n405) );
  CKNXD0 U427 ( .I(n406), .ZN(n407) );
  CKNXD0 U428 ( .I(n408), .ZN(n409) );
  CKNXD0 U429 ( .I(n410), .ZN(n411) );
  CKNXD0 U430 ( .I(n412), .ZN(n413) );
  CKNXD0 U431 ( .I(n418), .ZN(n419) );
  INVD0 U432 ( .I(n414), .ZN(n415) );
  CKNXD0 U433 ( .I(n416), .ZN(n417) );
  CKNXD0 U434 ( .I(n422), .ZN(n423) );
  INVD0 U435 ( .I(n420), .ZN(n421) );
  CKNXD16 U436 ( .I(InParDataB[8]), .ZN(n420) );
  CKNXD16 U437 ( .I(n421), .ZN(n422) );
  CKNXD0 U438 ( .I(n424), .ZN(n425) );
  CKNXD16 U439 ( .I(n423), .ZN(n424) );
  CKNXD0 U440 ( .I(n426), .ZN(n427) );
  CKNXD16 U441 ( .I(n425), .ZN(n426) );
  CKNXD0 U442 ( .I(n428), .ZN(n429) );
  CKNXD16 U443 ( .I(n427), .ZN(n428) );
  CKNXD0 U444 ( .I(n430), .ZN(n431) );
  CKNXD16 U445 ( .I(n429), .ZN(n430) );
  CKNXD0 U446 ( .I(n432), .ZN(n433) );
  CKNXD16 U447 ( .I(n431), .ZN(n432) );
  CKNXD0 U448 ( .I(n434), .ZN(n435) );
  CKNXD16 U449 ( .I(n433), .ZN(n434) );
  CKNXD0 U450 ( .I(n440), .ZN(n441) );
  INVD0 U451 ( .I(n436), .ZN(n437) );
  CKNXD16 U452 ( .I(n435), .ZN(n436) );
  CKNXD0 U453 ( .I(n438), .ZN(n439) );
  CKNXD16 U454 ( .I(n437), .ZN(n438) );
  CKNXD16 U455 ( .I(n439), .ZN(n440) );
  CKNXD0 U456 ( .I(n444), .ZN(n445) );
  INVD0 U457 ( .I(n442), .ZN(n443) );
  CKNXD16 U458 ( .I(InParDataB[7]), .ZN(n442) );
  CKNXD16 U459 ( .I(n443), .ZN(n444) );
  CKNXD0 U460 ( .I(n446), .ZN(n447) );
  CKNXD16 U461 ( .I(n445), .ZN(n446) );
  CKNXD0 U462 ( .I(n448), .ZN(n449) );
  CKNXD16 U463 ( .I(n447), .ZN(n448) );
  CKNXD0 U464 ( .I(n450), .ZN(n451) );
  CKNXD16 U465 ( .I(n449), .ZN(n450) );
  CKNXD0 U466 ( .I(n452), .ZN(n453) );
  CKNXD16 U467 ( .I(n451), .ZN(n452) );
  CKNXD0 U468 ( .I(n454), .ZN(n455) );
  CKNXD16 U469 ( .I(n453), .ZN(n454) );
  CKNXD0 U470 ( .I(n456), .ZN(n457) );
  CKNXD16 U471 ( .I(n455), .ZN(n456) );
  CKNXD0 U472 ( .I(n462), .ZN(n463) );
  INVD0 U473 ( .I(n458), .ZN(n459) );
  CKNXD16 U474 ( .I(n457), .ZN(n458) );
  CKNXD0 U475 ( .I(n460), .ZN(n461) );
  CKNXD16 U476 ( .I(n459), .ZN(n460) );
  CKNXD16 U477 ( .I(n461), .ZN(n462) );
  CKNXD0 U478 ( .I(n464), .ZN(n465) );
  INVD0 U479 ( .I(n466), .ZN(n467) );
  CKNXD0 U480 ( .I(n468), .ZN(n469) );
  CKNXD0 U481 ( .I(n470), .ZN(n471) );
  CKNXD0 U482 ( .I(n472), .ZN(n473) );
  CKNXD0 U483 ( .I(n474), .ZN(n475) );
  CKNXD0 U484 ( .I(n476), .ZN(n477) );
  CKNXD0 U485 ( .I(n478), .ZN(n479) );
  CKNXD0 U486 ( .I(n484), .ZN(n485) );
  INVD0 U487 ( .I(n480), .ZN(n481) );
  CKNXD0 U488 ( .I(n482), .ZN(n483) );
  CKNXD0 U489 ( .I(n486), .ZN(n487) );
  CKNXD16 U490 ( .I(InParDataB[5]), .ZN(n486) );
  CKNXD0 U491 ( .I(n488), .ZN(n489) );
  CKNXD16 U492 ( .I(n487), .ZN(n488) );
  INVD0 U493 ( .I(n490), .ZN(n491) );
  CKNXD16 U494 ( .I(n489), .ZN(n490) );
  CKNXD0 U495 ( .I(n492), .ZN(n493) );
  CKNXD16 U496 ( .I(n491), .ZN(n492) );
  CKNXD0 U497 ( .I(n494), .ZN(n495) );
  CKNXD16 U498 ( .I(n493), .ZN(n494) );
  CKNXD0 U499 ( .I(n496), .ZN(n497) );
  CKNXD16 U500 ( .I(n495), .ZN(n496) );
  CKNXD0 U501 ( .I(n498), .ZN(n499) );
  CKNXD16 U502 ( .I(n497), .ZN(n498) );
  CKNXD0 U503 ( .I(n500), .ZN(n501) );
  CKNXD16 U504 ( .I(n499), .ZN(n500) );
  CKNXD0 U505 ( .I(n502), .ZN(n503) );
  CKNXD16 U506 ( .I(n501), .ZN(n502) );
  CKNXD0 U507 ( .I(n508), .ZN(n509) );
  INVD0 U508 ( .I(n504), .ZN(n505) );
  CKNXD16 U509 ( .I(n503), .ZN(n504) );
  CKNXD0 U510 ( .I(n506), .ZN(n507) );
  CKNXD16 U511 ( .I(n505), .ZN(n506) );
  CKNXD16 U512 ( .I(n507), .ZN(n508) );
  CKNXD0 U513 ( .I(n514), .ZN(n515) );
  INVD0 U514 ( .I(n510), .ZN(n511) );
  CKNXD16 U515 ( .I(InParDataB[4]), .ZN(n510) );
  CKNXD0 U516 ( .I(n512), .ZN(n513) );
  CKNXD16 U517 ( .I(n511), .ZN(n512) );
  CKNXD16 U518 ( .I(n513), .ZN(n514) );
  CKNXD0 U519 ( .I(n516), .ZN(n517) );
  CKNXD16 U520 ( .I(n515), .ZN(n516) );
  CKNXD0 U521 ( .I(n518), .ZN(n519) );
  CKNXD16 U522 ( .I(n517), .ZN(n518) );
  CKNXD0 U523 ( .I(n520), .ZN(n521) );
  CKNXD16 U524 ( .I(n519), .ZN(n520) );
  CKNXD0 U525 ( .I(n522), .ZN(n523) );
  CKNXD16 U526 ( .I(n521), .ZN(n522) );
  CKNXD0 U527 ( .I(n524), .ZN(n525) );
  CKNXD16 U528 ( .I(n523), .ZN(n524) );
  CKNXD0 U529 ( .I(n526), .ZN(n527) );
  CKNXD16 U530 ( .I(n525), .ZN(n526) );
  CKNXD0 U531 ( .I(n532), .ZN(n533) );
  INVD0 U532 ( .I(n528), .ZN(n529) );
  CKNXD16 U533 ( .I(n527), .ZN(n528) );
  CKNXD0 U534 ( .I(n530), .ZN(n531) );
  CKNXD16 U535 ( .I(n529), .ZN(n530) );
  CKNXD16 U536 ( .I(n531), .ZN(n532) );
  CKNXD0 U537 ( .I(n536), .ZN(n537) );
  INVD0 U538 ( .I(n534), .ZN(n535) );
  CKNXD16 U539 ( .I(InParDataB[3]), .ZN(n534) );
  CKNXD16 U540 ( .I(n535), .ZN(n536) );
  CKNXD0 U541 ( .I(n538), .ZN(n539) );
  CKNXD16 U542 ( .I(n537), .ZN(n538) );
  CKNXD0 U543 ( .I(n540), .ZN(n541) );
  CKNXD16 U544 ( .I(n539), .ZN(n540) );
  CKNXD0 U545 ( .I(n542), .ZN(n543) );
  CKNXD16 U546 ( .I(n541), .ZN(n542) );
  CKNXD0 U547 ( .I(n544), .ZN(n545) );
  CKNXD16 U548 ( .I(n543), .ZN(n544) );
  CKNXD0 U549 ( .I(n546), .ZN(n547) );
  CKNXD16 U550 ( .I(n545), .ZN(n546) );
  CKNXD0 U551 ( .I(n548), .ZN(n549) );
  CKNXD16 U552 ( .I(n547), .ZN(n548) );
  CKNXD0 U553 ( .I(n554), .ZN(n555) );
  INVD0 U554 ( .I(n550), .ZN(n551) );
  CKNXD16 U555 ( .I(n549), .ZN(n550) );
  CKNXD0 U556 ( .I(n552), .ZN(n553) );
  CKNXD16 U557 ( .I(n551), .ZN(n552) );
  CKNXD16 U558 ( .I(n553), .ZN(n554) );
  CKNXD0 U559 ( .I(n556), .ZN(n557) );
  CKNXD16 U560 ( .I(InParDataB[2]), .ZN(n556) );
  CKNXD0 U561 ( .I(n558), .ZN(n559) );
  CKNXD16 U562 ( .I(n557), .ZN(n558) );
  INVD0 U563 ( .I(n560), .ZN(n561) );
  CKNXD16 U564 ( .I(n559), .ZN(n560) );
  CKNXD0 U565 ( .I(n562), .ZN(n563) );
  CKNXD16 U566 ( .I(n561), .ZN(n562) );
  CKNXD0 U567 ( .I(n564), .ZN(n565) );
  CKNXD16 U568 ( .I(n563), .ZN(n564) );
  CKNXD0 U569 ( .I(n566), .ZN(n567) );
  CKNXD16 U570 ( .I(n565), .ZN(n566) );
  CKNXD0 U571 ( .I(n568), .ZN(n569) );
  CKNXD16 U572 ( .I(n567), .ZN(n568) );
  CKNXD0 U573 ( .I(n570), .ZN(n571) );
  CKNXD16 U574 ( .I(n569), .ZN(n570) );
  CKNXD0 U575 ( .I(n572), .ZN(n573) );
  CKNXD16 U576 ( .I(n571), .ZN(n572) );
  CKNXD0 U577 ( .I(n578), .ZN(n579) );
  INVD0 U578 ( .I(n574), .ZN(n575) );
  CKNXD16 U579 ( .I(n573), .ZN(n574) );
  CKNXD0 U580 ( .I(n576), .ZN(n577) );
  CKNXD16 U581 ( .I(n575), .ZN(n576) );
  CKNXD16 U582 ( .I(n577), .ZN(n578) );
  CKNXD0 U583 ( .I(n580), .ZN(n581) );
  CKNXD16 U584 ( .I(InParDataB[1]), .ZN(n580) );
  CKNXD0 U585 ( .I(n582), .ZN(n583) );
  CKNXD16 U586 ( .I(n581), .ZN(n582) );
  INVD0 U587 ( .I(n584), .ZN(n585) );
  CKNXD16 U588 ( .I(n583), .ZN(n584) );
  CKNXD0 U589 ( .I(n586), .ZN(n587) );
  CKNXD16 U590 ( .I(n585), .ZN(n586) );
  CKNXD0 U591 ( .I(n588), .ZN(n589) );
  CKNXD16 U592 ( .I(n587), .ZN(n588) );
  CKNXD0 U593 ( .I(n590), .ZN(n591) );
  CKNXD16 U594 ( .I(n589), .ZN(n590) );
  CKNXD0 U595 ( .I(n592), .ZN(n593) );
  CKNXD16 U596 ( .I(n591), .ZN(n592) );
  CKNXD0 U597 ( .I(n594), .ZN(n595) );
  CKNXD16 U598 ( .I(n593), .ZN(n594) );
  CKNXD0 U599 ( .I(n596), .ZN(n597) );
  CKNXD16 U600 ( .I(n595), .ZN(n596) );
  CKNXD0 U601 ( .I(n602), .ZN(n603) );
  INVD0 U602 ( .I(n598), .ZN(n599) );
  CKNXD16 U603 ( .I(n597), .ZN(n598) );
  CKNXD0 U604 ( .I(n600), .ZN(n601) );
  CKNXD16 U605 ( .I(n599), .ZN(n600) );
  CKNXD16 U606 ( .I(n601), .ZN(n602) );
  CKNXD0 U607 ( .I(n604), .ZN(n605) );
  CKNXD16 U608 ( .I(InParDataB[0]), .ZN(n604) );
  CKNXD0 U609 ( .I(n606), .ZN(n607) );
  CKNXD16 U610 ( .I(n605), .ZN(n606) );
  INVD0 U611 ( .I(n608), .ZN(n609) );
  CKNXD16 U612 ( .I(n607), .ZN(n608) );
  CKNXD0 U613 ( .I(n610), .ZN(n611) );
  CKNXD16 U614 ( .I(n609), .ZN(n610) );
  CKNXD0 U615 ( .I(n612), .ZN(n613) );
  CKNXD16 U616 ( .I(n611), .ZN(n612) );
  CKNXD0 U617 ( .I(n614), .ZN(n615) );
  CKNXD16 U618 ( .I(n613), .ZN(n614) );
  CKNXD0 U619 ( .I(n616), .ZN(n617) );
  CKNXD16 U620 ( .I(n615), .ZN(n616) );
  CKNXD0 U621 ( .I(n618), .ZN(n619) );
  CKNXD16 U622 ( .I(n617), .ZN(n618) );
  CKNXD0 U623 ( .I(n620), .ZN(n621) );
  CKNXD16 U624 ( .I(n619), .ZN(n620) );
  CKNXD0 U625 ( .I(n626), .ZN(n627) );
  INVD0 U626 ( .I(n622), .ZN(n623) );
  CKNXD16 U627 ( .I(n621), .ZN(n622) );
  CKNXD0 U628 ( .I(n624), .ZN(n625) );
  CKNXD16 U629 ( .I(n623), .ZN(n624) );
  CKNXD16 U630 ( .I(n625), .ZN(n626) );
  CKNXD0 U631 ( .I(n628), .ZN(n629) );
  CKNXD16 U632 ( .I(InParDataA[2]), .ZN(n628) );
  CKNXD0 U633 ( .I(n630), .ZN(n631) );
  INVD0 U634 ( .I(n632), .ZN(n633) );
  CKNXD16 U635 ( .I(n631), .ZN(n632) );
  CKNXD0 U636 ( .I(n634), .ZN(n635) );
  CKNXD16 U637 ( .I(n633), .ZN(n634) );
  CKNXD0 U638 ( .I(n636), .ZN(n637) );
  CKNXD16 U639 ( .I(n635), .ZN(n636) );
  CKNXD0 U640 ( .I(n638), .ZN(n639) );
  CKNXD16 U641 ( .I(n637), .ZN(n638) );
  CKNXD0 U642 ( .I(n640), .ZN(n641) );
  CKNXD16 U643 ( .I(n639), .ZN(n640) );
  CKNXD0 U644 ( .I(n642), .ZN(n643) );
  CKNXD16 U645 ( .I(n641), .ZN(n642) );
  CKNXD0 U646 ( .I(n644), .ZN(n645) );
  CKNXD16 U647 ( .I(n643), .ZN(n644) );
  CKNXD0 U648 ( .I(n646), .ZN(n647) );
  CKNXD16 U649 ( .I(n645), .ZN(n646) );
  CKNXD0 U650 ( .I(n648), .ZN(n649) );
  CKNXD16 U651 ( .I(n647), .ZN(n648) );
  CKNXD0 U652 ( .I(n762), .ZN(n763) );
  CKNXD0 U653 ( .I(n650), .ZN(n651) );
  CKNXD16 U654 ( .I(InParDataA[0]), .ZN(n650) );
  CKNXD0 U655 ( .I(n652), .ZN(n653) );
  INVD0 U656 ( .I(n654), .ZN(n655) );
  CKNXD16 U657 ( .I(n653), .ZN(n654) );
  CKNXD0 U658 ( .I(n656), .ZN(n657) );
  CKNXD16 U659 ( .I(n655), .ZN(n656) );
  CKNXD0 U660 ( .I(n658), .ZN(n659) );
  CKNXD16 U661 ( .I(n657), .ZN(n658) );
  CKNXD0 U662 ( .I(n660), .ZN(n661) );
  CKNXD16 U663 ( .I(n659), .ZN(n660) );
  CKNXD0 U664 ( .I(n662), .ZN(n663) );
  CKNXD16 U665 ( .I(n661), .ZN(n662) );
  CKNXD0 U666 ( .I(n664), .ZN(n665) );
  CKNXD16 U667 ( .I(n663), .ZN(n664) );
  CKNXD0 U668 ( .I(n666), .ZN(n667) );
  CKNXD16 U669 ( .I(n665), .ZN(n666) );
  CKNXD0 U670 ( .I(n668), .ZN(n669) );
  CKNXD16 U671 ( .I(n667), .ZN(n668) );
  CKNXD0 U672 ( .I(n670), .ZN(n671) );
  CKNXD16 U673 ( .I(n669), .ZN(n670) );
  INVD0 U674 ( .I(n672), .ZN(n673) );
  CKNXD16 U675 ( .I(n671), .ZN(n672) );
  INVD0 U676 ( .I(n674), .ZN(n675) );
  CKNXD16 U677 ( .I(InParDataB[28]), .ZN(n674) );
  CKNXD0 U678 ( .I(n676), .ZN(n677) );
  CKNXD16 U679 ( .I(n675), .ZN(n676) );
  CKNXD0 U680 ( .I(n678), .ZN(n679) );
  CKNXD16 U681 ( .I(n677), .ZN(n678) );
  CKNXD0 U682 ( .I(n680), .ZN(n681) );
  CKNXD16 U683 ( .I(n679), .ZN(n680) );
  CKNXD0 U684 ( .I(n682), .ZN(n683) );
  CKNXD16 U685 ( .I(n681), .ZN(n682) );
  CKNXD0 U686 ( .I(n684), .ZN(n685) );
  CKNXD16 U687 ( .I(n683), .ZN(n684) );
  CKNXD0 U688 ( .I(n686), .ZN(n687) );
  CKNXD16 U689 ( .I(n685), .ZN(n686) );
  CKNXD0 U690 ( .I(n692), .ZN(n693) );
  INVD0 U691 ( .I(n688), .ZN(n689) );
  CKNXD16 U692 ( .I(n687), .ZN(n688) );
  CKNXD0 U693 ( .I(n690), .ZN(n691) );
  CKNXD16 U694 ( .I(n689), .ZN(n690) );
  CKNXD16 U695 ( .I(n691), .ZN(n692) );
  INVD0 U696 ( .I(n694), .ZN(n695) );
  CKNXD16 U697 ( .I(InParDataB[27]), .ZN(n694) );
  CKNXD0 U698 ( .I(n696), .ZN(n697) );
  CKNXD16 U699 ( .I(n695), .ZN(n696) );
  CKNXD0 U700 ( .I(n698), .ZN(n699) );
  CKNXD16 U701 ( .I(n697), .ZN(n698) );
  CKNXD0 U702 ( .I(n700), .ZN(n701) );
  CKNXD16 U703 ( .I(n699), .ZN(n700) );
  CKNXD0 U704 ( .I(n702), .ZN(n703) );
  CKNXD16 U705 ( .I(n701), .ZN(n702) );
  CKNXD0 U706 ( .I(n704), .ZN(n705) );
  CKNXD16 U707 ( .I(n703), .ZN(n704) );
  CKNXD0 U708 ( .I(n706), .ZN(n707) );
  CKNXD16 U709 ( .I(n705), .ZN(n706) );
  CKNXD0 U710 ( .I(n708), .ZN(n709) );
  CKNXD16 U711 ( .I(n707), .ZN(n708) );
  CKNXD0 U712 ( .I(n710), .ZN(n711) );
  CKNXD16 U713 ( .I(n709), .ZN(n710) );
  INVD0 U714 ( .I(n712), .ZN(n713) );
  CKNXD16 U715 ( .I(n711), .ZN(n712) );
  CKNXD0 U716 ( .I(n714), .ZN(n715) );
  CKNXD16 U717 ( .I(n713), .ZN(n714) );
  INVD0 U718 ( .I(n716), .ZN(n717) );
  CKNXD16 U719 ( .I(n715), .ZN(n716) );
  CKNXD0 U720 ( .I(n732), .ZN(n733) );
  CKNXD0 U721 ( .I(n718), .ZN(n719) );
  CKNXD16 U722 ( .I(InParDataB[26]), .ZN(n718) );
  CKNXD0 U723 ( .I(n720), .ZN(n721) );
  CKNXD16 U724 ( .I(n719), .ZN(n720) );
  CKNXD0 U725 ( .I(n722), .ZN(n723) );
  CKNXD16 U726 ( .I(n721), .ZN(n722) );
  CKNXD0 U727 ( .I(n724), .ZN(n725) );
  CKNXD16 U728 ( .I(n723), .ZN(n724) );
  CKNXD0 U729 ( .I(n726), .ZN(n727) );
  CKNXD16 U730 ( .I(n725), .ZN(n726) );
  CKNXD0 U731 ( .I(n728), .ZN(n729) );
  CKNXD16 U732 ( .I(n727), .ZN(n728) );
  CKNXD0 U733 ( .I(n730), .ZN(n731) );
  CKNXD16 U734 ( .I(n729), .ZN(n730) );
  CKNXD0 U735 ( .I(n736), .ZN(n737) );
  CKNXD16 U736 ( .I(n731), .ZN(n732) );
  CKNXD0 U737 ( .I(n734), .ZN(n735) );
  CKNXD16 U738 ( .I(n733), .ZN(n734) );
  CKNXD16 U739 ( .I(n735), .ZN(n736) );
  INVD0 U740 ( .I(n738), .ZN(n739) );
  CKNXD16 U741 ( .I(InParDataB[25]), .ZN(n738) );
  CKNXD0 U742 ( .I(n740), .ZN(n741) );
  CKNXD16 U743 ( .I(n739), .ZN(n740) );
  CKNXD0 U744 ( .I(n742), .ZN(n743) );
  CKNXD16 U745 ( .I(n741), .ZN(n742) );
  CKNXD0 U746 ( .I(n744), .ZN(n745) );
  CKNXD16 U747 ( .I(n743), .ZN(n744) );
  CKNXD0 U748 ( .I(n746), .ZN(n747) );
  CKNXD16 U749 ( .I(n745), .ZN(n746) );
  CKNXD0 U750 ( .I(n748), .ZN(n749) );
  CKNXD16 U751 ( .I(n747), .ZN(n748) );
  CKNXD0 U752 ( .I(n750), .ZN(n751) );
  CKNXD16 U753 ( .I(n749), .ZN(n750) );
  CKNXD0 U754 ( .I(n752), .ZN(n753) );
  CKNXD16 U755 ( .I(n751), .ZN(n752) );
  CKNXD0 U756 ( .I(n754), .ZN(n755) );
  CKNXD16 U757 ( .I(n753), .ZN(n754) );
  INVD0 U758 ( .I(n756), .ZN(n757) );
  CKNXD16 U759 ( .I(n755), .ZN(n756) );
  CKNXD0 U760 ( .I(n758), .ZN(n759) );
  CKNXD16 U761 ( .I(n757), .ZN(n758) );
  INVD0 U762 ( .I(n760), .ZN(n761) );
  CKNXD16 U763 ( .I(n759), .ZN(n760) );
  CKNXD16 U764 ( .I(InParDataA[1]), .ZN(n762) );
  INVD0 U765 ( .I(n764), .ZN(n765) );
  CKNXD16 U766 ( .I(n649), .ZN(n764) );
  CKNXD0 U767 ( .I(n766), .ZN(n767) );
  CKNXD16 U768 ( .I(InParDataA[17]), .ZN(n766) );
  CKNXD0 U769 ( .I(n768), .ZN(n769) );
  CKNXD16 U770 ( .I(InParDataA[22]), .ZN(n768) );
  CKNXD0 U771 ( .I(n770), .ZN(n771) );
  CKNXD16 U772 ( .I(InParDataA[23]), .ZN(n770) );
  CKNXD0 U773 ( .I(n772), .ZN(n773) );
  CKNXD16 U774 ( .I(InParDataA[10]), .ZN(n772) );
  CKNXD0 U775 ( .I(n774), .ZN(n775) );
  CKNXD16 U776 ( .I(InParDataA[14]), .ZN(n774) );
  CKNXD0 U777 ( .I(n776), .ZN(n777) );
  CKNXD16 U778 ( .I(InParDataA[13]), .ZN(n776) );
  CKNXD0 U779 ( .I(n778), .ZN(n779) );
  CKNXD16 U780 ( .I(InParDataA[15]), .ZN(n778) );
  CKNXD0 U781 ( .I(n780), .ZN(n781) );
  CKNXD16 U782 ( .I(InParDataA[16]), .ZN(n780) );
  CKNXD0 U783 ( .I(n782), .ZN(n783) );
  CKNXD16 U784 ( .I(InParDataA[11]), .ZN(n782) );
  CKNXD0 U785 ( .I(n784), .ZN(n785) );
  CKNXD16 U786 ( .I(InParDataA[12]), .ZN(n784) );
  CKNXD0 U787 ( .I(n786), .ZN(n787) );
  CKNXD16 U788 ( .I(InParDataA[3]), .ZN(n786) );
  CKNXD0 U789 ( .I(n788), .ZN(n789) );
  CKNXD16 U790 ( .I(InParDataA[7]), .ZN(n788) );
  CKNXD0 U791 ( .I(n790), .ZN(n791) );
  CKNXD16 U792 ( .I(InParDataA[8]), .ZN(n790) );
  CKNXD0 U793 ( .I(n792), .ZN(n793) );
  CKNXD16 U794 ( .I(InParDataA[9]), .ZN(n792) );
  CKNXD0 U795 ( .I(n794), .ZN(n795) );
  CKNXD16 U796 ( .I(InParDataA[6]), .ZN(n794) );
  CKNXD0 U797 ( .I(n796), .ZN(n797) );
  CKNXD16 U798 ( .I(InParDataA[4]), .ZN(n796) );
  CKNXD0 U799 ( .I(n798), .ZN(n799) );
  CKNXD16 U800 ( .I(InParDataA[5]), .ZN(n798) );
  CKNXD0 U801 ( .I(n800), .ZN(n801) );
  CKNXD16 U802 ( .I(n673), .ZN(n800) );
  CKNXD0 U803 ( .I(n802), .ZN(n803) );
  CKNXD16 U804 ( .I(n763), .ZN(n802) );
  CKNXD0 U805 ( .I(n804), .ZN(n805) );
  CKNXD16 U806 ( .I(n765), .ZN(n804) );
  CKNXD0 U807 ( .I(n806), .ZN(n807) );
  CKNXD16 U808 ( .I(InParDataA[31]), .ZN(n806) );
  CKNXD0 U809 ( .I(n808), .ZN(n809) );
  CKNXD16 U810 ( .I(n807), .ZN(n808) );
  CKNXD0 U811 ( .I(n810), .ZN(n811) );
  CKNXD16 U812 ( .I(n809), .ZN(n810) );
  CKNXD0 U813 ( .I(n812), .ZN(n813) );
  CKNXD16 U814 ( .I(n811), .ZN(n812) );
  CKNXD0 U815 ( .I(n814), .ZN(n815) );
  CKNXD16 U816 ( .I(n813), .ZN(n814) );
  CKNXD0 U817 ( .I(n816), .ZN(n817) );
  CKNXD16 U818 ( .I(n815), .ZN(n816) );
  CKNXD0 U819 ( .I(n818), .ZN(n819) );
  CKNXD16 U820 ( .I(n817), .ZN(n818) );
  CKNXD0 U821 ( .I(n820), .ZN(n821) );
  CKNXD16 U822 ( .I(n819), .ZN(n820) );
  INVD0 U823 ( .I(n822), .ZN(n823) );
  CKNXD16 U824 ( .I(n821), .ZN(n822) );
  CKNXD0 U825 ( .I(n824), .ZN(n825) );
  CKNXD16 U826 ( .I(n823), .ZN(n824) );
  CKNXD12 U827 ( .I(n829), .ZN(n830) );
  CKNXD0 U828 ( .I(n826), .ZN(n827) );
  CKNXD16 U829 ( .I(InParDataA[30]), .ZN(n826) );
  CKNXD0 U830 ( .I(n828), .ZN(n829) );
  CKNXD16 U831 ( .I(n827), .ZN(n828) );
  CKNXD0 U832 ( .I(n830), .ZN(n831) );
  CKNXD0 U833 ( .I(n832), .ZN(n833) );
  CKNXD16 U834 ( .I(n831), .ZN(n832) );
  CKNXD0 U835 ( .I(n834), .ZN(n835) );
  CKNXD16 U836 ( .I(n833), .ZN(n834) );
  CKNXD0 U837 ( .I(n836), .ZN(n837) );
  CKNXD16 U838 ( .I(n835), .ZN(n836) );
  CKNXD0 U839 ( .I(n838), .ZN(n839) );
  CKNXD16 U840 ( .I(n837), .ZN(n838) );
  CKNXD0 U841 ( .I(n840), .ZN(n841) );
  CKNXD16 U842 ( .I(n839), .ZN(n840) );
  INVD0 U843 ( .I(n842), .ZN(n843) );
  CKNXD16 U844 ( .I(n841), .ZN(n842) );
  CKNXD0 U845 ( .I(n844), .ZN(n845) );
  CKNXD16 U846 ( .I(n843), .ZN(n844) );
  CKNXD0 U847 ( .I(n846), .ZN(n847) );
  CKNXD16 U848 ( .I(InParDataA[29]), .ZN(n846) );
  CKNXD0 U849 ( .I(n848), .ZN(n849) );
  CKNXD16 U850 ( .I(n847), .ZN(n848) );
  CKNXD0 U851 ( .I(n850), .ZN(n851) );
  CKNXD16 U852 ( .I(n849), .ZN(n850) );
  CKNXD0 U853 ( .I(n852), .ZN(n853) );
  CKNXD16 U854 ( .I(n851), .ZN(n852) );
  CKNXD0 U855 ( .I(n854), .ZN(n855) );
  CKNXD16 U856 ( .I(n853), .ZN(n854) );
  CKNXD0 U857 ( .I(n856), .ZN(n857) );
  CKNXD16 U858 ( .I(n855), .ZN(n856) );
  CKNXD0 U859 ( .I(n858), .ZN(n859) );
  CKNXD16 U860 ( .I(n857), .ZN(n858) );
  CKNXD0 U861 ( .I(n860), .ZN(n861) );
  CKNXD16 U862 ( .I(n859), .ZN(n860) );
  INVD0 U863 ( .I(n862), .ZN(n863) );
  CKNXD16 U864 ( .I(n861), .ZN(n862) );
  CKNXD0 U865 ( .I(n864), .ZN(n865) );
  CKNXD16 U866 ( .I(n863), .ZN(n864) );
  CKNXD0 U867 ( .I(n866), .ZN(n867) );
  CKNXD16 U868 ( .I(InParDataA[28]), .ZN(n866) );
  CKNXD0 U869 ( .I(n868), .ZN(n869) );
  CKNXD16 U870 ( .I(n867), .ZN(n868) );
  CKNXD0 U871 ( .I(n870), .ZN(n871) );
  CKNXD16 U872 ( .I(n869), .ZN(n870) );
  CKNXD0 U873 ( .I(n872), .ZN(n873) );
  CKNXD16 U874 ( .I(n871), .ZN(n872) );
  CKNXD0 U875 ( .I(n874), .ZN(n875) );
  CKNXD16 U876 ( .I(n873), .ZN(n874) );
  CKNXD0 U877 ( .I(n876), .ZN(n877) );
  CKNXD16 U878 ( .I(n875), .ZN(n876) );
  CKNXD0 U879 ( .I(n878), .ZN(n879) );
  CKNXD16 U880 ( .I(n877), .ZN(n878) );
  CKNXD0 U881 ( .I(n880), .ZN(n881) );
  CKNXD16 U882 ( .I(n879), .ZN(n880) );
  INVD0 U883 ( .I(n882), .ZN(n883) );
  CKNXD16 U884 ( .I(n881), .ZN(n882) );
  CKNXD0 U885 ( .I(n884), .ZN(n885) );
  CKNXD16 U886 ( .I(n883), .ZN(n884) );
  CKNXD0 U887 ( .I(n886), .ZN(n887) );
  CKNXD16 U888 ( .I(InParDataA[27]), .ZN(n886) );
  CKNXD0 U889 ( .I(n888), .ZN(n889) );
  CKNXD16 U890 ( .I(n887), .ZN(n888) );
  CKNXD0 U891 ( .I(n890), .ZN(n891) );
  CKNXD16 U892 ( .I(n889), .ZN(n890) );
  CKNXD0 U893 ( .I(n892), .ZN(n893) );
  CKNXD16 U894 ( .I(n891), .ZN(n892) );
  CKNXD0 U895 ( .I(n894), .ZN(n895) );
  CKNXD16 U896 ( .I(n893), .ZN(n894) );
  CKNXD0 U897 ( .I(n896), .ZN(n897) );
  CKNXD16 U898 ( .I(n895), .ZN(n896) );
  CKNXD0 U899 ( .I(n898), .ZN(n899) );
  CKNXD16 U900 ( .I(n897), .ZN(n898) );
  CKNXD0 U901 ( .I(n900), .ZN(n901) );
  CKNXD16 U902 ( .I(n899), .ZN(n900) );
  INVD0 U903 ( .I(n902), .ZN(n903) );
  CKNXD16 U904 ( .I(n901), .ZN(n902) );
  CKNXD0 U905 ( .I(n904), .ZN(n905) );
  CKNXD16 U906 ( .I(n903), .ZN(n904) );
  CKNXD0 U907 ( .I(n906), .ZN(n907) );
  CKNXD16 U908 ( .I(InParDataA[26]), .ZN(n906) );
  CKNXD0 U909 ( .I(n908), .ZN(n909) );
  CKNXD16 U910 ( .I(n907), .ZN(n908) );
  CKNXD0 U911 ( .I(n910), .ZN(n911) );
  CKNXD16 U912 ( .I(n909), .ZN(n910) );
  CKNXD0 U913 ( .I(n912), .ZN(n913) );
  CKNXD16 U914 ( .I(n911), .ZN(n912) );
  CKNXD0 U915 ( .I(n914), .ZN(n915) );
  CKNXD16 U916 ( .I(n913), .ZN(n914) );
  CKNXD0 U917 ( .I(n916), .ZN(n917) );
  CKNXD16 U918 ( .I(n915), .ZN(n916) );
  CKNXD0 U919 ( .I(n918), .ZN(n919) );
  CKNXD16 U920 ( .I(n917), .ZN(n918) );
  CKNXD0 U921 ( .I(n920), .ZN(n921) );
  CKNXD16 U922 ( .I(n919), .ZN(n920) );
  INVD0 U923 ( .I(n922), .ZN(n923) );
  CKNXD16 U924 ( .I(n921), .ZN(n922) );
  CKNXD0 U925 ( .I(n924), .ZN(n925) );
  CKNXD16 U926 ( .I(n923), .ZN(n924) );
  CKNXD0 U927 ( .I(n926), .ZN(n927) );
  CKNXD16 U928 ( .I(InParDataA[25]), .ZN(n926) );
  CKNXD0 U929 ( .I(n928), .ZN(n929) );
  CKNXD16 U930 ( .I(n927), .ZN(n928) );
  CKNXD0 U931 ( .I(n930), .ZN(n931) );
  CKNXD16 U932 ( .I(n929), .ZN(n930) );
  CKNXD0 U933 ( .I(n932), .ZN(n933) );
  CKNXD16 U934 ( .I(n931), .ZN(n932) );
  CKNXD0 U935 ( .I(n934), .ZN(n935) );
  CKNXD16 U936 ( .I(n933), .ZN(n934) );
  CKNXD0 U937 ( .I(n936), .ZN(n937) );
  CKNXD16 U938 ( .I(n935), .ZN(n936) );
  CKNXD0 U939 ( .I(n938), .ZN(n939) );
  CKNXD16 U940 ( .I(n937), .ZN(n938) );
  CKNXD0 U941 ( .I(n940), .ZN(n941) );
  CKNXD16 U942 ( .I(n939), .ZN(n940) );
  INVD0 U943 ( .I(n942), .ZN(n943) );
  CKNXD16 U944 ( .I(n941), .ZN(n942) );
  CKNXD0 U945 ( .I(n944), .ZN(n945) );
  CKNXD16 U946 ( .I(n943), .ZN(n944) );
  CKNXD0 U947 ( .I(n946), .ZN(n947) );
  CKNXD16 U948 ( .I(InParDataA[24]), .ZN(n946) );
  CKNXD0 U949 ( .I(n948), .ZN(n949) );
  CKNXD16 U950 ( .I(n947), .ZN(n948) );
  CKNXD0 U951 ( .I(n950), .ZN(n951) );
  CKNXD16 U952 ( .I(n949), .ZN(n950) );
  CKNXD0 U953 ( .I(n952), .ZN(n953) );
  CKNXD16 U954 ( .I(n951), .ZN(n952) );
  CKNXD0 U955 ( .I(n954), .ZN(n955) );
  CKNXD16 U956 ( .I(n953), .ZN(n954) );
  CKNXD0 U957 ( .I(n956), .ZN(n957) );
  CKNXD16 U958 ( .I(n955), .ZN(n956) );
  CKNXD0 U959 ( .I(n958), .ZN(n959) );
  CKNXD16 U960 ( .I(n957), .ZN(n958) );
  CKNXD0 U961 ( .I(n960), .ZN(n961) );
  CKNXD16 U962 ( .I(n959), .ZN(n960) );
  CKNXD0 U963 ( .I(n962), .ZN(n963) );
  CKNXD16 U964 ( .I(n961), .ZN(n962) );
  INVD0 U965 ( .I(n964), .ZN(n965) );
  CKNXD16 U966 ( .I(n963), .ZN(n964) );
  CKNXD0 U967 ( .I(n966), .ZN(n967) );
  CKNXD16 U968 ( .I(n965), .ZN(n966) );
  INVD0 U969 ( .I(n968), .ZN(n969) );
  CKNXD16 U970 ( .I(InParDataA[21]), .ZN(n968) );
  CKNXD0 U971 ( .I(n970), .ZN(n971) );
  CKNXD16 U972 ( .I(n969), .ZN(n970) );
  CKNXD0 U973 ( .I(n972), .ZN(n973) );
  CKNXD16 U974 ( .I(n971), .ZN(n972) );
  CKNXD0 U975 ( .I(n974), .ZN(n975) );
  CKNXD16 U976 ( .I(n973), .ZN(n974) );
  CKNXD0 U977 ( .I(n976), .ZN(n977) );
  CKNXD16 U978 ( .I(n975), .ZN(n976) );
  CKNXD0 U979 ( .I(n978), .ZN(n979) );
  CKNXD16 U980 ( .I(n977), .ZN(n978) );
  CKNXD0 U981 ( .I(n980), .ZN(n981) );
  CKNXD16 U982 ( .I(n979), .ZN(n980) );
  CKNXD0 U983 ( .I(n982), .ZN(n983) );
  CKNXD16 U984 ( .I(n981), .ZN(n982) );
  CKNXD0 U985 ( .I(n984), .ZN(n985) );
  CKNXD16 U986 ( .I(n983), .ZN(n984) );
  INVD0 U987 ( .I(n986), .ZN(n987) );
  CKNXD16 U988 ( .I(n985), .ZN(n986) );
  CKNXD0 U989 ( .I(n988), .ZN(n989) );
  CKNXD16 U990 ( .I(n987), .ZN(n988) );
  INVD0 U991 ( .I(n990), .ZN(n991) );
  CKNXD16 U992 ( .I(InParDataA[20]), .ZN(n990) );
  CKNXD0 U993 ( .I(n992), .ZN(n993) );
  CKNXD16 U994 ( .I(n991), .ZN(n992) );
  CKNXD0 U995 ( .I(n994), .ZN(n995) );
  CKNXD16 U996 ( .I(n993), .ZN(n994) );
  CKNXD0 U997 ( .I(n996), .ZN(n997) );
  CKNXD16 U998 ( .I(n995), .ZN(n996) );
  CKNXD0 U999 ( .I(n998), .ZN(n999) );
  CKNXD16 U1000 ( .I(n997), .ZN(n998) );
  CKNXD0 U1001 ( .I(n1000), .ZN(n1001) );
  CKNXD16 U1002 ( .I(n999), .ZN(n1000) );
  CKNXD0 U1003 ( .I(n1002), .ZN(n1003) );
  CKNXD16 U1004 ( .I(n1001), .ZN(n1002) );
  CKNXD0 U1005 ( .I(n1004), .ZN(n1005) );
  CKNXD16 U1006 ( .I(n1003), .ZN(n1004) );
  CKNXD0 U1007 ( .I(n1006), .ZN(n1007) );
  CKNXD16 U1008 ( .I(n1005), .ZN(n1006) );
  INVD0 U1009 ( .I(n1008), .ZN(n1009) );
  CKNXD16 U1010 ( .I(n1007), .ZN(n1008) );
  CKNXD0 U1011 ( .I(n1010), .ZN(n1011) );
  CKNXD16 U1012 ( .I(n1009), .ZN(n1010) );
  CKNXD0 U1013 ( .I(n1012), .ZN(n1013) );
  CKNXD16 U1014 ( .I(InParDataA[19]), .ZN(n1012) );
  CKNXD0 U1015 ( .I(n1014), .ZN(n1015) );
  CKNXD16 U1016 ( .I(n1013), .ZN(n1014) );
  CKNXD0 U1017 ( .I(n1016), .ZN(n1017) );
  CKNXD16 U1018 ( .I(n1015), .ZN(n1016) );
  CKNXD0 U1019 ( .I(n1018), .ZN(n1019) );
  CKNXD16 U1020 ( .I(n1017), .ZN(n1018) );
  CKNXD0 U1021 ( .I(n1020), .ZN(n1021) );
  CKNXD16 U1022 ( .I(n1019), .ZN(n1020) );
  CKNXD0 U1023 ( .I(n1022), .ZN(n1023) );
  CKNXD16 U1024 ( .I(n1021), .ZN(n1022) );
  CKNXD0 U1025 ( .I(n1024), .ZN(n1025) );
  CKNXD16 U1026 ( .I(n1023), .ZN(n1024) );
  CKNXD0 U1027 ( .I(n1026), .ZN(n1027) );
  CKNXD16 U1028 ( .I(n1025), .ZN(n1026) );
  CKNXD0 U1029 ( .I(n1028), .ZN(n1029) );
  CKNXD16 U1030 ( .I(n1027), .ZN(n1028) );
  INVD0 U1031 ( .I(n1030), .ZN(n1031) );
  CKNXD16 U1032 ( .I(n1029), .ZN(n1030) );
  CKNXD0 U1033 ( .I(n1032), .ZN(n1033) );
  CKNXD16 U1034 ( .I(n1031), .ZN(n1032) );
  INVD0 U1035 ( .I(n1034), .ZN(n1035) );
  CKNXD16 U1036 ( .I(InParDataA[18]), .ZN(n1034) );
  CKNXD0 U1037 ( .I(n1036), .ZN(n1037) );
  CKNXD16 U1038 ( .I(n1035), .ZN(n1036) );
  CKNXD0 U1039 ( .I(n1038), .ZN(n1039) );
  CKNXD16 U1040 ( .I(n1037), .ZN(n1038) );
  CKNXD0 U1041 ( .I(n1040), .ZN(n1041) );
  CKNXD16 U1042 ( .I(n1039), .ZN(n1040) );
  CKNXD0 U1043 ( .I(n1042), .ZN(n1043) );
  CKNXD16 U1044 ( .I(n1041), .ZN(n1042) );
  CKNXD0 U1045 ( .I(n1044), .ZN(n1045) );
  CKNXD16 U1046 ( .I(n1043), .ZN(n1044) );
  CKNXD0 U1047 ( .I(n1046), .ZN(n1047) );
  CKNXD16 U1048 ( .I(n1045), .ZN(n1046) );
  CKNXD0 U1049 ( .I(n1048), .ZN(n1049) );
  CKNXD16 U1050 ( .I(n1047), .ZN(n1048) );
  CKNXD0 U1051 ( .I(n1050), .ZN(n1051) );
  CKNXD16 U1052 ( .I(n1049), .ZN(n1050) );
  INVD0 U1053 ( .I(n1052), .ZN(n1053) );
  CKNXD16 U1054 ( .I(n1051), .ZN(n1052) );
  CKNXD0 U1055 ( .I(n1054), .ZN(n1055) );
  CKNXD16 U1056 ( .I(n1053), .ZN(n1054) );
  CKNXD0 U1057 ( .I(n1056), .ZN(n1057) );
  CKNXD16 U1058 ( .I(InParValidB), .ZN(n1056) );
  CKNXD0 U1059 ( .I(n1058), .ZN(n1059) );
  CKNXD16 U1060 ( .I(InParValidA), .ZN(n1058) );
  BUFFD1 U1061 ( .I(ClockB), .Z(n1060) );
  BUFFD1 U1062 ( .I(ClockA), .Z(n1061) );
  TIEH U1063 ( .Z(\*Logic1* ) );
endmodule


module SerDes_DWid32_RxLogDepth4_TxLogDepth3 ( ParOutRxClk, SerLineXfer, 
        ParDataIn, InParClk, InParValid, OutParClk, RxRequest, TxRequest, 
        Reset );
  output [31:0] ParOutRxClk;
  input [31:0] ParDataIn;
  input InParClk, InParValid, OutParClk, RxRequest, TxRequest, Reset;
  output SerLineXfer;
  wire   SerLineValid, Tx_F_Empty, Tx_F_Full, Rx_F_Empty, Rx_F_Full, n1, n2,
         n3, n4;

  Serializer_DWid32_AWid3 Ser_U1 ( .SerOut(SerLineXfer), .SerValid(
        SerLineValid), .FIFOEmpty(Tx_F_Empty), .FIFOFull(Tx_F_Full), .ParIn(
        ParDataIn), .InParValid(InParValid), .ParInClk(n4), .SendSerial(
        TxRequest), .Reset(n1) );
  Deserializer_AWid4_DWid32 Des_U1 ( .ParOut(ParOutRxClk), .FIFOEmpty(
        Rx_F_Empty), .FIFOFull(Rx_F_Full), .ParOutClk(n3), .SerialIn(
        SerLineXfer), .ReadReq(RxRequest), .SerValid(SerLineValid), .Reset(n1)
         );
  BUFFD2 U1 ( .I(OutParClk), .Z(n3) );
  INVD1 U2 ( .I(n2), .ZN(n1) );
  INVD1 U3 ( .I(Reset), .ZN(n2) );
  BUFFD1 U4 ( .I(InParClk), .Z(n4) );
endmodule


module SerDes_DWid32_RxLogDepth3_TxLogDepth4 ( ParOutRxClk, SerLineXfer, 
        ParDataIn, InParClk, InParValid, OutParClk, RxRequest, TxRequest, 
        Reset );
  output [31:0] ParOutRxClk;
  input [31:0] ParDataIn;
  input InParClk, InParValid, OutParClk, RxRequest, TxRequest, Reset;
  output SerLineXfer;
  wire   SerLineValid, Tx_F_Empty, Tx_F_Full, Rx_F_Empty, Rx_F_Full, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  Serializer_DWid32_AWid4 Ser_U1 ( .SerOut(SerLineXfer), .SerValid(
        SerLineValid), .FIFOEmpty(Tx_F_Empty), .FIFOFull(Tx_F_Full), .ParIn(
        ParDataIn), .InParValid(InParValid), .ParInClk(n15), .SendSerial(
        TxRequest), .Reset(n1) );
  Deserializer_AWid3_DWid32 Des_U1 ( .ParOut(ParOutRxClk), .FIFOEmpty(
        Rx_F_Empty), .FIFOFull(Rx_F_Full), .ParOutClk(n16), .SerialIn(
        SerLineXfer), .ReadReq(RxRequest), .SerValid(SerLineValid), .Reset(n1)
         );
  BUFFD0 U1 ( .I(n2), .Z(n1) );
  BUFFD0 U2 ( .I(n3), .Z(n2) );
  BUFFD0 U3 ( .I(n4), .Z(n3) );
  BUFFD0 U4 ( .I(n5), .Z(n4) );
  BUFFD0 U5 ( .I(n6), .Z(n5) );
  BUFFD0 U6 ( .I(n7), .Z(n6) );
  BUFFD0 U7 ( .I(n8), .Z(n7) );
  BUFFD0 U8 ( .I(n9), .Z(n8) );
  BUFFD0 U9 ( .I(n10), .Z(n9) );
  BUFFD0 U10 ( .I(n11), .Z(n10) );
  BUFFD0 U11 ( .I(n12), .Z(n11) );
  BUFFD0 U12 ( .I(n13), .Z(n12) );
  BUFFD2 U13 ( .I(OutParClk), .Z(n16) );
  INVD1 U14 ( .I(n14), .ZN(n13) );
  INVD1 U15 ( .I(Reset), .ZN(n14) );
  BUFFD1 U16 ( .I(InParClk), .Z(n15) );
endmodule


module Serializer_DWid32_AWid3 ( SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk, 
        ParIn, InParValid, ParInClk, SendSerial, Reset );
  input [31:0] ParIn;
  input InParValid, ParInClk, SendSerial, Reset;
  output SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk;
  wire   F_Valid, SerEncReadReq, F_ReadReq, F_WriteReq, EncD_ToTx, n2, n1, n3,
         n4;
  wire   [31:0] FIFO_Out;

  FIFOTop_AWid3_DWid32_0 FIFO_Tx1 ( .Dout(FIFO_Out), .Din(ParIn), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(n1), .WriteIn(F_WriteReq), 
        .ClkR(ParInClk), .ClkW(ParInClk), .Reseter(n3) );
  SerEncoder_DWid32_0 SerEnc_Tx1 ( .SerOut(EncD_ToTx), .SerValid(SerValid), 
        .FIFO_ReadReq(SerEncReadReq), .ParIn(FIFO_Out), .F_Empty(FIFOEmpty), 
        .ParClk(ParInClk), .SerClk(SerClk), .ParValid(F_Valid), .Reset(n3) );
  SerialTx_0 SerTx_Tx1 ( .SerOut(SerOut), .SerClk(SerClk), .SerIn(EncD_ToTx), 
        .ParClk(ParInClk), .Reset(n3) );
  INR2XD0 U1 ( .A1(InParValid), .B1(FIFOFull), .ZN(F_WriteReq) );
  BUFFD0 U2 ( .I(F_ReadReq), .Z(n1) );
  INVD1 U3 ( .I(n4), .ZN(n3) );
  INVD1 U4 ( .I(Reset), .ZN(n4) );
  AN3D1 U5 ( .A1(n2), .A2(SendSerial), .A3(SerEncReadReq), .Z(F_ReadReq) );
  INVD1 U6 ( .I(FIFOEmpty), .ZN(n2) );
  NR2D1 U7 ( .A1(n3), .A2(FIFOEmpty), .ZN(F_Valid) );
endmodule


module Deserializer_AWid4_DWid32 ( ParOut, ParValid, DecoderParClk, FIFOEmpty, 
        FIFOFull, ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, N3, N4,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, ParValidDecode, SerialClk, SerRxToDecode, n3, n1, n2, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n61, n63,
         n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91,
         n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, n113, n115,
         n117, n119, n121, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid4_DWid32_0 FIFO_Rx1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), 
        .Full(FIFOFull), .Empty(FIFOEmpty), .ReadIn(ReadReq), .WriteIn(
        ParValidDecode), .ClkR(ParOutClk), .ClkW(DecoderParClk), .Reseter(n155) );
  DesDecoder_DWid32_0 DesDec_Rx1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(n155) );
  SerialRx_0 SerRx_Rx1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(n155) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(n1), .CP(ParOutClk), .CDN(n157), .Q(n158) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(n2), .CP(ParOutClk), .CDN(n157), .Q(n159) );
  DFCNQD1 \ParBuf_reg[29]  ( .D(n4), .CP(ParOutClk), .CDN(n157), .Q(n160) );
  DFCNQD1 \ParBuf_reg[28]  ( .D(n5), .CP(ParOutClk), .CDN(n157), .Q(n161) );
  DFCNQD1 \ParBuf_reg[27]  ( .D(n6), .CP(ParOutClk), .CDN(n157), .Q(n162) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(n7), .CP(ParOutClk), .CDN(n157), .Q(n163) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(n8), .CP(ParOutClk), .CDN(n156), .Q(n164) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(n9), .CP(ParOutClk), .CDN(n157), .Q(n165) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(n10), .CP(ParOutClk), .CDN(n157), .Q(n166) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(n11), .CP(ParOutClk), .CDN(n157), .Q(n167) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(n12), .CP(ParOutClk), .CDN(n157), .Q(n168) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(n13), .CP(ParOutClk), .CDN(n157), .Q(n169) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(n14), .CP(ParOutClk), .CDN(n157), .Q(n170) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(n15), .CP(ParOutClk), .CDN(n157), .Q(n171) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(n16), .CP(ParOutClk), .CDN(n156), .Q(n172) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(n17), .CP(ParOutClk), .CDN(n156), .Q(n173) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(n18), .CP(ParOutClk), .CDN(n156), .Q(n174) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(n19), .CP(ParOutClk), .CDN(n156), .Q(n175) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(n20), .CP(ParOutClk), .CDN(n156), .Q(n176) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(n21), .CP(ParOutClk), .CDN(n156), .Q(n177) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(n22), .CP(ParOutClk), .CDN(n156), .Q(n178) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(n23), .CP(ParOutClk), .CDN(n157), .Q(n179) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(n24), .CP(ParOutClk), .CDN(n157), .Q(n180) );
  DFCNQD1 \ParBuf_reg[8]  ( .D(n25), .CP(ParOutClk), .CDN(n157), .Q(n181) );
  DFCNQD1 \ParBuf_reg[7]  ( .D(n26), .CP(ParOutClk), .CDN(n157), .Q(n182) );
  DFCNQD1 \ParBuf_reg[6]  ( .D(n27), .CP(ParOutClk), .CDN(n157), .Q(n183) );
  DFCNQD1 \ParBuf_reg[5]  ( .D(n28), .CP(ParOutClk), .CDN(n157), .Q(n184) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(n29), .CP(ParOutClk), .CDN(n156), .Q(n185) );
  DFCNQD1 \ParBuf_reg[3]  ( .D(n30), .CP(ParOutClk), .CDN(n156), .Q(n186) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(n31), .CP(ParOutClk), .CDN(n156), .Q(n187) );
  DFCNQD1 \ParBuf_reg[1]  ( .D(n32), .CP(ParOutClk), .CDN(n156), .Q(n188) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(n33), .CP(ParOutClk), .CDN(n156), .Q(n189) );
  DFCNQD1 ParValidr_reg ( .D(n34), .CP(ParOutClk), .CDN(n156), .Q(ParValid) );
  CKBD0 U3 ( .CLK(N34), .C(n1) );
  CKBD0 U4 ( .CLK(N33), .C(n2) );
  CKBD0 U5 ( .CLK(N32), .C(n4) );
  CKBD0 U6 ( .CLK(N31), .C(n5) );
  CKBD0 U7 ( .CLK(N30), .C(n6) );
  CKBD0 U8 ( .CLK(N29), .C(n7) );
  CKBD0 U9 ( .CLK(N28), .C(n8) );
  CKBD0 U10 ( .CLK(N27), .C(n9) );
  CKBD0 U11 ( .CLK(N26), .C(n10) );
  CKBD0 U12 ( .CLK(N25), .C(n11) );
  CKBD0 U13 ( .CLK(N24), .C(n12) );
  CKBD0 U14 ( .CLK(N23), .C(n13) );
  CKBD0 U15 ( .CLK(N22), .C(n14) );
  CKBD0 U16 ( .CLK(N21), .C(n15) );
  CKBD0 U17 ( .CLK(N20), .C(n16) );
  CKBD0 U18 ( .CLK(N19), .C(n17) );
  CKBD0 U19 ( .CLK(N18), .C(n18) );
  CKBD0 U20 ( .CLK(N17), .C(n19) );
  CKBD0 U21 ( .CLK(N16), .C(n20) );
  CKBD0 U22 ( .CLK(N15), .C(n21) );
  CKBD0 U23 ( .CLK(N14), .C(n22) );
  CKBD0 U24 ( .CLK(N13), .C(n23) );
  CKBD0 U25 ( .CLK(N12), .C(n24) );
  CKBD0 U26 ( .CLK(N11), .C(n25) );
  CKBD0 U27 ( .CLK(N10), .C(n26) );
  CKBD0 U28 ( .CLK(N9), .C(n27) );
  CKBD0 U29 ( .CLK(N8), .C(n28) );
  BUFFD0 U30 ( .I(N7), .Z(n29) );
  BUFFD0 U31 ( .I(N6), .Z(n30) );
  BUFFD0 U32 ( .I(N5), .Z(n31) );
  BUFFD0 U33 ( .I(N4), .Z(n32) );
  BUFFD0 U34 ( .I(N3), .Z(n33) );
  BUFFD0 U35 ( .I(n35), .Z(n34) );
  BUFFD0 U36 ( .I(n36), .Z(n35) );
  BUFFD0 U37 ( .I(n37), .Z(n36) );
  BUFFD0 U38 ( .I(n38), .Z(n37) );
  BUFFD0 U39 ( .I(n39), .Z(n38) );
  BUFFD0 U40 ( .I(n40), .Z(n39) );
  BUFFD0 U41 ( .I(n41), .Z(n40) );
  BUFFD0 U42 ( .I(n42), .Z(n41) );
  BUFFD0 U43 ( .I(n43), .Z(n42) );
  BUFFD0 U44 ( .I(n44), .Z(n43) );
  BUFFD0 U45 ( .I(n45), .Z(n44) );
  BUFFD0 U46 ( .I(n46), .Z(n45) );
  BUFFD0 U47 ( .I(n47), .Z(n46) );
  BUFFD0 U48 ( .I(n48), .Z(n47) );
  BUFFD0 U49 ( .I(n49), .Z(n48) );
  BUFFD0 U50 ( .I(n50), .Z(n49) );
  BUFFD0 U51 ( .I(n51), .Z(n50) );
  BUFFD0 U52 ( .I(n52), .Z(n51) );
  BUFFD0 U53 ( .I(n53), .Z(n52) );
  BUFFD0 U54 ( .I(n54), .Z(n53) );
  BUFFD0 U55 ( .I(n55), .Z(n54) );
  BUFFD0 U56 ( .I(n56), .Z(n55) );
  BUFFD0 U57 ( .I(n57), .Z(n56) );
  BUFFD0 U58 ( .I(n58), .Z(n57) );
  BUFFD0 U59 ( .I(N35), .Z(n58) );
  CKBD0 U60 ( .CLK(n154), .C(n59) );
  CKNXD16 U61 ( .I(n59), .ZN(ParOut[31]) );
  CKBD0 U62 ( .CLK(n153), .C(n61) );
  CKNXD16 U63 ( .I(n61), .ZN(ParOut[30]) );
  CKBD0 U64 ( .CLK(n152), .C(n63) );
  CKNXD16 U65 ( .I(n63), .ZN(ParOut[29]) );
  CKBD0 U66 ( .CLK(n151), .C(n65) );
  CKNXD16 U67 ( .I(n65), .ZN(ParOut[28]) );
  CKBD0 U68 ( .CLK(n150), .C(n67) );
  CKNXD16 U69 ( .I(n67), .ZN(ParOut[27]) );
  CKBD0 U70 ( .CLK(n149), .C(n69) );
  CKNXD16 U71 ( .I(n69), .ZN(ParOut[26]) );
  CKBD0 U72 ( .CLK(n148), .C(n71) );
  CKNXD16 U73 ( .I(n71), .ZN(ParOut[25]) );
  CKBD0 U74 ( .CLK(n147), .C(n73) );
  CKNXD16 U75 ( .I(n73), .ZN(ParOut[24]) );
  CKBD0 U76 ( .CLK(n146), .C(n75) );
  CKNXD16 U77 ( .I(n75), .ZN(ParOut[23]) );
  CKBD0 U78 ( .CLK(n145), .C(n77) );
  CKNXD16 U79 ( .I(n77), .ZN(ParOut[22]) );
  CKBD0 U80 ( .CLK(n144), .C(n79) );
  CKNXD16 U81 ( .I(n79), .ZN(ParOut[21]) );
  CKBD0 U82 ( .CLK(n143), .C(n81) );
  CKNXD16 U83 ( .I(n81), .ZN(ParOut[20]) );
  CKBD0 U84 ( .CLK(n142), .C(n83) );
  CKNXD16 U85 ( .I(n83), .ZN(ParOut[19]) );
  CKBD0 U86 ( .CLK(n141), .C(n85) );
  CKNXD16 U87 ( .I(n85), .ZN(ParOut[18]) );
  CKBD0 U88 ( .CLK(n140), .C(n87) );
  CKNXD16 U89 ( .I(n87), .ZN(ParOut[17]) );
  CKBD0 U90 ( .CLK(n139), .C(n89) );
  CKNXD16 U91 ( .I(n89), .ZN(ParOut[16]) );
  CKBD0 U92 ( .CLK(n138), .C(n91) );
  CKNXD16 U93 ( .I(n91), .ZN(ParOut[15]) );
  CKBD0 U94 ( .CLK(n137), .C(n93) );
  CKNXD16 U95 ( .I(n93), .ZN(ParOut[14]) );
  CKBD0 U96 ( .CLK(n136), .C(n95) );
  CKNXD16 U97 ( .I(n95), .ZN(ParOut[13]) );
  CKBD0 U98 ( .CLK(n135), .C(n97) );
  CKNXD16 U99 ( .I(n97), .ZN(ParOut[12]) );
  CKBD0 U100 ( .CLK(n134), .C(n99) );
  CKNXD16 U101 ( .I(n99), .ZN(ParOut[11]) );
  CKBD0 U102 ( .CLK(n133), .C(n101) );
  CKNXD16 U103 ( .I(n101), .ZN(ParOut[10]) );
  CKBD0 U104 ( .CLK(n132), .C(n103) );
  CKNXD16 U105 ( .I(n103), .ZN(ParOut[9]) );
  CKBD0 U106 ( .CLK(n131), .C(n105) );
  CKNXD16 U107 ( .I(n105), .ZN(ParOut[8]) );
  CKBD0 U108 ( .CLK(n130), .C(n107) );
  CKNXD16 U109 ( .I(n107), .ZN(ParOut[7]) );
  CKBD0 U110 ( .CLK(n129), .C(n109) );
  CKNXD16 U111 ( .I(n109), .ZN(ParOut[6]) );
  CKBD0 U112 ( .CLK(n128), .C(n111) );
  CKNXD16 U113 ( .I(n111), .ZN(ParOut[5]) );
  CKBD0 U114 ( .CLK(n127), .C(n113) );
  CKNXD16 U115 ( .I(n113), .ZN(ParOut[4]) );
  CKBD0 U116 ( .CLK(n126), .C(n115) );
  CKNXD16 U117 ( .I(n115), .ZN(ParOut[3]) );
  CKBD0 U118 ( .CLK(n125), .C(n117) );
  CKNXD16 U119 ( .I(n117), .ZN(ParOut[2]) );
  CKBD0 U120 ( .CLK(n124), .C(n119) );
  CKNXD16 U121 ( .I(n119), .ZN(ParOut[1]) );
  CKBD0 U122 ( .CLK(n123), .C(n121) );
  CKNXD16 U123 ( .I(n121), .ZN(ParOut[0]) );
  INVD1 U124 ( .I(n156), .ZN(n155) );
  BUFFD1 U125 ( .I(n157), .Z(n156) );
  INVD1 U126 ( .I(Reset), .ZN(n157) );
  NR2D1 U127 ( .A1(FIFOEmpty), .A2(n3), .ZN(N35) );
  INVD0 U128 ( .I(ReadReq), .ZN(n3) );
  CKAN2D0 U129 ( .A1(FIFO_Out[0]), .A2(ReadReq), .Z(N3) );
  CKAN2D0 U130 ( .A1(FIFO_Out[1]), .A2(ReadReq), .Z(N4) );
  CKAN2D0 U131 ( .A1(FIFO_Out[2]), .A2(ReadReq), .Z(N5) );
  CKAN2D0 U132 ( .A1(FIFO_Out[3]), .A2(ReadReq), .Z(N6) );
  CKAN2D0 U133 ( .A1(FIFO_Out[4]), .A2(ReadReq), .Z(N7) );
  CKAN2D0 U134 ( .A1(FIFO_Out[5]), .A2(ReadReq), .Z(N8) );
  CKAN2D0 U135 ( .A1(FIFO_Out[6]), .A2(ReadReq), .Z(N9) );
  CKAN2D0 U136 ( .A1(FIFO_Out[7]), .A2(ReadReq), .Z(N10) );
  CKAN2D0 U137 ( .A1(FIFO_Out[8]), .A2(ReadReq), .Z(N11) );
  CKAN2D0 U138 ( .A1(FIFO_Out[9]), .A2(ReadReq), .Z(N12) );
  CKAN2D0 U139 ( .A1(FIFO_Out[10]), .A2(ReadReq), .Z(N13) );
  CKAN2D0 U140 ( .A1(FIFO_Out[11]), .A2(ReadReq), .Z(N14) );
  CKAN2D0 U141 ( .A1(FIFO_Out[12]), .A2(ReadReq), .Z(N15) );
  CKAN2D0 U142 ( .A1(FIFO_Out[13]), .A2(ReadReq), .Z(N16) );
  CKAN2D0 U143 ( .A1(FIFO_Out[14]), .A2(ReadReq), .Z(N17) );
  CKAN2D0 U144 ( .A1(FIFO_Out[15]), .A2(ReadReq), .Z(N18) );
  CKAN2D0 U145 ( .A1(FIFO_Out[16]), .A2(ReadReq), .Z(N19) );
  CKAN2D0 U146 ( .A1(FIFO_Out[17]), .A2(ReadReq), .Z(N20) );
  CKAN2D0 U147 ( .A1(FIFO_Out[18]), .A2(ReadReq), .Z(N21) );
  CKAN2D0 U148 ( .A1(FIFO_Out[19]), .A2(ReadReq), .Z(N22) );
  CKAN2D0 U149 ( .A1(FIFO_Out[20]), .A2(ReadReq), .Z(N23) );
  CKAN2D0 U150 ( .A1(FIFO_Out[21]), .A2(ReadReq), .Z(N24) );
  CKAN2D0 U151 ( .A1(FIFO_Out[22]), .A2(ReadReq), .Z(N25) );
  CKAN2D0 U152 ( .A1(FIFO_Out[23]), .A2(ReadReq), .Z(N26) );
  CKAN2D0 U153 ( .A1(FIFO_Out[24]), .A2(ReadReq), .Z(N27) );
  CKAN2D0 U154 ( .A1(FIFO_Out[25]), .A2(ReadReq), .Z(N28) );
  CKAN2D0 U155 ( .A1(FIFO_Out[26]), .A2(ReadReq), .Z(N29) );
  CKAN2D0 U156 ( .A1(FIFO_Out[27]), .A2(ReadReq), .Z(N30) );
  CKAN2D0 U157 ( .A1(FIFO_Out[28]), .A2(ReadReq), .Z(N31) );
  CKAN2D0 U158 ( .A1(FIFO_Out[29]), .A2(ReadReq), .Z(N32) );
  CKAN2D0 U159 ( .A1(FIFO_Out[30]), .A2(ReadReq), .Z(N33) );
  CKAN2D0 U160 ( .A1(FIFO_Out[31]), .A2(ReadReq), .Z(N34) );
  CKND0 U161 ( .CLK(n189), .CN(n123) );
  CKND0 U162 ( .CLK(n188), .CN(n124) );
  CKND0 U163 ( .CLK(n187), .CN(n125) );
  CKND0 U164 ( .CLK(n186), .CN(n126) );
  CKND0 U165 ( .CLK(n185), .CN(n127) );
  CKND0 U166 ( .CLK(n184), .CN(n128) );
  CKND0 U167 ( .CLK(n183), .CN(n129) );
  CKND0 U168 ( .CLK(n182), .CN(n130) );
  CKND0 U169 ( .CLK(n181), .CN(n131) );
  CKND0 U170 ( .CLK(n180), .CN(n132) );
  CKND0 U171 ( .CLK(n179), .CN(n133) );
  CKND0 U172 ( .CLK(n178), .CN(n134) );
  CKND0 U173 ( .CLK(n177), .CN(n135) );
  CKND0 U174 ( .CLK(n176), .CN(n136) );
  CKND0 U175 ( .CLK(n175), .CN(n137) );
  CKND0 U176 ( .CLK(n174), .CN(n138) );
  CKND0 U177 ( .CLK(n173), .CN(n139) );
  CKND0 U178 ( .CLK(n172), .CN(n140) );
  CKND0 U179 ( .CLK(n171), .CN(n141) );
  CKND0 U180 ( .CLK(n170), .CN(n142) );
  CKND0 U181 ( .CLK(n169), .CN(n143) );
  CKND0 U182 ( .CLK(n168), .CN(n144) );
  CKND0 U183 ( .CLK(n167), .CN(n145) );
  CKND0 U184 ( .CLK(n166), .CN(n146) );
  CKND0 U185 ( .CLK(n165), .CN(n147) );
  CKND0 U186 ( .CLK(n164), .CN(n148) );
  CKND0 U187 ( .CLK(n163), .CN(n149) );
  CKND0 U188 ( .CLK(n162), .CN(n150) );
  CKND0 U189 ( .CLK(n161), .CN(n151) );
  CKND0 U190 ( .CLK(n160), .CN(n152) );
  CKND0 U191 ( .CLK(n159), .CN(n153) );
  CKND0 U192 ( .CLK(n158), .CN(n154) );
endmodule


module Serializer_DWid32_AWid4 ( SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk, 
        ParIn, InParValid, ParInClk, SendSerial, Reset );
  input [31:0] ParIn;
  input InParValid, ParInClk, SendSerial, Reset;
  output SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk;
  wire   F_Valid, SerEncReadReq, F_ReadReq, F_WriteReq, EncD_ToTx, n2, n1, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [31:0] FIFO_Out;

  FIFOTop_AWid4_DWid32_1 FIFO_Tx1 ( .Dout(FIFO_Out), .Din(ParIn), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(n1), .WriteIn(F_WriteReq), 
        .ClkR(ParInClk), .ClkW(ParInClk), .Reseter(n29) );
  SerEncoder_DWid32_1 SerEnc_Tx1 ( .SerOut(EncD_ToTx), .SerValid(SerValid), 
        .FIFO_ReadReq(SerEncReadReq), .ParIn(FIFO_Out), .F_Empty(FIFOEmpty), 
        .ParClk(ParInClk), .SerClk(SerClk), .ParValid(F_Valid), .Reset(n29) );
  SerialTx_1 SerTx_Tx1 ( .SerOut(SerOut), .SerClk(SerClk), .SerIn(EncD_ToTx), 
        .ParClk(ParInClk), .Reset(n29) );
  INR2XD0 U1 ( .A1(InParValid), .B1(FIFOFull), .ZN(F_WriteReq) );
  BUFFD0 U2 ( .I(n3), .Z(n1) );
  BUFFD0 U3 ( .I(n4), .Z(n3) );
  BUFFD0 U4 ( .I(n5), .Z(n4) );
  BUFFD0 U5 ( .I(n6), .Z(n5) );
  BUFFD0 U6 ( .I(n7), .Z(n6) );
  BUFFD0 U7 ( .I(n8), .Z(n7) );
  BUFFD0 U8 ( .I(n9), .Z(n8) );
  BUFFD0 U9 ( .I(n10), .Z(n9) );
  BUFFD0 U10 ( .I(n11), .Z(n10) );
  BUFFD0 U11 ( .I(n12), .Z(n11) );
  BUFFD0 U12 ( .I(n13), .Z(n12) );
  BUFFD0 U13 ( .I(n14), .Z(n13) );
  BUFFD0 U14 ( .I(n15), .Z(n14) );
  BUFFD0 U15 ( .I(n16), .Z(n15) );
  BUFFD0 U16 ( .I(n17), .Z(n16) );
  BUFFD0 U17 ( .I(n18), .Z(n17) );
  BUFFD0 U18 ( .I(n19), .Z(n18) );
  BUFFD0 U19 ( .I(n20), .Z(n19) );
  BUFFD0 U20 ( .I(n21), .Z(n20) );
  BUFFD0 U21 ( .I(n22), .Z(n21) );
  BUFFD0 U22 ( .I(n23), .Z(n22) );
  BUFFD0 U23 ( .I(n24), .Z(n23) );
  BUFFD0 U24 ( .I(n25), .Z(n24) );
  BUFFD0 U25 ( .I(n26), .Z(n25) );
  BUFFD0 U26 ( .I(n27), .Z(n26) );
  BUFFD0 U27 ( .I(n28), .Z(n27) );
  BUFFD0 U28 ( .I(F_ReadReq), .Z(n28) );
  INVD1 U29 ( .I(n30), .ZN(n29) );
  INVD1 U30 ( .I(Reset), .ZN(n30) );
  AN3D1 U31 ( .A1(n2), .A2(SendSerial), .A3(SerEncReadReq), .Z(F_ReadReq) );
  INVD1 U32 ( .I(FIFOEmpty), .ZN(n2) );
  NR2D1 U33 ( .A1(n29), .A2(FIFOEmpty), .ZN(F_Valid) );
endmodule


module Deserializer_AWid3_DWid32 ( ParOut, ParValid, DecoderParClk, FIFOEmpty, 
        FIFOFull, ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, N3, N4,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, ParValidDecode, SerialClk, SerRxToDecode, n3, n1, n2, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n55, n57, n59, n61, n63, n65, n67, n69,
         n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97,
         n99, n101, n103, n105, n107, n109, n111, n113, n115, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid3_DWid32_1 FIFO_Rx1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), 
        .Full(FIFOFull), .Empty(FIFOEmpty), .ReadIn(ReadReq), .WriteIn(
        ParValidDecode), .ClkR(ParOutClk), .ClkW(DecoderParClk), .Reseter(n149) );
  DesDecoder_DWid32_1 DesDec_Rx1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(n149) );
  SerialRx_1 SerRx_Rx1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(n149) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(n1), .CP(ParOutClk), .CDN(n151), .Q(n152) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(n2), .CP(ParOutClk), .CDN(n151), .Q(n153) );
  DFCNQD1 \ParBuf_reg[29]  ( .D(n4), .CP(ParOutClk), .CDN(n151), .Q(n154) );
  DFCNQD1 \ParBuf_reg[28]  ( .D(n5), .CP(ParOutClk), .CDN(n151), .Q(n155) );
  DFCNQD1 \ParBuf_reg[27]  ( .D(n6), .CP(ParOutClk), .CDN(n151), .Q(n156) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(n7), .CP(ParOutClk), .CDN(n151), .Q(n157) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(n8), .CP(ParOutClk), .CDN(n150), .Q(n158) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(n9), .CP(ParOutClk), .CDN(n151), .Q(n159) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(n10), .CP(ParOutClk), .CDN(n151), .Q(n160) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(n11), .CP(ParOutClk), .CDN(n151), .Q(n161) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(n12), .CP(ParOutClk), .CDN(n151), .Q(n162) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(n13), .CP(ParOutClk), .CDN(n151), .Q(n163) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(n14), .CP(ParOutClk), .CDN(n151), .Q(n164) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(n15), .CP(ParOutClk), .CDN(n151), .Q(n165) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(n16), .CP(ParOutClk), .CDN(n150), .Q(n166) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(n17), .CP(ParOutClk), .CDN(n150), .Q(n167) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(n18), .CP(ParOutClk), .CDN(n150), .Q(n168) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(n19), .CP(ParOutClk), .CDN(n150), .Q(n169) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(n20), .CP(ParOutClk), .CDN(n150), .Q(n170) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(n21), .CP(ParOutClk), .CDN(n150), .Q(n171) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(n22), .CP(ParOutClk), .CDN(n150), .Q(n172) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(n23), .CP(ParOutClk), .CDN(n151), .Q(n173) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(n24), .CP(ParOutClk), .CDN(n151), .Q(n174) );
  DFCNQD1 \ParBuf_reg[8]  ( .D(n25), .CP(ParOutClk), .CDN(n151), .Q(n175) );
  DFCNQD1 \ParBuf_reg[7]  ( .D(n26), .CP(ParOutClk), .CDN(n151), .Q(n176) );
  DFCNQD1 \ParBuf_reg[6]  ( .D(n27), .CP(ParOutClk), .CDN(n151), .Q(n177) );
  DFCNQD1 \ParBuf_reg[5]  ( .D(n28), .CP(ParOutClk), .CDN(n151), .Q(n178) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(n29), .CP(ParOutClk), .CDN(n150), .Q(n179) );
  DFCNQD1 \ParBuf_reg[3]  ( .D(n30), .CP(ParOutClk), .CDN(n150), .Q(n180) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(n31), .CP(ParOutClk), .CDN(n150), .Q(n181) );
  DFCNQD1 \ParBuf_reg[1]  ( .D(n32), .CP(ParOutClk), .CDN(n150), .Q(n182) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(n33), .CP(ParOutClk), .CDN(n150), .Q(n183) );
  DFCNQD1 ParValidr_reg ( .D(n34), .CP(ParOutClk), .CDN(n150), .Q(ParValid) );
  CKBD0 U3 ( .CLK(N34), .C(n1) );
  CKBD0 U4 ( .CLK(N33), .C(n2) );
  CKBD0 U5 ( .CLK(N32), .C(n4) );
  CKBD0 U6 ( .CLK(N31), .C(n5) );
  CKBD0 U7 ( .CLK(N30), .C(n6) );
  CKBD0 U8 ( .CLK(N29), .C(n7) );
  CKBD0 U9 ( .CLK(N28), .C(n8) );
  CKBD0 U10 ( .CLK(N27), .C(n9) );
  CKBD0 U11 ( .CLK(N26), .C(n10) );
  CKBD0 U12 ( .CLK(N25), .C(n11) );
  CKBD0 U13 ( .CLK(N24), .C(n12) );
  CKBD0 U14 ( .CLK(N23), .C(n13) );
  CKBD0 U15 ( .CLK(N22), .C(n14) );
  CKBD0 U16 ( .CLK(N21), .C(n15) );
  CKBD0 U17 ( .CLK(N20), .C(n16) );
  CKBD0 U18 ( .CLK(N19), .C(n17) );
  CKBD0 U19 ( .CLK(N18), .C(n18) );
  CKBD0 U20 ( .CLK(N17), .C(n19) );
  CKBD0 U21 ( .CLK(N16), .C(n20) );
  CKBD0 U22 ( .CLK(N15), .C(n21) );
  CKBD0 U23 ( .CLK(N14), .C(n22) );
  CKBD0 U24 ( .CLK(N13), .C(n23) );
  CKBD0 U25 ( .CLK(N12), .C(n24) );
  CKBD0 U26 ( .CLK(N11), .C(n25) );
  CKBD0 U27 ( .CLK(N10), .C(n26) );
  CKBD0 U28 ( .CLK(N9), .C(n27) );
  CKBD0 U29 ( .CLK(N8), .C(n28) );
  BUFFD0 U30 ( .I(N7), .Z(n29) );
  BUFFD0 U31 ( .I(N6), .Z(n30) );
  BUFFD0 U32 ( .I(N5), .Z(n31) );
  BUFFD0 U33 ( .I(N4), .Z(n32) );
  BUFFD0 U34 ( .I(N3), .Z(n33) );
  NR2D0 U35 ( .A1(FIFOEmpty), .A2(n3), .ZN(N35) );
  BUFFD0 U36 ( .I(n35), .Z(n34) );
  BUFFD0 U37 ( .I(n36), .Z(n35) );
  BUFFD0 U38 ( .I(n37), .Z(n36) );
  BUFFD0 U39 ( .I(n38), .Z(n37) );
  BUFFD0 U40 ( .I(n39), .Z(n38) );
  BUFFD0 U41 ( .I(n40), .Z(n39) );
  BUFFD0 U42 ( .I(n41), .Z(n40) );
  BUFFD0 U43 ( .I(n42), .Z(n41) );
  BUFFD0 U44 ( .I(n43), .Z(n42) );
  BUFFD0 U45 ( .I(n44), .Z(n43) );
  BUFFD0 U46 ( .I(n45), .Z(n44) );
  BUFFD0 U47 ( .I(n46), .Z(n45) );
  BUFFD0 U48 ( .I(n47), .Z(n46) );
  BUFFD0 U49 ( .I(n48), .Z(n47) );
  BUFFD0 U50 ( .I(n49), .Z(n48) );
  BUFFD0 U51 ( .I(n50), .Z(n49) );
  BUFFD0 U52 ( .I(n51), .Z(n50) );
  BUFFD0 U53 ( .I(n52), .Z(n51) );
  BUFFD0 U54 ( .I(N35), .Z(n52) );
  CKBD0 U55 ( .CLK(n148), .C(n53) );
  CKNXD16 U56 ( .I(n53), .ZN(ParOut[31]) );
  CKBD0 U57 ( .CLK(n147), .C(n55) );
  CKNXD16 U58 ( .I(n55), .ZN(ParOut[30]) );
  CKBD0 U59 ( .CLK(n146), .C(n57) );
  CKNXD16 U60 ( .I(n57), .ZN(ParOut[29]) );
  CKBD0 U61 ( .CLK(n145), .C(n59) );
  CKNXD16 U62 ( .I(n59), .ZN(ParOut[28]) );
  CKBD0 U63 ( .CLK(n144), .C(n61) );
  CKNXD16 U64 ( .I(n61), .ZN(ParOut[27]) );
  CKBD0 U65 ( .CLK(n143), .C(n63) );
  CKNXD16 U66 ( .I(n63), .ZN(ParOut[26]) );
  CKBD0 U67 ( .CLK(n142), .C(n65) );
  CKNXD16 U68 ( .I(n65), .ZN(ParOut[25]) );
  CKBD0 U69 ( .CLK(n141), .C(n67) );
  CKNXD16 U70 ( .I(n67), .ZN(ParOut[24]) );
  CKBD0 U71 ( .CLK(n140), .C(n69) );
  CKNXD16 U72 ( .I(n69), .ZN(ParOut[23]) );
  CKBD0 U73 ( .CLK(n139), .C(n71) );
  CKNXD16 U74 ( .I(n71), .ZN(ParOut[22]) );
  CKBD0 U75 ( .CLK(n138), .C(n73) );
  CKNXD16 U76 ( .I(n73), .ZN(ParOut[21]) );
  CKBD0 U77 ( .CLK(n137), .C(n75) );
  CKNXD16 U78 ( .I(n75), .ZN(ParOut[20]) );
  CKBD0 U79 ( .CLK(n136), .C(n77) );
  CKNXD16 U80 ( .I(n77), .ZN(ParOut[19]) );
  CKBD0 U81 ( .CLK(n135), .C(n79) );
  CKNXD16 U82 ( .I(n79), .ZN(ParOut[18]) );
  CKBD0 U83 ( .CLK(n134), .C(n81) );
  CKNXD16 U84 ( .I(n81), .ZN(ParOut[17]) );
  CKBD0 U85 ( .CLK(n133), .C(n83) );
  CKNXD16 U86 ( .I(n83), .ZN(ParOut[16]) );
  CKBD0 U87 ( .CLK(n132), .C(n85) );
  CKNXD16 U88 ( .I(n85), .ZN(ParOut[15]) );
  CKBD0 U89 ( .CLK(n131), .C(n87) );
  CKNXD16 U90 ( .I(n87), .ZN(ParOut[14]) );
  CKBD0 U91 ( .CLK(n130), .C(n89) );
  CKNXD16 U92 ( .I(n89), .ZN(ParOut[13]) );
  CKBD0 U93 ( .CLK(n129), .C(n91) );
  CKNXD16 U94 ( .I(n91), .ZN(ParOut[12]) );
  CKBD0 U95 ( .CLK(n128), .C(n93) );
  CKNXD16 U96 ( .I(n93), .ZN(ParOut[11]) );
  CKBD0 U97 ( .CLK(n127), .C(n95) );
  CKNXD16 U98 ( .I(n95), .ZN(ParOut[10]) );
  CKBD0 U99 ( .CLK(n126), .C(n97) );
  CKNXD16 U100 ( .I(n97), .ZN(ParOut[9]) );
  CKBD0 U101 ( .CLK(n125), .C(n99) );
  CKNXD16 U102 ( .I(n99), .ZN(ParOut[8]) );
  CKBD0 U103 ( .CLK(n124), .C(n101) );
  CKNXD16 U104 ( .I(n101), .ZN(ParOut[7]) );
  CKBD0 U105 ( .CLK(n123), .C(n103) );
  CKNXD16 U106 ( .I(n103), .ZN(ParOut[6]) );
  CKBD0 U107 ( .CLK(n122), .C(n105) );
  CKNXD16 U108 ( .I(n105), .ZN(ParOut[5]) );
  CKBD0 U109 ( .CLK(n121), .C(n107) );
  CKNXD16 U110 ( .I(n107), .ZN(ParOut[4]) );
  CKBD0 U111 ( .CLK(n120), .C(n109) );
  CKNXD16 U112 ( .I(n109), .ZN(ParOut[3]) );
  CKBD0 U113 ( .CLK(n119), .C(n111) );
  CKNXD16 U114 ( .I(n111), .ZN(ParOut[2]) );
  CKBD0 U115 ( .CLK(n118), .C(n113) );
  CKNXD16 U116 ( .I(n113), .ZN(ParOut[1]) );
  CKBD0 U117 ( .CLK(n117), .C(n115) );
  CKNXD16 U118 ( .I(n115), .ZN(ParOut[0]) );
  INVD1 U119 ( .I(n150), .ZN(n149) );
  BUFFD1 U120 ( .I(n151), .Z(n150) );
  INVD1 U121 ( .I(Reset), .ZN(n151) );
  INVD0 U122 ( .I(ReadReq), .ZN(n3) );
  CKAN2D0 U123 ( .A1(FIFO_Out[0]), .A2(ReadReq), .Z(N3) );
  CKAN2D0 U124 ( .A1(FIFO_Out[1]), .A2(ReadReq), .Z(N4) );
  CKAN2D0 U125 ( .A1(FIFO_Out[2]), .A2(ReadReq), .Z(N5) );
  CKAN2D0 U126 ( .A1(FIFO_Out[3]), .A2(ReadReq), .Z(N6) );
  CKAN2D0 U127 ( .A1(FIFO_Out[4]), .A2(ReadReq), .Z(N7) );
  CKAN2D0 U128 ( .A1(FIFO_Out[5]), .A2(ReadReq), .Z(N8) );
  CKAN2D0 U129 ( .A1(FIFO_Out[6]), .A2(ReadReq), .Z(N9) );
  CKAN2D0 U130 ( .A1(FIFO_Out[7]), .A2(ReadReq), .Z(N10) );
  CKAN2D0 U131 ( .A1(FIFO_Out[8]), .A2(ReadReq), .Z(N11) );
  CKAN2D0 U132 ( .A1(FIFO_Out[9]), .A2(ReadReq), .Z(N12) );
  CKAN2D0 U133 ( .A1(FIFO_Out[10]), .A2(ReadReq), .Z(N13) );
  CKAN2D0 U134 ( .A1(FIFO_Out[11]), .A2(ReadReq), .Z(N14) );
  CKAN2D0 U135 ( .A1(FIFO_Out[12]), .A2(ReadReq), .Z(N15) );
  CKAN2D0 U136 ( .A1(FIFO_Out[13]), .A2(ReadReq), .Z(N16) );
  CKAN2D0 U137 ( .A1(FIFO_Out[14]), .A2(ReadReq), .Z(N17) );
  CKAN2D0 U138 ( .A1(FIFO_Out[15]), .A2(ReadReq), .Z(N18) );
  CKAN2D0 U139 ( .A1(FIFO_Out[16]), .A2(ReadReq), .Z(N19) );
  CKAN2D0 U140 ( .A1(FIFO_Out[17]), .A2(ReadReq), .Z(N20) );
  CKAN2D0 U141 ( .A1(FIFO_Out[18]), .A2(ReadReq), .Z(N21) );
  CKAN2D0 U142 ( .A1(FIFO_Out[19]), .A2(ReadReq), .Z(N22) );
  CKAN2D0 U143 ( .A1(FIFO_Out[20]), .A2(ReadReq), .Z(N23) );
  CKAN2D0 U144 ( .A1(FIFO_Out[21]), .A2(ReadReq), .Z(N24) );
  CKAN2D0 U145 ( .A1(FIFO_Out[22]), .A2(ReadReq), .Z(N25) );
  CKAN2D0 U146 ( .A1(FIFO_Out[23]), .A2(ReadReq), .Z(N26) );
  CKAN2D0 U147 ( .A1(FIFO_Out[24]), .A2(ReadReq), .Z(N27) );
  CKAN2D0 U148 ( .A1(FIFO_Out[25]), .A2(ReadReq), .Z(N28) );
  CKAN2D0 U149 ( .A1(FIFO_Out[26]), .A2(ReadReq), .Z(N29) );
  CKAN2D0 U150 ( .A1(FIFO_Out[27]), .A2(ReadReq), .Z(N30) );
  CKAN2D0 U151 ( .A1(FIFO_Out[28]), .A2(ReadReq), .Z(N31) );
  CKAN2D0 U152 ( .A1(FIFO_Out[29]), .A2(ReadReq), .Z(N32) );
  CKAN2D0 U153 ( .A1(FIFO_Out[30]), .A2(ReadReq), .Z(N33) );
  CKAN2D0 U154 ( .A1(FIFO_Out[31]), .A2(ReadReq), .Z(N34) );
  CKND0 U155 ( .CLK(n183), .CN(n117) );
  CKND0 U156 ( .CLK(n182), .CN(n118) );
  CKND0 U157 ( .CLK(n181), .CN(n119) );
  CKND0 U158 ( .CLK(n180), .CN(n120) );
  CKND0 U159 ( .CLK(n179), .CN(n121) );
  CKND0 U160 ( .CLK(n178), .CN(n122) );
  CKND0 U161 ( .CLK(n177), .CN(n123) );
  CKND0 U162 ( .CLK(n176), .CN(n124) );
  CKND0 U163 ( .CLK(n175), .CN(n125) );
  CKND0 U164 ( .CLK(n174), .CN(n126) );
  CKND0 U165 ( .CLK(n173), .CN(n127) );
  CKND0 U166 ( .CLK(n172), .CN(n128) );
  CKND0 U167 ( .CLK(n171), .CN(n129) );
  CKND0 U168 ( .CLK(n170), .CN(n130) );
  CKND0 U169 ( .CLK(n169), .CN(n131) );
  CKND0 U170 ( .CLK(n168), .CN(n132) );
  CKND0 U171 ( .CLK(n167), .CN(n133) );
  CKND0 U172 ( .CLK(n166), .CN(n134) );
  CKND0 U173 ( .CLK(n165), .CN(n135) );
  CKND0 U174 ( .CLK(n164), .CN(n136) );
  CKND0 U175 ( .CLK(n163), .CN(n137) );
  CKND0 U176 ( .CLK(n162), .CN(n138) );
  CKND0 U177 ( .CLK(n161), .CN(n139) );
  CKND0 U178 ( .CLK(n160), .CN(n140) );
  CKND0 U179 ( .CLK(n159), .CN(n141) );
  CKND0 U180 ( .CLK(n158), .CN(n142) );
  CKND0 U181 ( .CLK(n157), .CN(n143) );
  CKND0 U182 ( .CLK(n156), .CN(n144) );
  CKND0 U183 ( .CLK(n155), .CN(n145) );
  CKND0 U184 ( .CLK(n154), .CN(n146) );
  CKND0 U185 ( .CLK(n153), .CN(n147) );
  CKND0 U186 ( .CLK(n152), .CN(n148) );
endmodule


module FIFOTop_AWid3_DWid32_0 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [2:0] SM_ReadAddr;
  wire   [2:0] SM_WriteAddr;

  FIFOStateM_AWid3_0 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid3_DWid32_0 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  INVD1 U2 ( .I(n3), .ZN(n2) );
  INVD1 U3 ( .I(Reseter), .ZN(n3) );
  BUFFD1 U4 ( .I(SM_MemReadCmd), .Z(n1) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module SerEncoder_DWid32_0 ( SerOut, SerValid, FIFO_ReadReq, ParIn, F_Empty, 
        ParClk, SerClk, ParValid, Reset );
  input [31:0] ParIn;
  input F_Empty, ParClk, SerClk, ParValid, Reset;
  output SerOut, SerValid, FIFO_ReadReq;
  wire   N2, N3, N4, N5, N6, HalfParClkr, \Sh_N[5] , N8, N9, N10, N11, N12,
         N13, N23, N24, N25, N26, N27, N28, N29, N31, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87;
  wire   [31:0] InBuf;

  SerEncoder_DWid32_0_DW01_dec_0 \ShifterBlock/sub_132  ( .A({n27, n48, n42, 
        n29, n45, n44}), .SUM({N13, N12, N11, N10, N9, N8}) );
  DFCNQD1 SerValidr_reg ( .D(n62), .CP(n20), .CDN(n69), .Q(SerValid) );
  DFCNQD1 HalfParClkr_reg ( .D(n5), .CP(ParClk), .CDN(n67), .Q(HalfParClkr) );
  DFCNQD1 \InBuf_reg[30]  ( .D(N83), .CP(HalfParClkr), .CDN(n67), .Q(InBuf[30]) );
  DFCNQD1 \InBuf_reg[29]  ( .D(N82), .CP(n20), .CDN(n67), .Q(InBuf[29]) );
  DFCNQD1 \InBuf_reg[26]  ( .D(N79), .CP(n20), .CDN(n68), .Q(InBuf[26]) );
  DFCNQD1 \InBuf_reg[25]  ( .D(N78), .CP(n20), .CDN(n68), .Q(InBuf[25]) );
  DFCNQD1 \InBuf_reg[22]  ( .D(N75), .CP(n64), .CDN(n68), .Q(InBuf[22]) );
  DFCNQD1 \InBuf_reg[21]  ( .D(N74), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[21]) );
  DFCNQD1 \InBuf_reg[18]  ( .D(N71), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[18]) );
  DFCNQD1 \InBuf_reg[17]  ( .D(N70), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[17]) );
  DFCNQD1 \InBuf_reg[14]  ( .D(N67), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[14]) );
  DFCNQD1 \InBuf_reg[13]  ( .D(N66), .CP(n64), .CDN(n69), .Q(InBuf[13]) );
  DFCNQD1 \InBuf_reg[10]  ( .D(N63), .CP(n20), .CDN(n69), .Q(InBuf[10]) );
  DFCNQD1 \InBuf_reg[9]  ( .D(N62), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[9])
         );
  DFCNQD1 \InBuf_reg[6]  ( .D(N59), .CP(n20), .CDN(n68), .Q(InBuf[6]) );
  DFCNQD1 \InBuf_reg[5]  ( .D(N58), .CP(HalfParClkr), .CDN(n67), .Q(InBuf[5])
         );
  DFCNQD1 \InBuf_reg[2]  ( .D(N55), .CP(n20), .CDN(n68), .Q(InBuf[2]) );
  DFCNQD1 \InBuf_reg[1]  ( .D(N54), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[1])
         );
  DFCNQD1 \InBuf_reg[31]  ( .D(N84), .CP(HalfParClkr), .CDN(n67), .Q(InBuf[31]) );
  DFCNQD1 \InBuf_reg[28]  ( .D(N81), .CP(n20), .CDN(n68), .Q(InBuf[28]) );
  DFCNQD1 \InBuf_reg[27]  ( .D(N80), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[27]) );
  DFCNQD1 \InBuf_reg[24]  ( .D(N77), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[24]) );
  DFCNQD1 \InBuf_reg[23]  ( .D(N76), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[23]) );
  DFCNQD1 \InBuf_reg[20]  ( .D(N73), .CP(n20), .CDN(n68), .Q(InBuf[20]) );
  DFCNQD1 \InBuf_reg[19]  ( .D(N72), .CP(n20), .CDN(n68), .Q(InBuf[19]) );
  DFCNQD1 \InBuf_reg[16]  ( .D(N69), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[16]) );
  DFCNQD1 \InBuf_reg[15]  ( .D(N68), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[15]) );
  DFCNQD1 \InBuf_reg[12]  ( .D(N65), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[12]) );
  DFCNQD1 \InBuf_reg[11]  ( .D(N64), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[11]) );
  DFCNQD1 \InBuf_reg[8]  ( .D(N61), .CP(HalfParClkr), .CDN(n67), .Q(InBuf[8])
         );
  DFCNQD1 \InBuf_reg[7]  ( .D(N60), .CP(n20), .CDN(n68), .Q(InBuf[7]) );
  DFCNQD1 \InBuf_reg[4]  ( .D(N57), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[4])
         );
  DFCNQD1 \InBuf_reg[3]  ( .D(N56), .CP(n20), .CDN(n67), .Q(InBuf[3]) );
  DFCNQD1 \InBuf_reg[0]  ( .D(N53), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[0])
         );
  DFCNQD1 \Sh_N_reg[5]  ( .D(N13), .CP(SerClk), .CDN(n67), .Q(\Sh_N[5] ) );
  DFCNQD1 \Sh_N_reg[4]  ( .D(N12), .CP(SerClk), .CDN(n67), .Q(N6) );
  DFCNQD1 \Sh_N_reg[2]  ( .D(N10), .CP(SerClk), .CDN(n67), .Q(N4) );
  DFCNQD1 \Sh_N_reg[3]  ( .D(N11), .CP(SerClk), .CDN(n67), .Q(N5) );
  DFCNQD1 \Sh_N_reg[1]  ( .D(N9), .CP(SerClk), .CDN(n67), .Q(N3) );
  DFCNQD1 \Sh_N_reg[0]  ( .D(N8), .CP(SerClk), .CDN(n67), .Q(N2) );
  DFCNQD1 SerOutr_reg ( .D(n41), .CP(SerClk), .CDN(n69), .Q(SerOut) );
  INVD0 U3 ( .I(n65), .ZN(n64) );
  INR2D1 U4 ( .A1(ParValid), .B1(F_Empty), .ZN(N85) );
  CKND0 U5 ( .CLK(n39), .CN(n66) );
  MUX2ND0 U6 ( .I0(n56), .I1(n57), .S(n47), .ZN(n1) );
  MUX2ND0 U7 ( .I0(n52), .I1(n53), .S(n47), .ZN(n2) );
  MUX2ND0 U8 ( .I0(n54), .I1(n55), .S(n47), .ZN(n3) );
  MUX2ND0 U9 ( .I0(n50), .I1(n51), .S(n47), .ZN(n4) );
  CKBD0 U10 ( .CLK(HalfParClkr), .C(n20) );
  BUFFD0 U11 ( .I(n7), .Z(n5) );
  BUFFD0 U12 ( .I(n64), .Z(n6) );
  BUFFD0 U13 ( .I(n8), .Z(n7) );
  BUFFD0 U14 ( .I(n10), .Z(n8) );
  BUFFD0 U15 ( .I(n6), .Z(n9) );
  BUFFD0 U16 ( .I(n12), .Z(n10) );
  BUFFD0 U17 ( .I(n9), .Z(n11) );
  BUFFD0 U18 ( .I(n16), .Z(n12) );
  BUFFD0 U19 ( .I(n11), .Z(n13) );
  BUFFD0 U20 ( .I(n66), .Z(n14) );
  BUFFD0 U21 ( .I(n13), .Z(n15) );
  BUFFD0 U22 ( .I(n18), .Z(n16) );
  BUFFD0 U23 ( .I(n15), .Z(n17) );
  BUFFD0 U24 ( .I(n21), .Z(n18) );
  BUFFD0 U25 ( .I(n17), .Z(n19) );
  BUFFD0 U26 ( .I(n37), .Z(n21) );
  BUFFD0 U27 ( .I(n20), .Z(n22) );
  BUFFD0 U28 ( .I(n22), .Z(n23) );
  BUFFD0 U29 ( .I(n23), .Z(n24) );
  BUFFD0 U30 ( .I(n24), .Z(n25) );
  CKBD0 U31 ( .CLK(\Sh_N[5] ), .C(n26) );
  BUFFD0 U32 ( .I(n43), .Z(n27) );
  BUFFD0 U33 ( .I(N6), .Z(n28) );
  CKBD0 U34 ( .CLK(n49), .C(n42) );
  CKBXD0 U35 ( .I(N5), .Z(n49) );
  BUFFD0 U36 ( .I(n47), .Z(n29) );
  CKBXD0 U37 ( .I(N4), .Z(n47) );
  CKBD0 U38 ( .CLK(N3), .C(n30) );
  CKBD0 U39 ( .CLK(n30), .C(n31) );
  CKBD0 U40 ( .CLK(n31), .C(n32) );
  CKBD0 U41 ( .CLK(N2), .C(n33) );
  CKBD0 U42 ( .CLK(n33), .C(n34) );
  CKBD0 U43 ( .CLK(n34), .C(n35) );
  CKBD0 U44 ( .CLK(n35), .C(n36) );
  BUFFD0 U45 ( .I(n40), .Z(n37) );
  BUFFD0 U46 ( .I(n25), .Z(n38) );
  BUFFD0 U47 ( .I(n19), .Z(n39) );
  BUFFD0 U48 ( .I(n14), .Z(n40) );
  BUFFD0 U49 ( .I(N31), .Z(n41) );
  CKBD0 U50 ( .CLK(n46), .C(n43) );
  CKBXD0 U51 ( .I(n26), .Z(n46) );
  CKBD0 U52 ( .CLK(n36), .C(n44) );
  CKBD0 U53 ( .CLK(n32), .C(n45) );
  OR2D0 U54 ( .A1(n44), .A2(n45), .Z(n71) );
  CKND2D0 U55 ( .A1(n45), .A2(n44), .ZN(n72) );
  CKBXD0 U56 ( .I(n28), .Z(n48) );
  INVD1 U57 ( .I(Reset), .ZN(n69) );
  INVD1 U58 ( .I(Reset), .ZN(n68) );
  INVD1 U59 ( .I(Reset), .ZN(n67) );
  INVD1 U60 ( .I(n63), .ZN(n62) );
  INVD1 U61 ( .I(n71), .ZN(n70) );
  AN2D1 U62 ( .A1(n47), .A2(n70), .Z(N26) );
  MUX4ND0 U63 ( .I0(InBuf[8]), .I1(InBuf[9]), .I2(InBuf[10]), .I3(InBuf[11]), 
        .S0(N2), .S1(N3), .ZN(n50) );
  MUX4ND0 U64 ( .I0(InBuf[12]), .I1(InBuf[13]), .I2(InBuf[14]), .I3(InBuf[15]), 
        .S0(N2), .S1(N3), .ZN(n51) );
  MUX4ND0 U65 ( .I0(InBuf[16]), .I1(InBuf[17]), .I2(InBuf[18]), .I3(InBuf[19]), 
        .S0(N2), .S1(N3), .ZN(n52) );
  MUX4ND0 U66 ( .I0(InBuf[20]), .I1(InBuf[21]), .I2(InBuf[22]), .I3(InBuf[23]), 
        .S0(N2), .S1(N3), .ZN(n53) );
  MUX4ND0 U67 ( .I0(InBuf[24]), .I1(InBuf[25]), .I2(InBuf[26]), .I3(InBuf[27]), 
        .S0(N2), .S1(N3), .ZN(n54) );
  MUX4ND0 U68 ( .I0(InBuf[28]), .I1(InBuf[29]), .I2(InBuf[30]), .I3(InBuf[31]), 
        .S0(N2), .S1(N3), .ZN(n55) );
  MUX4ND0 U69 ( .I0(InBuf[0]), .I1(InBuf[1]), .I2(InBuf[2]), .I3(InBuf[3]), 
        .S0(N2), .S1(N3), .ZN(n56) );
  MUX4ND0 U70 ( .I0(InBuf[4]), .I1(InBuf[5]), .I2(InBuf[6]), .I3(InBuf[7]), 
        .S0(N2), .S1(N3), .ZN(n57) );
  NR2D1 U71 ( .A1(n72), .A2(n47), .ZN(N24) );
  INVD1 U72 ( .I(N85), .ZN(n63) );
  INVD1 U73 ( .I(n38), .ZN(n65) );
  MUX2ND0 U74 ( .I0(n58), .I1(n59), .S(n48), .ZN(N29) );
  MUX2ND0 U75 ( .I0(n60), .I1(n61), .S(n48), .ZN(N27) );
  MUX2ND0 U76 ( .I0(n59), .I1(n58), .S(n48), .ZN(N25) );
  MUX2ND0 U77 ( .I0(n61), .I1(n60), .S(n48), .ZN(N23) );
  MUX2ND0 U78 ( .I0(n2), .I1(n3), .S(n49), .ZN(n59) );
  MUX2ND0 U79 ( .I0(n1), .I1(n4), .S(n49), .ZN(n58) );
  MUX2ND0 U80 ( .I0(n3), .I1(n1), .S(n49), .ZN(n61) );
  MUX2ND0 U81 ( .I0(n4), .I1(n2), .S(n49), .ZN(n60) );
  MUX2ND0 U82 ( .I0(n72), .I1(n71), .S(n47), .ZN(N28) );
  AN2D0 U83 ( .A1(ParIn[31]), .A2(N85), .Z(N84) );
  AN2D0 U84 ( .A1(ParIn[30]), .A2(n62), .Z(N83) );
  AN2D0 U85 ( .A1(ParIn[29]), .A2(N85), .Z(N82) );
  AN2D0 U86 ( .A1(ParIn[28]), .A2(n62), .Z(N81) );
  AN2D0 U87 ( .A1(ParIn[27]), .A2(N85), .Z(N80) );
  AN2D0 U88 ( .A1(ParIn[26]), .A2(N85), .Z(N79) );
  AN2D0 U89 ( .A1(ParIn[25]), .A2(N85), .Z(N78) );
  AN2D0 U90 ( .A1(ParIn[24]), .A2(N85), .Z(N77) );
  AN2D0 U91 ( .A1(ParIn[23]), .A2(n62), .Z(N76) );
  AN2D0 U92 ( .A1(ParIn[22]), .A2(n62), .Z(N75) );
  AN2D0 U93 ( .A1(ParIn[21]), .A2(n62), .Z(N74) );
  AN2D0 U94 ( .A1(ParIn[20]), .A2(n62), .Z(N73) );
  AN2D0 U95 ( .A1(ParIn[19]), .A2(n62), .Z(N72) );
  AN2D0 U96 ( .A1(ParIn[18]), .A2(n62), .Z(N71) );
  AN2D0 U97 ( .A1(ParIn[17]), .A2(n62), .Z(N70) );
  AN2D0 U98 ( .A1(ParIn[16]), .A2(N85), .Z(N69) );
  AN2D0 U99 ( .A1(ParIn[15]), .A2(N85), .Z(N68) );
  AN2D0 U100 ( .A1(ParIn[14]), .A2(N85), .Z(N67) );
  AN2D0 U101 ( .A1(ParIn[13]), .A2(N85), .Z(N66) );
  AN2D0 U102 ( .A1(ParIn[12]), .A2(N85), .Z(N65) );
  AN2D0 U103 ( .A1(ParIn[11]), .A2(N85), .Z(N64) );
  AN2D0 U104 ( .A1(ParIn[10]), .A2(n62), .Z(N63) );
  AN2D0 U105 ( .A1(ParIn[9]), .A2(N85), .Z(N62) );
  AN2D0 U106 ( .A1(ParIn[8]), .A2(N85), .Z(N61) );
  AN2D0 U107 ( .A1(ParIn[7]), .A2(n62), .Z(N60) );
  AN2D0 U108 ( .A1(ParIn[6]), .A2(n62), .Z(N59) );
  AN2D0 U109 ( .A1(ParIn[5]), .A2(n62), .Z(N58) );
  AN2D0 U110 ( .A1(ParIn[4]), .A2(n62), .Z(N57) );
  AN2D0 U111 ( .A1(ParIn[3]), .A2(n62), .Z(N56) );
  AN2D0 U112 ( .A1(ParIn[2]), .A2(n62), .Z(N55) );
  AN2D0 U113 ( .A1(ParIn[1]), .A2(n62), .Z(N54) );
  AN2D0 U114 ( .A1(ParIn[0]), .A2(n62), .Z(N53) );
  IND2D0 U115 ( .A1(n73), .B1(n74), .ZN(N31) );
  OAI21D0 U116 ( .A1(N23), .A2(n75), .B(n76), .ZN(n74) );
  MUX2ND0 U117 ( .I0(n77), .I1(n78), .S(n75), .ZN(n76) );
  MUX3ND0 U118 ( .I0(N25), .I1(n79), .I2(N24), .S0(n43), .S1(n80), .ZN(n78) );
  NR2D0 U119 ( .A1(n43), .A2(n49), .ZN(n80) );
  MUX2D0 U120 ( .I0(n81), .I1(N26), .S(n82), .Z(n79) );
  NR2D0 U121 ( .A1(n48), .A2(n49), .ZN(n82) );
  INR2D0 U122 ( .A1(N27), .B1(n48), .ZN(n81) );
  CKND0 U123 ( .CLK(n42), .CN(n77) );
  CKND2D0 U124 ( .A1(n83), .A2(n84), .ZN(n75) );
  MUX2ND0 U125 ( .I0(n85), .I1(n86), .S(n42), .ZN(n73) );
  CKND2D0 U126 ( .A1(N29), .A2(n87), .ZN(n86) );
  CKND2D0 U127 ( .A1(N28), .A2(n87), .ZN(n85) );
  NR2D0 U128 ( .A1(n84), .A2(n83), .ZN(n87) );
  CKND0 U129 ( .CLK(n48), .CN(n83) );
  CKND0 U130 ( .CLK(n43), .CN(n84) );
  INR3D0 U131 ( .A1(n62), .B1(Reset), .B2(n37), .ZN(FIFO_ReadReq) );
endmodule


module SerialTx_0 ( SerOut, SerClk, SerIn, ParClk, Reset );
  input SerIn, ParClk, Reset;
  output SerOut, SerClk;
  wire   n2;

  PLLTop_0 PLL_TxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerIn), .Z(SerOut) );
endmodule


module FIFOTop_AWid4_DWid32_0 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4;
  wire   [3:0] SM_ReadAddr;
  wire   [3:0] SM_WriteAddr;

  FIFOStateM_AWid4_0 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(n1), .ClkW(ClkW), .Reset(n3) );
  DPMem1kx32_AWid4_DWid32_0 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(n1), .ClkW(ClkW), .ChipEna(
        \*Logic1* ), .Read(n2), .Write(SM_MemWriteCmd), .Reset(n3) );
  CKBD0 U2 ( .CLK(SM_MemReadCmd), .C(n2) );
  BUFFD0 U3 ( .I(ClkR), .Z(n1) );
  INVD1 U4 ( .I(n4), .ZN(n3) );
  INVD1 U5 ( .I(Reseter), .ZN(n4) );
  TIEH U6 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32_0 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   SerClock, N30, N31, N32, N33, N34, N37, N38, N39, N40, N41, N42, N43,
         N47, n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n230, n231, n232, n1, n4, n5, n30, n31, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9026, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164;
  wire   [3:0] ParValidTimer;
  wire   [31:0] Decoder;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  MOAI22D1 U39 ( .A1(n9127), .A2(n54), .B1(n9129), .B2(Decoder[9]), .ZN(n123)
         );
  MOAI22D1 U40 ( .A1(n9127), .A2(n55), .B1(n9129), .B2(Decoder[8]), .ZN(n124)
         );
  OR3D1 U92 ( .A1(n8214), .A2(n8437), .A3(n8357), .Z(n22) );
  OR3D1 U94 ( .A1(n8342), .A2(n8345), .A3(n8359), .Z(n23) );
  OR3D1 U96 ( .A1(n8539), .A2(n8180), .A3(n8254), .Z(n24) );
  OA21D1 U99 ( .A1(n26), .A2(n27), .B(SerValid), .Z(N43) );
  OR2D1 U101 ( .A1(Count32[1]), .A2(Count32[0]), .Z(n28) );
  DesDecoder_DWid32_0_DW01_inc_0 \ClkGen/add_206  ( .A({Count32[4:2], n6727, 
        n6735}), .SUM({N34, N33, N32, N31, N30}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(n4), .CPN(n9149), .CDN(n9162), .Q(FrameSR[63]) );
  DFNCND1 \FrameSR_reg[22]  ( .D(n30), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[22]) );
  DFNCND1 \FrameSR_reg[23]  ( .D(n220), .CPN(n9154), .CDN(n9157), .Q(
        FrameSR[23]) );
  DFNCND1 \FrameSR_reg[37]  ( .D(n313), .CPN(n9152), .CDN(n9159), .Q(
        FrameSR[37]) );
  DFNCND1 \FrameSR_reg[38]  ( .D(n402), .CPN(n9152), .CDN(n9159), .Q(
        FrameSR[38]) );
  DFNCND1 \FrameSR_reg[53]  ( .D(n492), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[53]) );
  DFNCND1 \FrameSR_reg[54]  ( .D(n581), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[54]) );
  DFNCND1 \FrameSR_reg[32]  ( .D(n671), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[32]) );
  DFNCND1 \FrameSR_reg[39]  ( .D(n673), .CPN(n9152), .CDN(n9159), .Q(
        FrameSR[39]) );
  DFNCND1 \FrameSR_reg[55]  ( .D(n763), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[55]) );
  DFNCND1 \FrameSR_reg[8]  ( .D(n853), .CPN(n9155), .CDN(n9157), .Q(FrameSR[8]) );
  DFNCND1 \FrameSR_reg[9]  ( .D(n857), .CPN(n9155), .CDN(n9157), .Q(FrameSR[9]) );
  DFNCND1 \FrameSR_reg[10]  ( .D(n859), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[10]) );
  DFNCND1 \FrameSR_reg[11]  ( .D(n861), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[11]) );
  DFNCND1 \FrameSR_reg[12]  ( .D(n863), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[12]) );
  DFNCND1 \FrameSR_reg[13]  ( .D(n865), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[13]) );
  DFNCND1 \FrameSR_reg[14]  ( .D(n867), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[14]) );
  DFNCND1 \FrameSR_reg[15]  ( .D(n869), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[15]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(n871), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[19]) );
  DFNCND1 \FrameSR_reg[24]  ( .D(n960), .CPN(n9153), .CDN(n9160), .Q(
        FrameSR[24]) );
  DFNCND1 \FrameSR_reg[25]  ( .D(n1050), .CPN(n9153), .CDN(n9163), .Q(
        FrameSR[25]) );
  DFNCND1 \FrameSR_reg[26]  ( .D(n1052), .CPN(n9153), .CDN(n9162), .Q(
        FrameSR[26]) );
  DFNCND1 \FrameSR_reg[27]  ( .D(n1054), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[27]) );
  DFNCND1 \FrameSR_reg[28]  ( .D(n1056), .CPN(n9153), .CDN(n9161), .Q(
        FrameSR[28]) );
  DFNCND1 \FrameSR_reg[29]  ( .D(n1058), .CPN(n9153), .CDN(n9164), .Q(
        FrameSR[29]) );
  DFNCND1 \FrameSR_reg[30]  ( .D(n1060), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[30]) );
  DFNCND1 \FrameSR_reg[31]  ( .D(n1062), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[31]) );
  DFNCND1 \FrameSR_reg[40]  ( .D(n1064), .CPN(n9152), .CDN(n9163), .Q(
        FrameSR[40]) );
  DFNCND1 \FrameSR_reg[41]  ( .D(n1154), .CPN(n9152), .CDN(n9161), .Q(
        FrameSR[41]) );
  DFNCND1 \FrameSR_reg[42]  ( .D(n1156), .CPN(n9151), .CDN(n9159), .Q(
        FrameSR[42]) );
  DFNCND1 \FrameSR_reg[43]  ( .D(n1158), .CPN(n9151), .CDN(n9161), .Q(
        FrameSR[43]) );
  DFNCND1 \FrameSR_reg[44]  ( .D(n1160), .CPN(n9151), .CDN(n9162), .Q(
        FrameSR[44]) );
  DFNCND1 \FrameSR_reg[45]  ( .D(n1162), .CPN(n9151), .CDN(n9164), .Q(
        FrameSR[45]) );
  DFNCND1 \FrameSR_reg[46]  ( .D(n1164), .CPN(n9151), .CDN(n9162), .Q(
        FrameSR[46]) );
  DFNCND1 \FrameSR_reg[47]  ( .D(n1166), .CPN(n9151), .CDN(n9157), .Q(
        FrameSR[47]) );
  DFNCND1 \FrameSR_reg[56]  ( .D(n1168), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[56]) );
  DFNCND1 \FrameSR_reg[57]  ( .D(n1258), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[57]) );
  DFNCND1 \FrameSR_reg[58]  ( .D(n1260), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[58]) );
  DFNCND1 \FrameSR_reg[59]  ( .D(n1262), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[59]) );
  DFNCND1 \FrameSR_reg[60]  ( .D(n1264), .CPN(n9149), .CDN(n9160), .Q(
        FrameSR[60]) );
  DFNCND1 \FrameSR_reg[61]  ( .D(n1266), .CPN(n9149), .CDN(n9164), .Q(
        FrameSR[61]) );
  DFNCND1 \FrameSR_reg[62]  ( .D(n1268), .CPN(n9149), .CDN(n9162), .Q(
        FrameSR[62]) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[0]) );
  DFNCND1 \FrameSR_reg[4]  ( .D(n1270), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(n1273), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(n1361), .CPN(n9152), .CDN(n9159), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(n1450), .CPN(n9151), .CDN(n9158), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(n1539), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(n1542), .CPN(n9155), .CDN(n9157), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(n1546), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(n1635), .CPN(n9152), .CDN(n9159), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(n1725), .CPN(n9151), .CDN(n9160), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(n1727), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(n1730), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(n1733), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(n1736), .CPN(n9155), .CDN(n9157), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(n1740), .CPN(n9154), .CDN(n9157), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(n1829), .CPN(n9152), .CDN(n9159), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(n1918), .CPN(n9151), .CDN(n9160), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[51]  ( .D(n2007), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[51]) );
  DFNCND1 \FrameSR_reg[36]  ( .D(n2096), .CPN(n9152), .CDN(n9159), .Q(
        FrameSR[36]) );
  DFNCND1 \FrameSR_reg[52]  ( .D(n2185), .CPN(n9150), .CDN(n9160), .Q(
        FrameSR[52]) );
  DFNCND1 \FrameSR_reg[17]  ( .D(n2273), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[17]) );
  DFNCND1 \FrameSR_reg[16]  ( .D(n2362), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[16]) );
  EDFCNQD1 \Count32_reg[4]  ( .D(n2364), .E(SerValid), .CP(n9141), .CDN(n9163), 
        .Q(Count32[4]) );
  DFNCND1 \Decoder_reg[31]  ( .D(n2365), .CPN(n9149), .CDN(n9157), .Q(
        Decoder[31]) );
  DFNCND1 \Decoder_reg[30]  ( .D(n2499), .CPN(n9149), .CDN(n9163), .Q(
        Decoder[30]) );
  DFNCND1 \Decoder_reg[29]  ( .D(n2635), .CPN(n9149), .CDN(n9159), .Q(
        Decoder[29]) );
  DFNCND1 \Decoder_reg[28]  ( .D(n2771), .CPN(n9149), .CDN(n9161), .Q(
        Decoder[28]) );
  DFNCND1 \Decoder_reg[27]  ( .D(n2907), .CPN(n9149), .CDN(n9159), .Q(
        Decoder[27]) );
  DFNCND1 \Decoder_reg[26]  ( .D(n3043), .CPN(n9148), .CDN(n9164), .Q(
        Decoder[26]) );
  DFNCND1 \Decoder_reg[25]  ( .D(n3179), .CPN(n9148), .CDN(n9163), .Q(
        Decoder[25]) );
  DFNCND1 \Decoder_reg[24]  ( .D(n3315), .CPN(n9148), .CDN(n9157), .Q(
        Decoder[24]) );
  DFNCND1 \Decoder_reg[23]  ( .D(n3451), .CPN(n9148), .CDN(n9163), .Q(
        Decoder[23]) );
  DFNCND1 \Decoder_reg[22]  ( .D(n3587), .CPN(n9148), .CDN(n9163), .Q(
        Decoder[22]) );
  DFNCND1 \Decoder_reg[21]  ( .D(n3723), .CPN(n9148), .CDN(n9161), .Q(
        Decoder[21]) );
  DFNCND1 \Decoder_reg[20]  ( .D(n3859), .CPN(n9148), .CDN(n9161), .Q(
        Decoder[20]) );
  DFNCND1 \Decoder_reg[19]  ( .D(n3995), .CPN(n9148), .CDN(n9164), .Q(
        Decoder[19]) );
  DFNCND1 \Decoder_reg[18]  ( .D(n4131), .CPN(n9148), .CDN(n9158), .Q(
        Decoder[18]) );
  DFNCND1 \Decoder_reg[17]  ( .D(n4267), .CPN(n9147), .CDN(n9162), .Q(
        Decoder[17]) );
  DFNCND1 \Decoder_reg[16]  ( .D(n4403), .CPN(n9147), .CDN(n9163), .Q(
        Decoder[16]) );
  DFNCND1 \Decoder_reg[15]  ( .D(n4539), .CPN(n9147), .CDN(n9162), .Q(
        Decoder[15]) );
  DFNCND1 \Decoder_reg[14]  ( .D(n4675), .CPN(n9147), .CDN(n9163), .Q(
        Decoder[14]) );
  DFNCND1 \Decoder_reg[13]  ( .D(n4811), .CPN(n9147), .CDN(n9164), .Q(
        Decoder[13]) );
  DFNCND1 \Decoder_reg[12]  ( .D(n4947), .CPN(n9147), .CDN(n9164), .Q(
        Decoder[12]) );
  DFNCND1 \Decoder_reg[11]  ( .D(n5083), .CPN(n9147), .CDN(n9161), .Q(
        Decoder[11]) );
  DFNCND1 \Decoder_reg[10]  ( .D(n5219), .CPN(n9147), .CDN(n9158), .Q(
        Decoder[10]) );
  DFNCND1 \Decoder_reg[9]  ( .D(n5355), .CPN(n9147), .CDN(n9163), .Q(
        Decoder[9]) );
  DFNCND1 \Decoder_reg[8]  ( .D(n5492), .CPN(n9146), .CDN(n9161), .Q(
        Decoder[8]) );
  DFNCND1 \Decoder_reg[7]  ( .D(n5629), .CPN(n9146), .CDN(n9161), .Q(
        Decoder[7]) );
  DFNCND1 \Decoder_reg[6]  ( .D(n5765), .CPN(n9146), .CDN(n9162), .Q(
        Decoder[6]) );
  DFNCND1 \Decoder_reg[5]  ( .D(n5902), .CPN(n9146), .CDN(n9160), .Q(
        Decoder[5]) );
  DFNCND1 \Decoder_reg[4]  ( .D(n6039), .CPN(n9146), .CDN(n9160), .Q(
        Decoder[4]) );
  DFNCND1 \Decoder_reg[3]  ( .D(n6176), .CPN(n9146), .CDN(n9161), .Q(
        Decoder[3]) );
  DFNCND1 \Decoder_reg[2]  ( .D(n6313), .CPN(n9146), .CDN(n9159), .Q(
        Decoder[2]) );
  DFNCND1 \Decoder_reg[1]  ( .D(n6450), .CPN(n9146), .CDN(n9163), .Q(
        Decoder[1]) );
  DFNCND1 \Decoder_reg[0]  ( .D(n6587), .CPN(n9146), .CDN(n9158), .Q(
        Decoder[0]) );
  DFNCND1 \ParValidTimer_reg[1]  ( .D(n6724), .CPN(n9142), .CDN(n9163), .Q(
        ParValidTimer[1]) );
  EDFCNQD1 \Count32_reg[1]  ( .D(n6726), .E(SerValid), .CP(n9141), .CDN(n9163), 
        .Q(Count32[1]) );
  DFNCND1 \ParValidTimer_reg[0]  ( .D(n6728), .CPN(n9142), .CDN(n9160), .Q(
        ParValidTimer[0]) );
  EDFCNQD1 \Count32_reg[3]  ( .D(n6730), .E(SerValid), .CP(n9141), .CDN(n9158), 
        .Q(Count32[3]) );
  EDFCNQD1 \Count32_reg[2]  ( .D(n6732), .E(SerValid), .CP(n9141), .CDN(n9157), 
        .Q(Count32[2]) );
  EDFCNQD1 \Count32_reg[0]  ( .D(n6734), .E(SerValid), .CP(n9141), .CDN(n9159), 
        .Q(Count32[0]) );
  DFNCND1 \ParOutr_reg[0]  ( .D(n6736), .CPN(n9145), .CDN(n9163), .Q(ParOut[0]), .QN(n63) );
  DFNCND1 \ParOutr_reg[1]  ( .D(n6740), .CPN(n9145), .CDN(n9164), .Q(ParOut[1]), .QN(n62) );
  DFNCND1 \ParOutr_reg[2]  ( .D(n6744), .CPN(n9145), .CDN(n9161), .Q(ParOut[2]), .QN(n61) );
  DFNCND1 \ParOutr_reg[3]  ( .D(n6748), .CPN(n9145), .CDN(n9162), .Q(ParOut[3]), .QN(n60) );
  DFNCND1 \ParOutr_reg[4]  ( .D(n6752), .CPN(n9145), .CDN(n9161), .Q(ParOut[4]), .QN(n59) );
  DFNCND1 \ParOutr_reg[5]  ( .D(n6756), .CPN(n9145), .CDN(n9160), .Q(ParOut[5]), .QN(n58) );
  DFNCND1 \ParOutr_reg[6]  ( .D(n6760), .CPN(n9145), .CDN(n9164), .Q(ParOut[6]), .QN(n57) );
  DFNCND1 \ParOutr_reg[7]  ( .D(n6764), .CPN(n9144), .CDN(n9162), .Q(ParOut[7]), .QN(n56) );
  DFNCND1 \ParOutr_reg[8]  ( .D(n6768), .CPN(n9144), .CDN(n9164), .Q(ParOut[8]), .QN(n55) );
  DFNCND1 \ParOutr_reg[9]  ( .D(n6772), .CPN(n9144), .CDN(n9157), .Q(ParOut[9]), .QN(n54) );
  DFNCND1 \ParOutr_reg[10]  ( .D(n6776), .CPN(n9144), .CDN(n9163), .Q(
        ParOut[10]), .QN(n53) );
  DFNCND1 \ParOutr_reg[11]  ( .D(n6780), .CPN(n9144), .CDN(n9162), .Q(
        ParOut[11]), .QN(n52) );
  DFNCND1 \ParOutr_reg[12]  ( .D(n6784), .CPN(n9144), .CDN(n9160), .Q(
        ParOut[12]), .QN(n51) );
  DFNCND1 \ParOutr_reg[13]  ( .D(n6788), .CPN(n9144), .CDN(n9163), .Q(
        ParOut[13]), .QN(n50) );
  DFNCND1 \ParOutr_reg[14]  ( .D(n6792), .CPN(n9144), .CDN(n9161), .Q(
        ParOut[14]), .QN(n49) );
  DFNCND1 \ParOutr_reg[15]  ( .D(n6796), .CPN(n9144), .CDN(n9162), .Q(
        ParOut[15]), .QN(n48) );
  DFNCND1 \ParOutr_reg[16]  ( .D(n6800), .CPN(n9143), .CDN(n9164), .Q(
        ParOut[16]), .QN(n47) );
  DFNCND1 \ParOutr_reg[17]  ( .D(n6804), .CPN(n9143), .CDN(n9159), .Q(
        ParOut[17]), .QN(n46) );
  DFNCND1 \ParOutr_reg[18]  ( .D(n6808), .CPN(n9143), .CDN(n9159), .Q(
        ParOut[18]), .QN(n45) );
  DFNCND1 \ParOutr_reg[19]  ( .D(n6812), .CPN(n9143), .CDN(n9158), .Q(
        ParOut[19]), .QN(n44) );
  DFNCND1 \ParOutr_reg[20]  ( .D(n6816), .CPN(n9143), .CDN(n9157), .Q(
        ParOut[20]), .QN(n43) );
  DFNCND1 \ParOutr_reg[21]  ( .D(n6820), .CPN(n9143), .CDN(n9164), .Q(
        ParOut[21]), .QN(n42) );
  DFNCND1 \ParOutr_reg[22]  ( .D(n6824), .CPN(n9143), .CDN(n9162), .Q(
        ParOut[22]), .QN(n41) );
  DFNCND1 \ParOutr_reg[23]  ( .D(n6828), .CPN(n9143), .CDN(n9161), .Q(
        ParOut[23]), .QN(n40) );
  DFNCND1 \ParOutr_reg[24]  ( .D(n6832), .CPN(n9143), .CDN(n9161), .Q(
        ParOut[24]), .QN(n39) );
  DFNCND1 \ParOutr_reg[25]  ( .D(n6836), .CPN(n9142), .CDN(n9164), .Q(
        ParOut[25]), .QN(n38) );
  DFNCND1 \ParOutr_reg[26]  ( .D(n6840), .CPN(n9142), .CDN(n9161), .Q(
        ParOut[26]), .QN(n37) );
  DFNCND1 \ParOutr_reg[27]  ( .D(n6844), .CPN(n9142), .CDN(n9162), .Q(
        ParOut[27]), .QN(n36) );
  DFNCND1 \ParOutr_reg[28]  ( .D(n6848), .CPN(n9142), .CDN(n9162), .Q(
        ParOut[28]), .QN(n35) );
  DFNCND1 \ParOutr_reg[29]  ( .D(n6852), .CPN(n9142), .CDN(n9161), .Q(
        ParOut[29]), .QN(n34) );
  DFNCND1 \ParOutr_reg[30]  ( .D(n6856), .CPN(n9142), .CDN(n9162), .Q(
        ParOut[30]), .QN(n33) );
  DFNCND1 \ParOutr_reg[31]  ( .D(n6860), .CPN(n9142), .CDN(n9163), .Q(
        ParOut[31]), .QN(n32) );
  EDFCNQD1 ParClkr_reg ( .D(n6864), .E(n6866), .CP(n9141), .CDN(n9161), .Q(
        ParClk) );
  DFNCND1 ParValidr_reg ( .D(n6868), .CPN(n9141), .CDN(n9162), .Q(ParValid), 
        .QN(n29) );
  DFNCND1 doParSync_reg ( .D(N47), .CPN(n9145), .CDN(n9164), .Q(n27), .QN(n2)
         );
  DFNCND1 UnLoad_reg ( .D(n9001), .CPN(n9145), .CDN(n9164), .Q(n1), .QN(n231)
         );
  DFNCND1 \ParValidTimer_reg[3]  ( .D(n9018), .CPN(n9141), .CDN(n9164), .QN(
        n232) );
  DFNCND1 \ParValidTimer_reg[2]  ( .D(n9021), .CPN(n9141), .CDN(n9164), .QN(
        n230) );
  IOA22D0 U3 ( .B1(n9128), .B2(n32), .A1(n1), .A2(Decoder[31]), .ZN(n101) );
  AO22D0 U4 ( .A1(n5491), .A2(n9125), .B1(Decoder[9]), .B2(n9126), .Z(n142) );
  CKAN2D0 U5 ( .A1(N30), .A2(n2), .Z(N38) );
  INVD0 U6 ( .I(ParValidTimer[0]), .ZN(n6) );
  BUFFD0 U7 ( .I(n2634), .Z(n4) );
  CKBD0 U8 ( .CLK(FrameSR[62]), .C(n5) );
  BUFFD0 U9 ( .I(n8398), .Z(n30) );
  CKBD0 U10 ( .CLK(FrameSR[21]), .C(n31) );
  BUFFD0 U11 ( .I(n31), .Z(n64) );
  CKBD0 U12 ( .CLK(n64), .C(n65) );
  CKBD0 U13 ( .CLK(n65), .C(n66) );
  CKBD0 U14 ( .CLK(n66), .C(n67) );
  CKBD0 U15 ( .CLK(n67), .C(n68) );
  CKBD0 U16 ( .CLK(n68), .C(n69) );
  CKBD0 U17 ( .CLK(n69), .C(n70) );
  CKBD0 U18 ( .CLK(n70), .C(n71) );
  CKBD0 U19 ( .CLK(n71), .C(n72) );
  CKBD0 U20 ( .CLK(n72), .C(n73) );
  CKBD0 U21 ( .CLK(n73), .C(n74) );
  BUFFD0 U22 ( .I(n74), .Z(n75) );
  CKBD0 U23 ( .CLK(n75), .C(n76) );
  CKBD0 U24 ( .CLK(n76), .C(n77) );
  CKBD0 U25 ( .CLK(n77), .C(n78) );
  CKBD0 U26 ( .CLK(n78), .C(n79) );
  CKBD0 U27 ( .CLK(n79), .C(n80) );
  CKBD0 U28 ( .CLK(n80), .C(n81) );
  CKBD0 U29 ( .CLK(n81), .C(n82) );
  CKBD0 U30 ( .CLK(n82), .C(n83) );
  CKBD0 U31 ( .CLK(n83), .C(n84) );
  CKBD0 U32 ( .CLK(n84), .C(n85) );
  BUFFD0 U33 ( .I(n85), .Z(n86) );
  CKBD0 U34 ( .CLK(n86), .C(n87) );
  CKBD0 U35 ( .CLK(n87), .C(n88) );
  CKBD0 U36 ( .CLK(n88), .C(n89) );
  CKBD0 U37 ( .CLK(n89), .C(n90) );
  CKBD0 U38 ( .CLK(n90), .C(n91) );
  CKBD0 U41 ( .CLK(n91), .C(n92) );
  CKBD0 U42 ( .CLK(n92), .C(n93) );
  CKBD0 U43 ( .CLK(n93), .C(n94) );
  CKBD0 U44 ( .CLK(n94), .C(n95) );
  CKBD0 U45 ( .CLK(n95), .C(n165) );
  BUFFD0 U46 ( .I(n165), .Z(n166) );
  CKBD0 U47 ( .CLK(n166), .C(n167) );
  CKBD0 U48 ( .CLK(n167), .C(n168) );
  CKBD0 U49 ( .CLK(n168), .C(n169) );
  CKBD0 U50 ( .CLK(n169), .C(n170) );
  CKBD0 U51 ( .CLK(n170), .C(n171) );
  CKBD0 U52 ( .CLK(n171), .C(n172) );
  CKBD0 U53 ( .CLK(n172), .C(n173) );
  CKBD0 U54 ( .CLK(n173), .C(n174) );
  CKBD0 U55 ( .CLK(n174), .C(n175) );
  CKBD0 U56 ( .CLK(n175), .C(n176) );
  BUFFD0 U57 ( .I(n176), .Z(n177) );
  CKBD0 U58 ( .CLK(n177), .C(n178) );
  CKBD0 U59 ( .CLK(n178), .C(n179) );
  CKBD0 U60 ( .CLK(n179), .C(n180) );
  CKBD0 U61 ( .CLK(n180), .C(n181) );
  CKBD0 U62 ( .CLK(n181), .C(n182) );
  CKBD0 U63 ( .CLK(n182), .C(n183) );
  CKBD0 U64 ( .CLK(n183), .C(n184) );
  CKBD0 U65 ( .CLK(n184), .C(n185) );
  CKBD0 U66 ( .CLK(n185), .C(n186) );
  CKBD0 U67 ( .CLK(n186), .C(n187) );
  BUFFD0 U68 ( .I(n187), .Z(n188) );
  CKBD0 U69 ( .CLK(n188), .C(n189) );
  CKBD0 U70 ( .CLK(n189), .C(n190) );
  CKBD0 U71 ( .CLK(n190), .C(n191) );
  CKBD0 U72 ( .CLK(n191), .C(n192) );
  CKBD0 U73 ( .CLK(n192), .C(n193) );
  CKBD0 U74 ( .CLK(n193), .C(n194) );
  CKBD0 U75 ( .CLK(n194), .C(n195) );
  CKBD0 U76 ( .CLK(n195), .C(n196) );
  CKBD0 U77 ( .CLK(n196), .C(n197) );
  BUFFD0 U78 ( .I(n197), .Z(n198) );
  CKBD0 U79 ( .CLK(n198), .C(n199) );
  CKBD0 U80 ( .CLK(n199), .C(n200) );
  CKBD0 U81 ( .CLK(n200), .C(n201) );
  CKBD0 U82 ( .CLK(n201), .C(n202) );
  CKBD0 U83 ( .CLK(n202), .C(n203) );
  CKBD0 U84 ( .CLK(n203), .C(n204) );
  CKBD0 U85 ( .CLK(n204), .C(n205) );
  CKBD0 U86 ( .CLK(n205), .C(n206) );
  CKBD0 U87 ( .CLK(n206), .C(n207) );
  CKBD0 U88 ( .CLK(n207), .C(n208) );
  BUFFD0 U89 ( .I(n208), .Z(n209) );
  CKBD0 U90 ( .CLK(n209), .C(n210) );
  CKBD0 U91 ( .CLK(n210), .C(n211) );
  CKBD0 U93 ( .CLK(n211), .C(n212) );
  CKBD0 U95 ( .CLK(n212), .C(n213) );
  CKBD0 U97 ( .CLK(n213), .C(n214) );
  CKBD0 U98 ( .CLK(n214), .C(n215) );
  CKBD0 U100 ( .CLK(n215), .C(n216) );
  CKBD0 U102 ( .CLK(n216), .C(n217) );
  CKBD0 U103 ( .CLK(n217), .C(n218) );
  CKBD0 U104 ( .CLK(n218), .C(n219) );
  BUFFD0 U105 ( .I(n8254), .Z(n220) );
  CKBD0 U106 ( .CLK(FrameSR[22]), .C(n221) );
  CKBD0 U107 ( .CLK(n221), .C(n222) );
  CKBD0 U108 ( .CLK(n222), .C(n223) );
  CKBD0 U109 ( .CLK(n223), .C(n224) );
  CKBD0 U110 ( .CLK(n224), .C(n225) );
  CKBD0 U111 ( .CLK(n225), .C(n226) );
  CKBD0 U112 ( .CLK(n226), .C(n227) );
  BUFFD0 U113 ( .I(n227), .Z(n228) );
  CKBD0 U114 ( .CLK(n228), .C(n229) );
  CKBD0 U115 ( .CLK(n229), .C(n233) );
  CKBD0 U116 ( .CLK(n233), .C(n234) );
  CKBD0 U117 ( .CLK(n234), .C(n235) );
  CKBD0 U118 ( .CLK(n235), .C(n236) );
  CKBD0 U119 ( .CLK(n236), .C(n237) );
  CKBD0 U120 ( .CLK(n237), .C(n238) );
  CKBD0 U121 ( .CLK(n238), .C(n239) );
  CKBD0 U122 ( .CLK(n239), .C(n240) );
  CKBD0 U123 ( .CLK(n240), .C(n241) );
  BUFFD0 U124 ( .I(n241), .Z(n242) );
  CKBD0 U125 ( .CLK(n242), .C(n243) );
  CKBD0 U126 ( .CLK(n243), .C(n244) );
  CKBD0 U127 ( .CLK(n244), .C(n245) );
  CKBD0 U128 ( .CLK(n245), .C(n246) );
  CKBD0 U129 ( .CLK(n246), .C(n247) );
  CKBD0 U130 ( .CLK(n247), .C(n248) );
  CKBD0 U131 ( .CLK(n248), .C(n249) );
  CKBD0 U132 ( .CLK(n249), .C(n250) );
  CKBD0 U133 ( .CLK(n250), .C(n251) );
  CKBD0 U134 ( .CLK(n251), .C(n252) );
  BUFFD0 U135 ( .I(n252), .Z(n253) );
  CKBD0 U136 ( .CLK(n253), .C(n254) );
  CKBD0 U137 ( .CLK(n254), .C(n255) );
  CKBD0 U138 ( .CLK(n255), .C(n256) );
  CKBD0 U139 ( .CLK(n256), .C(n257) );
  CKBD0 U140 ( .CLK(n257), .C(n258) );
  CKBD0 U141 ( .CLK(n258), .C(n259) );
  CKBD0 U142 ( .CLK(n259), .C(n260) );
  CKBD0 U143 ( .CLK(n260), .C(n261) );
  CKBD0 U144 ( .CLK(n261), .C(n262) );
  CKBD0 U145 ( .CLK(n262), .C(n263) );
  BUFFD0 U146 ( .I(n263), .Z(n264) );
  CKBD0 U147 ( .CLK(n264), .C(n265) );
  CKBD0 U148 ( .CLK(n265), .C(n266) );
  CKBD0 U149 ( .CLK(n266), .C(n267) );
  CKBD0 U150 ( .CLK(n267), .C(n268) );
  CKBD0 U151 ( .CLK(n268), .C(n269) );
  CKBD0 U152 ( .CLK(n269), .C(n270) );
  CKBD0 U153 ( .CLK(n270), .C(n271) );
  CKBD0 U154 ( .CLK(n271), .C(n272) );
  CKBD0 U155 ( .CLK(n272), .C(n273) );
  CKBD0 U156 ( .CLK(n273), .C(n274) );
  BUFFD0 U157 ( .I(n274), .Z(n275) );
  CKBD0 U158 ( .CLK(n275), .C(n276) );
  CKBD0 U159 ( .CLK(n276), .C(n277) );
  CKBD0 U160 ( .CLK(n277), .C(n278) );
  CKBD0 U161 ( .CLK(n278), .C(n279) );
  CKBD0 U162 ( .CLK(n279), .C(n280) );
  CKBD0 U163 ( .CLK(n280), .C(n281) );
  CKBD0 U164 ( .CLK(n281), .C(n282) );
  CKBD0 U165 ( .CLK(n282), .C(n283) );
  CKBD0 U166 ( .CLK(n283), .C(n284) );
  CKBD0 U167 ( .CLK(n284), .C(n285) );
  BUFFD0 U168 ( .I(n285), .Z(n286) );
  CKBD0 U169 ( .CLK(n286), .C(n287) );
  CKBD0 U170 ( .CLK(n287), .C(n288) );
  CKBD0 U171 ( .CLK(n288), .C(n289) );
  CKBD0 U172 ( .CLK(n289), .C(n290) );
  CKBD0 U173 ( .CLK(n290), .C(n291) );
  CKBD0 U174 ( .CLK(n291), .C(n292) );
  CKBD0 U175 ( .CLK(n292), .C(n293) );
  CKBD0 U176 ( .CLK(n293), .C(n294) );
  CKBD0 U177 ( .CLK(n294), .C(n295) );
  BUFFD0 U178 ( .I(n295), .Z(n296) );
  CKBD0 U179 ( .CLK(n296), .C(n297) );
  CKBD0 U180 ( .CLK(n297), .C(n298) );
  CKBD0 U181 ( .CLK(n298), .C(n299) );
  CKBD0 U182 ( .CLK(n299), .C(n300) );
  CKBD0 U183 ( .CLK(n300), .C(n301) );
  CKBD0 U184 ( .CLK(n301), .C(n302) );
  CKBD0 U185 ( .CLK(n302), .C(n303) );
  CKBD0 U186 ( .CLK(n303), .C(n304) );
  CKBD0 U187 ( .CLK(n304), .C(n305) );
  CKBD0 U188 ( .CLK(n305), .C(n306) );
  BUFFD0 U189 ( .I(n306), .Z(n307) );
  CKBD0 U190 ( .CLK(n307), .C(n308) );
  CKBD0 U191 ( .CLK(n308), .C(n309) );
  CKBD0 U192 ( .CLK(n309), .C(n310) );
  CKBD0 U193 ( .CLK(n310), .C(n311) );
  CKBD0 U194 ( .CLK(n311), .C(n312) );
  BUFFD0 U195 ( .I(n8373), .Z(n313) );
  CKBD0 U196 ( .CLK(FrameSR[36]), .C(n314) );
  CKBD0 U197 ( .CLK(n314), .C(n315) );
  CKBD0 U198 ( .CLK(n315), .C(n316) );
  CKBD0 U199 ( .CLK(n316), .C(n317) );
  CKBD0 U200 ( .CLK(n317), .C(n318) );
  CKBD0 U201 ( .CLK(n318), .C(n319) );
  CKBD0 U202 ( .CLK(n319), .C(n320) );
  BUFFD0 U203 ( .I(n320), .Z(n321) );
  CKBD0 U204 ( .CLK(n321), .C(n322) );
  CKBD0 U205 ( .CLK(n322), .C(n323) );
  CKBD0 U206 ( .CLK(n323), .C(n324) );
  CKBD0 U207 ( .CLK(n324), .C(n325) );
  CKBD0 U208 ( .CLK(n325), .C(n326) );
  CKBD0 U209 ( .CLK(n326), .C(n327) );
  CKBD0 U210 ( .CLK(n327), .C(n328) );
  CKBD0 U211 ( .CLK(n328), .C(n329) );
  CKBD0 U212 ( .CLK(n329), .C(n330) );
  CKBD0 U213 ( .CLK(n330), .C(n331) );
  BUFFD0 U214 ( .I(n331), .Z(n332) );
  CKBD0 U215 ( .CLK(n332), .C(n333) );
  CKBD0 U216 ( .CLK(n333), .C(n334) );
  CKBD0 U217 ( .CLK(n334), .C(n335) );
  CKBD0 U218 ( .CLK(n335), .C(n336) );
  CKBD0 U219 ( .CLK(n336), .C(n337) );
  CKBD0 U220 ( .CLK(n337), .C(n338) );
  CKBD0 U221 ( .CLK(n338), .C(n339) );
  CKBD0 U222 ( .CLK(n339), .C(n340) );
  CKBD0 U223 ( .CLK(n340), .C(n341) );
  CKBD0 U224 ( .CLK(n341), .C(n342) );
  BUFFD0 U225 ( .I(n342), .Z(n343) );
  CKBD0 U226 ( .CLK(n343), .C(n344) );
  CKBD0 U227 ( .CLK(n344), .C(n345) );
  CKBD0 U228 ( .CLK(n345), .C(n346) );
  CKBD0 U229 ( .CLK(n346), .C(n347) );
  CKBD0 U230 ( .CLK(n347), .C(n348) );
  CKBD0 U231 ( .CLK(n348), .C(n349) );
  CKBD0 U232 ( .CLK(n349), .C(n350) );
  CKBD0 U233 ( .CLK(n350), .C(n351) );
  CKBD0 U234 ( .CLK(n351), .C(n352) );
  CKBD0 U235 ( .CLK(n352), .C(n353) );
  BUFFD0 U236 ( .I(n353), .Z(n354) );
  CKBD0 U237 ( .CLK(n354), .C(n355) );
  CKBD0 U238 ( .CLK(n355), .C(n356) );
  CKBD0 U239 ( .CLK(n356), .C(n357) );
  CKBD0 U240 ( .CLK(n357), .C(n358) );
  CKBD0 U241 ( .CLK(n358), .C(n359) );
  CKBD0 U242 ( .CLK(n359), .C(n360) );
  CKBD0 U243 ( .CLK(n360), .C(n361) );
  CKBD0 U244 ( .CLK(n361), .C(n362) );
  CKBD0 U245 ( .CLK(n362), .C(n363) );
  CKBD0 U246 ( .CLK(n363), .C(n364) );
  BUFFD0 U247 ( .I(n364), .Z(n365) );
  CKBD0 U248 ( .CLK(n365), .C(n366) );
  CKBD0 U249 ( .CLK(n366), .C(n367) );
  CKBD0 U250 ( .CLK(n367), .C(n368) );
  CKBD0 U251 ( .CLK(n368), .C(n369) );
  CKBD0 U252 ( .CLK(n369), .C(n370) );
  CKBD0 U253 ( .CLK(n370), .C(n371) );
  CKBD0 U254 ( .CLK(n371), .C(n372) );
  CKBD0 U255 ( .CLK(n372), .C(n373) );
  CKBD0 U256 ( .CLK(n373), .C(n374) );
  CKBD0 U257 ( .CLK(n374), .C(n375) );
  BUFFD0 U258 ( .I(n375), .Z(n376) );
  CKBD0 U259 ( .CLK(n376), .C(n377) );
  CKBD0 U260 ( .CLK(n377), .C(n378) );
  CKBD0 U261 ( .CLK(n378), .C(n379) );
  CKBD0 U262 ( .CLK(n379), .C(n380) );
  CKBD0 U263 ( .CLK(n380), .C(n381) );
  CKBD0 U264 ( .CLK(n381), .C(n382) );
  CKBD0 U265 ( .CLK(n382), .C(n383) );
  CKBD0 U266 ( .CLK(n383), .C(n384) );
  CKBD0 U267 ( .CLK(n384), .C(n385) );
  BUFFD0 U268 ( .I(n385), .Z(n386) );
  CKBD0 U269 ( .CLK(n386), .C(n387) );
  CKBD0 U270 ( .CLK(n387), .C(n388) );
  CKBD0 U271 ( .CLK(n388), .C(n389) );
  CKBD0 U272 ( .CLK(n389), .C(n390) );
  CKBD0 U273 ( .CLK(n390), .C(n391) );
  CKBD0 U274 ( .CLK(n391), .C(n392) );
  CKBD0 U275 ( .CLK(n392), .C(n393) );
  CKBD0 U276 ( .CLK(n393), .C(n394) );
  CKBD0 U277 ( .CLK(n394), .C(n395) );
  CKBD0 U278 ( .CLK(n395), .C(n396) );
  BUFFD0 U279 ( .I(n396), .Z(n397) );
  CKBD0 U280 ( .CLK(n397), .C(n398) );
  CKBD0 U281 ( .CLK(n398), .C(n399) );
  CKBD0 U282 ( .CLK(n399), .C(n400) );
  CKBD0 U283 ( .CLK(n400), .C(n401) );
  BUFFD0 U284 ( .I(n8359), .Z(n402) );
  CKBD0 U285 ( .CLK(FrameSR[37]), .C(n403) );
  CKBD0 U286 ( .CLK(n403), .C(n404) );
  CKBD0 U287 ( .CLK(n404), .C(n405) );
  CKBD0 U288 ( .CLK(n405), .C(n406) );
  CKBD0 U289 ( .CLK(n406), .C(n407) );
  CKBD0 U290 ( .CLK(n407), .C(n408) );
  CKBD0 U291 ( .CLK(n408), .C(n409) );
  BUFFD0 U292 ( .I(n409), .Z(n410) );
  CKBD0 U293 ( .CLK(n410), .C(n411) );
  CKBD0 U294 ( .CLK(n411), .C(n412) );
  CKBD0 U295 ( .CLK(n412), .C(n413) );
  CKBD0 U296 ( .CLK(n413), .C(n414) );
  CKBD0 U297 ( .CLK(n414), .C(n415) );
  CKBD0 U298 ( .CLK(n415), .C(n416) );
  CKBD0 U299 ( .CLK(n416), .C(n417) );
  CKBD0 U300 ( .CLK(n417), .C(n418) );
  CKBD0 U301 ( .CLK(n418), .C(n419) );
  CKBD0 U302 ( .CLK(n419), .C(n420) );
  BUFFD0 U303 ( .I(n420), .Z(n421) );
  CKBD0 U304 ( .CLK(n421), .C(n422) );
  CKBD0 U305 ( .CLK(n422), .C(n423) );
  CKBD0 U306 ( .CLK(n423), .C(n424) );
  CKBD0 U307 ( .CLK(n424), .C(n425) );
  CKBD0 U308 ( .CLK(n425), .C(n426) );
  CKBD0 U309 ( .CLK(n426), .C(n427) );
  CKBD0 U310 ( .CLK(n427), .C(n428) );
  CKBD0 U311 ( .CLK(n428), .C(n429) );
  CKBD0 U312 ( .CLK(n429), .C(n430) );
  CKBD0 U313 ( .CLK(n430), .C(n431) );
  BUFFD0 U314 ( .I(n431), .Z(n432) );
  CKBD0 U315 ( .CLK(n432), .C(n433) );
  CKBD0 U316 ( .CLK(n433), .C(n434) );
  CKBD0 U317 ( .CLK(n434), .C(n435) );
  CKBD0 U318 ( .CLK(n435), .C(n436) );
  CKBD0 U319 ( .CLK(n436), .C(n437) );
  CKBD0 U320 ( .CLK(n437), .C(n438) );
  CKBD0 U321 ( .CLK(n438), .C(n439) );
  CKBD0 U322 ( .CLK(n439), .C(n440) );
  CKBD0 U323 ( .CLK(n440), .C(n441) );
  CKBD0 U324 ( .CLK(n441), .C(n442) );
  BUFFD0 U325 ( .I(n442), .Z(n443) );
  CKBD0 U326 ( .CLK(n443), .C(n444) );
  CKBD0 U327 ( .CLK(n444), .C(n445) );
  CKBD0 U328 ( .CLK(n445), .C(n446) );
  CKBD0 U329 ( .CLK(n446), .C(n447) );
  CKBD0 U330 ( .CLK(n447), .C(n448) );
  CKBD0 U331 ( .CLK(n448), .C(n449) );
  CKBD0 U332 ( .CLK(n449), .C(n450) );
  CKBD0 U333 ( .CLK(n450), .C(n451) );
  CKBD0 U334 ( .CLK(n451), .C(n452) );
  CKBD0 U335 ( .CLK(n452), .C(n453) );
  BUFFD0 U336 ( .I(n453), .Z(n454) );
  CKBD0 U337 ( .CLK(n454), .C(n455) );
  CKBD0 U338 ( .CLK(n455), .C(n456) );
  CKBD0 U339 ( .CLK(n456), .C(n457) );
  CKBD0 U340 ( .CLK(n457), .C(n458) );
  CKBD0 U341 ( .CLK(n458), .C(n459) );
  CKBD0 U342 ( .CLK(n459), .C(n460) );
  CKBD0 U343 ( .CLK(n460), .C(n461) );
  CKBD0 U344 ( .CLK(n461), .C(n462) );
  CKBD0 U345 ( .CLK(n462), .C(n463) );
  CKBD0 U346 ( .CLK(n463), .C(n464) );
  BUFFD0 U347 ( .I(n464), .Z(n465) );
  CKBD0 U348 ( .CLK(n465), .C(n466) );
  CKBD0 U349 ( .CLK(n466), .C(n467) );
  CKBD0 U350 ( .CLK(n467), .C(n468) );
  CKBD0 U351 ( .CLK(n468), .C(n469) );
  CKBD0 U352 ( .CLK(n469), .C(n470) );
  CKBD0 U353 ( .CLK(n470), .C(n471) );
  CKBD0 U354 ( .CLK(n471), .C(n472) );
  CKBD0 U355 ( .CLK(n472), .C(n473) );
  CKBD0 U356 ( .CLK(n473), .C(n474) );
  BUFFD0 U357 ( .I(n474), .Z(n475) );
  CKBD0 U358 ( .CLK(n475), .C(n476) );
  CKBD0 U359 ( .CLK(n476), .C(n477) );
  CKBD0 U360 ( .CLK(n477), .C(n478) );
  CKBD0 U361 ( .CLK(n478), .C(n479) );
  CKBD0 U362 ( .CLK(n479), .C(n480) );
  CKBD0 U363 ( .CLK(n480), .C(n481) );
  CKBD0 U364 ( .CLK(n481), .C(n482) );
  CKBD0 U365 ( .CLK(n482), .C(n483) );
  CKBD0 U366 ( .CLK(n483), .C(n484) );
  CKBD0 U367 ( .CLK(n484), .C(n485) );
  BUFFD0 U368 ( .I(n485), .Z(n486) );
  CKBD0 U369 ( .CLK(n486), .C(n487) );
  CKBD0 U370 ( .CLK(n487), .C(n488) );
  CKBD0 U371 ( .CLK(n488), .C(n489) );
  CKBD0 U372 ( .CLK(n489), .C(n490) );
  CKBD0 U373 ( .CLK(n490), .C(n491) );
  BUFFD0 U374 ( .I(n8680), .Z(n492) );
  CKBD0 U375 ( .CLK(FrameSR[52]), .C(n493) );
  CKBD0 U376 ( .CLK(n493), .C(n494) );
  CKBD0 U377 ( .CLK(n494), .C(n495) );
  CKBD0 U378 ( .CLK(n495), .C(n496) );
  CKBD0 U379 ( .CLK(n496), .C(n497) );
  CKBD0 U380 ( .CLK(n497), .C(n498) );
  BUFFD0 U381 ( .I(n498), .Z(n499) );
  CKBD0 U382 ( .CLK(n499), .C(n500) );
  CKBD0 U383 ( .CLK(n500), .C(n501) );
  CKBD0 U384 ( .CLK(n501), .C(n502) );
  CKBD0 U385 ( .CLK(n502), .C(n503) );
  CKBD0 U386 ( .CLK(n503), .C(n504) );
  CKBD0 U387 ( .CLK(n504), .C(n505) );
  CKBD0 U388 ( .CLK(n505), .C(n506) );
  CKBD0 U389 ( .CLK(n506), .C(n507) );
  CKBD0 U390 ( .CLK(n507), .C(n508) );
  CKBD0 U391 ( .CLK(n508), .C(n509) );
  BUFFD0 U392 ( .I(n509), .Z(n510) );
  CKBD0 U393 ( .CLK(n510), .C(n511) );
  CKBD0 U394 ( .CLK(n511), .C(n512) );
  CKBD0 U395 ( .CLK(n512), .C(n513) );
  CKBD0 U396 ( .CLK(n513), .C(n514) );
  CKBD0 U397 ( .CLK(n514), .C(n515) );
  CKBD0 U398 ( .CLK(n515), .C(n516) );
  CKBD0 U399 ( .CLK(n516), .C(n517) );
  CKBD0 U400 ( .CLK(n517), .C(n518) );
  CKBD0 U401 ( .CLK(n518), .C(n519) );
  BUFFD0 U402 ( .I(n519), .Z(n520) );
  CKBD0 U403 ( .CLK(n520), .C(n521) );
  CKBD0 U404 ( .CLK(n521), .C(n522) );
  CKBD0 U405 ( .CLK(n522), .C(n523) );
  CKBD0 U406 ( .CLK(n523), .C(n524) );
  CKBD0 U407 ( .CLK(n524), .C(n525) );
  CKBD0 U408 ( .CLK(n525), .C(n526) );
  CKBD0 U409 ( .CLK(n526), .C(n527) );
  CKBD0 U410 ( .CLK(n527), .C(n528) );
  CKBD0 U411 ( .CLK(n528), .C(n529) );
  CKBD0 U412 ( .CLK(n529), .C(n530) );
  BUFFD0 U413 ( .I(n530), .Z(n531) );
  CKBD0 U414 ( .CLK(n531), .C(n532) );
  CKBD0 U415 ( .CLK(n532), .C(n533) );
  CKBD0 U416 ( .CLK(n533), .C(n534) );
  CKBD0 U417 ( .CLK(n534), .C(n535) );
  CKBD0 U418 ( .CLK(n535), .C(n536) );
  CKBD0 U419 ( .CLK(n536), .C(n537) );
  CKBD0 U420 ( .CLK(n537), .C(n538) );
  CKBD0 U421 ( .CLK(n538), .C(n539) );
  CKBD0 U422 ( .CLK(n539), .C(n540) );
  CKBD0 U423 ( .CLK(n540), .C(n541) );
  BUFFD0 U424 ( .I(n541), .Z(n542) );
  CKBD0 U425 ( .CLK(n542), .C(n543) );
  CKBD0 U426 ( .CLK(n543), .C(n544) );
  CKBD0 U427 ( .CLK(n544), .C(n545) );
  CKBD0 U428 ( .CLK(n545), .C(n546) );
  CKBD0 U429 ( .CLK(n546), .C(n547) );
  CKBD0 U430 ( .CLK(n547), .C(n548) );
  CKBD0 U431 ( .CLK(n548), .C(n549) );
  CKBD0 U432 ( .CLK(n549), .C(n550) );
  CKBD0 U433 ( .CLK(n550), .C(n551) );
  CKBD0 U434 ( .CLK(n551), .C(n552) );
  BUFFD0 U435 ( .I(n552), .Z(n553) );
  CKBD0 U436 ( .CLK(n553), .C(n554) );
  CKBD0 U437 ( .CLK(n554), .C(n555) );
  CKBD0 U438 ( .CLK(n555), .C(n556) );
  CKBD0 U439 ( .CLK(n556), .C(n557) );
  CKBD0 U440 ( .CLK(n557), .C(n558) );
  CKBD0 U441 ( .CLK(n558), .C(n559) );
  CKBD0 U442 ( .CLK(n559), .C(n560) );
  CKBD0 U443 ( .CLK(n560), .C(n561) );
  CKBD0 U444 ( .CLK(n561), .C(n562) );
  CKBD0 U445 ( .CLK(n562), .C(n563) );
  BUFFD0 U446 ( .I(n563), .Z(n564) );
  CKBD0 U447 ( .CLK(n564), .C(n565) );
  CKBD0 U448 ( .CLK(n565), .C(n566) );
  CKBD0 U449 ( .CLK(n566), .C(n567) );
  CKBD0 U450 ( .CLK(n567), .C(n568) );
  CKBD0 U451 ( .CLK(n568), .C(n569) );
  CKBD0 U452 ( .CLK(n569), .C(n570) );
  CKBD0 U453 ( .CLK(n570), .C(n571) );
  CKBD0 U454 ( .CLK(n571), .C(n572) );
  CKBD0 U455 ( .CLK(n572), .C(n573) );
  CKBD0 U456 ( .CLK(n573), .C(n574) );
  BUFFD0 U457 ( .I(n574), .Z(n575) );
  CKBD0 U458 ( .CLK(n575), .C(n576) );
  CKBD0 U459 ( .CLK(n576), .C(n577) );
  CKBD0 U460 ( .CLK(n577), .C(n578) );
  CKBD0 U461 ( .CLK(n578), .C(n579) );
  CKBD0 U462 ( .CLK(n579), .C(n580) );
  BUFFD0 U463 ( .I(n8357), .Z(n581) );
  CKBD0 U464 ( .CLK(FrameSR[53]), .C(n582) );
  CKBD0 U465 ( .CLK(n582), .C(n583) );
  CKBD0 U466 ( .CLK(n583), .C(n584) );
  CKBD0 U467 ( .CLK(n584), .C(n585) );
  CKBD0 U468 ( .CLK(n585), .C(n586) );
  CKBD0 U469 ( .CLK(n586), .C(n587) );
  CKBD0 U470 ( .CLK(n587), .C(n588) );
  BUFFD0 U471 ( .I(n588), .Z(n589) );
  CKBD0 U472 ( .CLK(n589), .C(n590) );
  CKBD0 U473 ( .CLK(n590), .C(n591) );
  CKBD0 U474 ( .CLK(n591), .C(n592) );
  CKBD0 U475 ( .CLK(n592), .C(n593) );
  CKBD0 U476 ( .CLK(n593), .C(n594) );
  CKBD0 U477 ( .CLK(n594), .C(n595) );
  CKBD0 U478 ( .CLK(n595), .C(n596) );
  CKBD0 U479 ( .CLK(n596), .C(n597) );
  CKBD0 U480 ( .CLK(n597), .C(n598) );
  CKBD0 U481 ( .CLK(n598), .C(n599) );
  BUFFD0 U482 ( .I(n599), .Z(n600) );
  CKBD0 U483 ( .CLK(n600), .C(n601) );
  CKBD0 U484 ( .CLK(n601), .C(n602) );
  CKBD0 U485 ( .CLK(n602), .C(n603) );
  CKBD0 U486 ( .CLK(n603), .C(n604) );
  CKBD0 U487 ( .CLK(n604), .C(n605) );
  CKBD0 U488 ( .CLK(n605), .C(n606) );
  CKBD0 U489 ( .CLK(n606), .C(n607) );
  CKBD0 U490 ( .CLK(n607), .C(n608) );
  CKBD0 U491 ( .CLK(n608), .C(n609) );
  CKBD0 U492 ( .CLK(n609), .C(n610) );
  BUFFD0 U493 ( .I(n610), .Z(n611) );
  CKBD0 U494 ( .CLK(n611), .C(n612) );
  CKBD0 U495 ( .CLK(n612), .C(n613) );
  CKBD0 U496 ( .CLK(n613), .C(n614) );
  CKBD0 U497 ( .CLK(n614), .C(n615) );
  CKBD0 U498 ( .CLK(n615), .C(n616) );
  CKBD0 U499 ( .CLK(n616), .C(n617) );
  CKBD0 U500 ( .CLK(n617), .C(n618) );
  CKBD0 U501 ( .CLK(n618), .C(n619) );
  CKBD0 U502 ( .CLK(n619), .C(n620) );
  CKBD0 U503 ( .CLK(n620), .C(n621) );
  BUFFD0 U504 ( .I(n621), .Z(n622) );
  CKBD0 U505 ( .CLK(n622), .C(n623) );
  CKBD0 U506 ( .CLK(n623), .C(n624) );
  CKBD0 U507 ( .CLK(n624), .C(n625) );
  CKBD0 U508 ( .CLK(n625), .C(n626) );
  CKBD0 U509 ( .CLK(n626), .C(n627) );
  CKBD0 U510 ( .CLK(n627), .C(n628) );
  CKBD0 U511 ( .CLK(n628), .C(n629) );
  CKBD0 U512 ( .CLK(n629), .C(n630) );
  CKBD0 U513 ( .CLK(n630), .C(n631) );
  CKBD0 U514 ( .CLK(n631), .C(n632) );
  BUFFD0 U515 ( .I(n632), .Z(n633) );
  CKBD0 U516 ( .CLK(n633), .C(n634) );
  CKBD0 U517 ( .CLK(n634), .C(n635) );
  CKBD0 U518 ( .CLK(n635), .C(n636) );
  CKBD0 U519 ( .CLK(n636), .C(n637) );
  CKBD0 U520 ( .CLK(n637), .C(n638) );
  CKBD0 U521 ( .CLK(n638), .C(n639) );
  CKBD0 U522 ( .CLK(n639), .C(n640) );
  CKBD0 U523 ( .CLK(n640), .C(n641) );
  CKBD0 U524 ( .CLK(n641), .C(n642) );
  CKBD0 U525 ( .CLK(n642), .C(n643) );
  BUFFD0 U526 ( .I(n643), .Z(n644) );
  CKBD0 U527 ( .CLK(n644), .C(n645) );
  CKBD0 U528 ( .CLK(n645), .C(n646) );
  CKBD0 U529 ( .CLK(n646), .C(n647) );
  CKBD0 U530 ( .CLK(n647), .C(n648) );
  CKBD0 U531 ( .CLK(n648), .C(n649) );
  CKBD0 U532 ( .CLK(n649), .C(n650) );
  CKBD0 U533 ( .CLK(n650), .C(n651) );
  CKBD0 U534 ( .CLK(n651), .C(n652) );
  CKBD0 U535 ( .CLK(n652), .C(n653) );
  BUFFD0 U536 ( .I(n653), .Z(n654) );
  CKBD0 U537 ( .CLK(n654), .C(n655) );
  CKBD0 U538 ( .CLK(n655), .C(n656) );
  CKBD0 U539 ( .CLK(n656), .C(n657) );
  CKBD0 U540 ( .CLK(n657), .C(n658) );
  CKBD0 U541 ( .CLK(n658), .C(n659) );
  CKBD0 U542 ( .CLK(n659), .C(n660) );
  CKBD0 U543 ( .CLK(n660), .C(n661) );
  CKBD0 U544 ( .CLK(n661), .C(n662) );
  CKBD0 U545 ( .CLK(n662), .C(n663) );
  CKBD0 U546 ( .CLK(n663), .C(n664) );
  BUFFD0 U547 ( .I(n664), .Z(n665) );
  CKBD0 U548 ( .CLK(n665), .C(n666) );
  CKBD0 U549 ( .CLK(n666), .C(n667) );
  CKBD0 U550 ( .CLK(n667), .C(n668) );
  CKBD0 U551 ( .CLK(n668), .C(n669) );
  CKBD0 U552 ( .CLK(n669), .C(n670) );
  BUFFD0 U553 ( .I(n4674), .Z(n671) );
  CKBD0 U554 ( .CLK(FrameSR[31]), .C(n672) );
  BUFFD0 U555 ( .I(n8345), .Z(n673) );
  CKBD0 U556 ( .CLK(FrameSR[38]), .C(n674) );
  CKBD0 U557 ( .CLK(n674), .C(n675) );
  CKBD0 U558 ( .CLK(n675), .C(n676) );
  CKBD0 U559 ( .CLK(n676), .C(n677) );
  CKBD0 U560 ( .CLK(n677), .C(n678) );
  CKBD0 U561 ( .CLK(n678), .C(n679) );
  CKBD0 U562 ( .CLK(n679), .C(n680) );
  BUFFD0 U563 ( .I(n680), .Z(n681) );
  CKBD0 U564 ( .CLK(n681), .C(n682) );
  CKBD0 U565 ( .CLK(n682), .C(n683) );
  CKBD0 U566 ( .CLK(n683), .C(n684) );
  CKBD0 U567 ( .CLK(n684), .C(n685) );
  CKBD0 U568 ( .CLK(n685), .C(n686) );
  CKBD0 U569 ( .CLK(n686), .C(n687) );
  CKBD0 U570 ( .CLK(n687), .C(n688) );
  CKBD0 U571 ( .CLK(n688), .C(n689) );
  CKBD0 U572 ( .CLK(n689), .C(n690) );
  CKBD0 U573 ( .CLK(n690), .C(n691) );
  BUFFD0 U574 ( .I(n691), .Z(n692) );
  CKBD0 U575 ( .CLK(n692), .C(n693) );
  CKBD0 U576 ( .CLK(n693), .C(n694) );
  CKBD0 U577 ( .CLK(n694), .C(n695) );
  CKBD0 U578 ( .CLK(n695), .C(n696) );
  CKBD0 U579 ( .CLK(n696), .C(n697) );
  CKBD0 U580 ( .CLK(n697), .C(n698) );
  CKBD0 U581 ( .CLK(n698), .C(n699) );
  CKBD0 U582 ( .CLK(n699), .C(n700) );
  CKBD0 U583 ( .CLK(n700), .C(n701) );
  CKBD0 U584 ( .CLK(n701), .C(n702) );
  BUFFD0 U585 ( .I(n702), .Z(n703) );
  CKBD0 U586 ( .CLK(n703), .C(n704) );
  CKBD0 U587 ( .CLK(n704), .C(n705) );
  CKBD0 U588 ( .CLK(n705), .C(n706) );
  CKBD0 U589 ( .CLK(n706), .C(n707) );
  CKBD0 U590 ( .CLK(n707), .C(n708) );
  CKBD0 U591 ( .CLK(n708), .C(n709) );
  CKBD0 U592 ( .CLK(n709), .C(n710) );
  CKBD0 U593 ( .CLK(n710), .C(n711) );
  CKBD0 U594 ( .CLK(n711), .C(n712) );
  CKBD0 U595 ( .CLK(n712), .C(n713) );
  BUFFD0 U596 ( .I(n713), .Z(n714) );
  CKBD0 U597 ( .CLK(n714), .C(n715) );
  CKBD0 U598 ( .CLK(n715), .C(n716) );
  CKBD0 U599 ( .CLK(n716), .C(n717) );
  CKBD0 U600 ( .CLK(n717), .C(n718) );
  CKBD0 U601 ( .CLK(n718), .C(n719) );
  CKBD0 U602 ( .CLK(n719), .C(n720) );
  CKBD0 U603 ( .CLK(n720), .C(n721) );
  CKBD0 U604 ( .CLK(n721), .C(n722) );
  CKBD0 U605 ( .CLK(n722), .C(n723) );
  CKBD0 U606 ( .CLK(n723), .C(n724) );
  BUFFD0 U607 ( .I(n724), .Z(n725) );
  CKBD0 U608 ( .CLK(n725), .C(n726) );
  CKBD0 U609 ( .CLK(n726), .C(n727) );
  CKBD0 U610 ( .CLK(n727), .C(n728) );
  CKBD0 U611 ( .CLK(n728), .C(n729) );
  CKBD0 U612 ( .CLK(n729), .C(n730) );
  CKBD0 U613 ( .CLK(n730), .C(n731) );
  CKBD0 U614 ( .CLK(n731), .C(n732) );
  CKBD0 U615 ( .CLK(n732), .C(n733) );
  CKBD0 U616 ( .CLK(n733), .C(n734) );
  CKBD0 U617 ( .CLK(n734), .C(n735) );
  BUFFD0 U618 ( .I(n735), .Z(n736) );
  CKBD0 U619 ( .CLK(n736), .C(n737) );
  CKBD0 U620 ( .CLK(n737), .C(n738) );
  CKBD0 U621 ( .CLK(n738), .C(n739) );
  CKBD0 U622 ( .CLK(n739), .C(n740) );
  CKBD0 U623 ( .CLK(n740), .C(n741) );
  CKBD0 U624 ( .CLK(n741), .C(n742) );
  CKBD0 U625 ( .CLK(n742), .C(n743) );
  CKBD0 U626 ( .CLK(n743), .C(n744) );
  CKBD0 U627 ( .CLK(n744), .C(n745) );
  BUFFD0 U628 ( .I(n745), .Z(n746) );
  CKBD0 U629 ( .CLK(n746), .C(n747) );
  CKBD0 U630 ( .CLK(n747), .C(n748) );
  CKBD0 U631 ( .CLK(n748), .C(n749) );
  CKBD0 U632 ( .CLK(n749), .C(n750) );
  CKBD0 U633 ( .CLK(n750), .C(n751) );
  CKBD0 U634 ( .CLK(n751), .C(n752) );
  CKBD0 U635 ( .CLK(n752), .C(n753) );
  CKBD0 U636 ( .CLK(n753), .C(n754) );
  CKBD0 U637 ( .CLK(n754), .C(n755) );
  CKBD0 U638 ( .CLK(n755), .C(n756) );
  BUFFD0 U639 ( .I(n756), .Z(n757) );
  CKBD0 U640 ( .CLK(n757), .C(n758) );
  CKBD0 U641 ( .CLK(n758), .C(n759) );
  CKBD0 U642 ( .CLK(n759), .C(n760) );
  CKBD0 U643 ( .CLK(n760), .C(n761) );
  CKBD0 U644 ( .CLK(n761), .C(n762) );
  BUFFD0 U645 ( .I(n8437), .Z(n763) );
  CKBD0 U646 ( .CLK(FrameSR[54]), .C(n764) );
  BUFFD0 U647 ( .I(n764), .Z(n765) );
  CKBD0 U648 ( .CLK(n765), .C(n766) );
  CKBD0 U649 ( .CLK(n766), .C(n767) );
  CKBD0 U650 ( .CLK(n767), .C(n768) );
  CKBD0 U651 ( .CLK(n768), .C(n769) );
  CKBD0 U652 ( .CLK(n769), .C(n770) );
  CKBD0 U653 ( .CLK(n770), .C(n771) );
  CKBD0 U654 ( .CLK(n771), .C(n772) );
  CKBD0 U655 ( .CLK(n772), .C(n773) );
  CKBD0 U656 ( .CLK(n773), .C(n774) );
  BUFFD0 U657 ( .I(n774), .Z(n775) );
  CKBD0 U658 ( .CLK(n775), .C(n776) );
  CKBD0 U659 ( .CLK(n776), .C(n777) );
  CKBD0 U660 ( .CLK(n777), .C(n778) );
  CKBD0 U661 ( .CLK(n778), .C(n779) );
  CKBD0 U662 ( .CLK(n779), .C(n780) );
  CKBD0 U663 ( .CLK(n780), .C(n781) );
  CKBD0 U664 ( .CLK(n781), .C(n782) );
  CKBD0 U665 ( .CLK(n782), .C(n783) );
  CKBD0 U666 ( .CLK(n783), .C(n784) );
  CKBD0 U667 ( .CLK(n784), .C(n785) );
  BUFFD0 U668 ( .I(n785), .Z(n786) );
  CKBD0 U669 ( .CLK(n786), .C(n787) );
  CKBD0 U670 ( .CLK(n787), .C(n788) );
  CKBD0 U671 ( .CLK(n788), .C(n789) );
  CKBD0 U672 ( .CLK(n789), .C(n790) );
  CKBD0 U673 ( .CLK(n790), .C(n791) );
  CKBD0 U674 ( .CLK(n791), .C(n792) );
  CKBD0 U675 ( .CLK(n792), .C(n793) );
  CKBD0 U676 ( .CLK(n793), .C(n794) );
  CKBD0 U677 ( .CLK(n794), .C(n795) );
  CKBD0 U678 ( .CLK(n795), .C(n796) );
  BUFFD0 U679 ( .I(n796), .Z(n797) );
  CKBD0 U680 ( .CLK(n797), .C(n798) );
  CKBD0 U681 ( .CLK(n798), .C(n799) );
  CKBD0 U682 ( .CLK(n799), .C(n800) );
  CKBD0 U683 ( .CLK(n800), .C(n801) );
  CKBD0 U684 ( .CLK(n801), .C(n802) );
  CKBD0 U685 ( .CLK(n802), .C(n803) );
  CKBD0 U686 ( .CLK(n803), .C(n804) );
  CKBD0 U687 ( .CLK(n804), .C(n805) );
  CKBD0 U688 ( .CLK(n805), .C(n806) );
  CKBD0 U689 ( .CLK(n806), .C(n807) );
  BUFFD0 U690 ( .I(n807), .Z(n808) );
  CKBD0 U691 ( .CLK(n808), .C(n809) );
  CKBD0 U692 ( .CLK(n809), .C(n810) );
  CKBD0 U693 ( .CLK(n810), .C(n811) );
  CKBD0 U694 ( .CLK(n811), .C(n812) );
  CKBD0 U695 ( .CLK(n812), .C(n813) );
  CKBD0 U696 ( .CLK(n813), .C(n814) );
  CKBD0 U697 ( .CLK(n814), .C(n815) );
  CKBD0 U698 ( .CLK(n815), .C(n816) );
  CKBD0 U699 ( .CLK(n816), .C(n817) );
  CKBD0 U700 ( .CLK(n817), .C(n818) );
  BUFFD0 U701 ( .I(n818), .Z(n819) );
  CKBD0 U702 ( .CLK(n819), .C(n820) );
  CKBD0 U703 ( .CLK(n820), .C(n821) );
  CKBD0 U704 ( .CLK(n821), .C(n822) );
  CKBD0 U705 ( .CLK(n822), .C(n823) );
  CKBD0 U706 ( .CLK(n823), .C(n824) );
  CKBD0 U707 ( .CLK(n824), .C(n825) );
  CKBD0 U708 ( .CLK(n825), .C(n826) );
  CKBD0 U709 ( .CLK(n826), .C(n827) );
  CKBD0 U710 ( .CLK(n827), .C(n828) );
  CKBD0 U711 ( .CLK(n828), .C(n829) );
  BUFFD0 U712 ( .I(n829), .Z(n830) );
  CKBD0 U713 ( .CLK(n830), .C(n831) );
  CKBD0 U714 ( .CLK(n831), .C(n832) );
  CKBD0 U715 ( .CLK(n832), .C(n833) );
  CKBD0 U716 ( .CLK(n833), .C(n834) );
  CKBD0 U717 ( .CLK(n834), .C(n835) );
  CKBD0 U718 ( .CLK(n835), .C(n836) );
  CKBD0 U719 ( .CLK(n836), .C(n837) );
  CKBD0 U720 ( .CLK(n837), .C(n838) );
  CKBD0 U721 ( .CLK(n838), .C(n839) );
  CKBD0 U722 ( .CLK(n839), .C(n840) );
  BUFFD0 U723 ( .I(n840), .Z(n841) );
  CKBD0 U724 ( .CLK(n841), .C(n842) );
  CKBD0 U725 ( .CLK(n842), .C(n843) );
  CKBD0 U726 ( .CLK(n843), .C(n844) );
  CKBD0 U727 ( .CLK(n844), .C(n845) );
  CKBD0 U728 ( .CLK(n845), .C(n846) );
  CKBD0 U729 ( .CLK(n846), .C(n847) );
  CKBD0 U730 ( .CLK(n847), .C(n848) );
  CKBD0 U731 ( .CLK(n848), .C(n849) );
  CKBD0 U732 ( .CLK(n849), .C(n850) );
  CKBD0 U733 ( .CLK(n850), .C(n851) );
  CKBD0 U734 ( .CLK(n851), .C(n852) );
  BUFFD0 U735 ( .I(n8897), .Z(n853) );
  CKBD0 U736 ( .CLK(FrameSR[7]), .C(n854) );
  CKBD0 U737 ( .CLK(n854), .C(n855) );
  CKBD0 U738 ( .CLK(n855), .C(n856) );
  BUFFD0 U739 ( .I(n6723), .Z(n857) );
  CKBD0 U740 ( .CLK(FrameSR[8]), .C(n858) );
  BUFFD0 U741 ( .I(n6586), .Z(n859) );
  CKBD0 U742 ( .CLK(FrameSR[9]), .C(n860) );
  BUFFD0 U743 ( .I(n6449), .Z(n861) );
  CKBD0 U744 ( .CLK(FrameSR[10]), .C(n862) );
  BUFFD0 U745 ( .I(n6312), .Z(n863) );
  CKBD0 U746 ( .CLK(FrameSR[11]), .C(n864) );
  BUFFD0 U747 ( .I(n6175), .Z(n865) );
  CKBD0 U748 ( .CLK(FrameSR[12]), .C(n866) );
  BUFFD0 U749 ( .I(n6038), .Z(n867) );
  CKBD0 U750 ( .CLK(FrameSR[13]), .C(n868) );
  BUFFD0 U751 ( .I(n5901), .Z(n869) );
  CKBD0 U752 ( .CLK(FrameSR[14]), .C(n870) );
  BUFFD0 U753 ( .I(n8550), .Z(n871) );
  CKBD0 U754 ( .CLK(FrameSR[18]), .C(n872) );
  CKBD0 U755 ( .CLK(n872), .C(n873) );
  CKBD0 U756 ( .CLK(n873), .C(n874) );
  CKBD0 U757 ( .CLK(n874), .C(n875) );
  CKBD0 U758 ( .CLK(n875), .C(n876) );
  CKBD0 U759 ( .CLK(n876), .C(n877) );
  CKBD0 U760 ( .CLK(n877), .C(n878) );
  CKBD0 U761 ( .CLK(n878), .C(n879) );
  BUFFD0 U762 ( .I(n879), .Z(n880) );
  CKBD0 U763 ( .CLK(n880), .C(n881) );
  CKBD0 U764 ( .CLK(n881), .C(n882) );
  CKBD0 U765 ( .CLK(n882), .C(n883) );
  CKBD0 U766 ( .CLK(n883), .C(n884) );
  CKBD0 U767 ( .CLK(n884), .C(n885) );
  CKBD0 U768 ( .CLK(n885), .C(n886) );
  CKBD0 U769 ( .CLK(n886), .C(n887) );
  CKBD0 U770 ( .CLK(n887), .C(n888) );
  CKBD0 U771 ( .CLK(n888), .C(n889) );
  CKBD0 U772 ( .CLK(n889), .C(n890) );
  BUFFD0 U773 ( .I(n890), .Z(n891) );
  CKBD0 U774 ( .CLK(n891), .C(n892) );
  CKBD0 U775 ( .CLK(n892), .C(n893) );
  CKBD0 U776 ( .CLK(n893), .C(n894) );
  CKBD0 U777 ( .CLK(n894), .C(n895) );
  CKBD0 U778 ( .CLK(n895), .C(n896) );
  CKBD0 U779 ( .CLK(n896), .C(n897) );
  CKBD0 U780 ( .CLK(n897), .C(n898) );
  CKBD0 U781 ( .CLK(n898), .C(n899) );
  CKBD0 U782 ( .CLK(n899), .C(n900) );
  CKBD0 U783 ( .CLK(n900), .C(n901) );
  BUFFD0 U784 ( .I(n901), .Z(n902) );
  CKBD0 U785 ( .CLK(n902), .C(n903) );
  CKBD0 U786 ( .CLK(n903), .C(n904) );
  CKBD0 U787 ( .CLK(n904), .C(n905) );
  CKBD0 U788 ( .CLK(n905), .C(n906) );
  CKBD0 U789 ( .CLK(n906), .C(n907) );
  CKBD0 U790 ( .CLK(n907), .C(n908) );
  CKBD0 U791 ( .CLK(n908), .C(n909) );
  CKBD0 U792 ( .CLK(n909), .C(n910) );
  CKBD0 U793 ( .CLK(n910), .C(n911) );
  CKBD0 U794 ( .CLK(n911), .C(n912) );
  BUFFD0 U795 ( .I(n912), .Z(n913) );
  CKBD0 U796 ( .CLK(n913), .C(n914) );
  CKBD0 U797 ( .CLK(n914), .C(n915) );
  CKBD0 U798 ( .CLK(n915), .C(n916) );
  CKBD0 U799 ( .CLK(n916), .C(n917) );
  CKBD0 U800 ( .CLK(n917), .C(n918) );
  CKBD0 U801 ( .CLK(n918), .C(n919) );
  CKBD0 U802 ( .CLK(n919), .C(n920) );
  CKBD0 U803 ( .CLK(n920), .C(n921) );
  CKBD0 U804 ( .CLK(n921), .C(n922) );
  BUFFD0 U805 ( .I(n922), .Z(n923) );
  CKBD0 U806 ( .CLK(n923), .C(n924) );
  CKBD0 U807 ( .CLK(n924), .C(n925) );
  CKBD0 U808 ( .CLK(n925), .C(n926) );
  CKBD0 U809 ( .CLK(n926), .C(n927) );
  CKBD0 U810 ( .CLK(n927), .C(n928) );
  CKBD0 U811 ( .CLK(n928), .C(n929) );
  CKBD0 U812 ( .CLK(n929), .C(n930) );
  CKBD0 U813 ( .CLK(n930), .C(n931) );
  CKBD0 U814 ( .CLK(n931), .C(n932) );
  CKBD0 U815 ( .CLK(n932), .C(n933) );
  BUFFD0 U816 ( .I(n933), .Z(n934) );
  CKBD0 U817 ( .CLK(n934), .C(n935) );
  CKBD0 U818 ( .CLK(n935), .C(n936) );
  CKBD0 U819 ( .CLK(n936), .C(n937) );
  CKBD0 U820 ( .CLK(n937), .C(n938) );
  CKBD0 U821 ( .CLK(n938), .C(n939) );
  CKBD0 U822 ( .CLK(n939), .C(n940) );
  CKBD0 U823 ( .CLK(n940), .C(n941) );
  CKBD0 U824 ( .CLK(n941), .C(n942) );
  CKBD0 U825 ( .CLK(n942), .C(n943) );
  CKBD0 U826 ( .CLK(n943), .C(n944) );
  BUFFD0 U827 ( .I(n944), .Z(n945) );
  CKBD0 U828 ( .CLK(n945), .C(n946) );
  CKBD0 U829 ( .CLK(n946), .C(n947) );
  CKBD0 U830 ( .CLK(n947), .C(n948) );
  CKBD0 U831 ( .CLK(n948), .C(n949) );
  CKBD0 U832 ( .CLK(n949), .C(n950) );
  CKBD0 U833 ( .CLK(n950), .C(n951) );
  CKBD0 U834 ( .CLK(n951), .C(n952) );
  CKBD0 U835 ( .CLK(n952), .C(n953) );
  CKBD0 U836 ( .CLK(n953), .C(n954) );
  CKBD0 U837 ( .CLK(n954), .C(n955) );
  BUFFD0 U838 ( .I(n955), .Z(n956) );
  CKBD0 U839 ( .CLK(n956), .C(n957) );
  CKBD0 U840 ( .CLK(n957), .C(n958) );
  CKBD0 U841 ( .CLK(n958), .C(n959) );
  BUFFD0 U842 ( .I(n8180), .Z(n960) );
  CKBD0 U843 ( .CLK(FrameSR[23]), .C(n961) );
  CKBD0 U844 ( .CLK(n961), .C(n962) );
  CKBD0 U845 ( .CLK(n962), .C(n963) );
  CKBD0 U846 ( .CLK(n963), .C(n964) );
  CKBD0 U847 ( .CLK(n964), .C(n965) );
  BUFFD0 U848 ( .I(n965), .Z(n966) );
  CKBD0 U849 ( .CLK(n966), .C(n967) );
  CKBD0 U850 ( .CLK(n967), .C(n968) );
  CKBD0 U851 ( .CLK(n968), .C(n969) );
  CKBD0 U852 ( .CLK(n969), .C(n970) );
  CKBD0 U853 ( .CLK(n970), .C(n971) );
  CKBD0 U854 ( .CLK(n971), .C(n972) );
  CKBD0 U855 ( .CLK(n972), .C(n973) );
  CKBD0 U856 ( .CLK(n973), .C(n974) );
  CKBD0 U857 ( .CLK(n974), .C(n975) );
  CKBD0 U858 ( .CLK(n975), .C(n976) );
  BUFFD0 U859 ( .I(n976), .Z(n977) );
  CKBD0 U860 ( .CLK(n977), .C(n978) );
  CKBD0 U861 ( .CLK(n978), .C(n979) );
  CKBD0 U862 ( .CLK(n979), .C(n980) );
  CKBD0 U863 ( .CLK(n980), .C(n981) );
  CKBD0 U864 ( .CLK(n981), .C(n982) );
  CKBD0 U865 ( .CLK(n982), .C(n983) );
  CKBD0 U866 ( .CLK(n983), .C(n984) );
  CKBD0 U867 ( .CLK(n984), .C(n985) );
  CKBD0 U868 ( .CLK(n985), .C(n986) );
  CKBD0 U869 ( .CLK(n986), .C(n987) );
  BUFFD0 U870 ( .I(n987), .Z(n988) );
  CKBD0 U871 ( .CLK(n988), .C(n989) );
  CKBD0 U872 ( .CLK(n989), .C(n990) );
  CKBD0 U873 ( .CLK(n990), .C(n991) );
  CKBD0 U874 ( .CLK(n991), .C(n992) );
  CKBD0 U875 ( .CLK(n992), .C(n993) );
  CKBD0 U876 ( .CLK(n993), .C(n994) );
  CKBD0 U877 ( .CLK(n994), .C(n995) );
  CKBD0 U878 ( .CLK(n995), .C(n996) );
  CKBD0 U879 ( .CLK(n996), .C(n997) );
  CKBD0 U880 ( .CLK(n997), .C(n998) );
  BUFFD0 U881 ( .I(n998), .Z(n999) );
  CKBD0 U882 ( .CLK(n999), .C(n1000) );
  CKBD0 U883 ( .CLK(n1000), .C(n1001) );
  CKBD0 U884 ( .CLK(n1001), .C(n1002) );
  CKBD0 U885 ( .CLK(n1002), .C(n1003) );
  CKBD0 U886 ( .CLK(n1003), .C(n1004) );
  CKBD0 U887 ( .CLK(n1004), .C(n1005) );
  CKBD0 U888 ( .CLK(n1005), .C(n1006) );
  CKBD0 U889 ( .CLK(n1006), .C(n1007) );
  CKBD0 U890 ( .CLK(n1007), .C(n1008) );
  CKBD0 U891 ( .CLK(n1008), .C(n1009) );
  BUFFD0 U892 ( .I(n1009), .Z(n1010) );
  CKBD0 U893 ( .CLK(n1010), .C(n1011) );
  CKBD0 U894 ( .CLK(n1011), .C(n1012) );
  CKBD0 U895 ( .CLK(n1012), .C(n1013) );
  CKBD0 U896 ( .CLK(n1013), .C(n1014) );
  CKBD0 U897 ( .CLK(n1014), .C(n1015) );
  CKBD0 U898 ( .CLK(n1015), .C(n1016) );
  CKBD0 U899 ( .CLK(n1016), .C(n1017) );
  CKBD0 U900 ( .CLK(n1017), .C(n1018) );
  CKBD0 U901 ( .CLK(n1018), .C(n1019) );
  BUFFD0 U902 ( .I(n1019), .Z(n1020) );
  CKBD0 U903 ( .CLK(n1020), .C(n1021) );
  CKBD0 U904 ( .CLK(n1021), .C(n1022) );
  CKBD0 U905 ( .CLK(n1022), .C(n1023) );
  CKBD0 U906 ( .CLK(n1023), .C(n1024) );
  CKBD0 U907 ( .CLK(n1024), .C(n1025) );
  CKBD0 U908 ( .CLK(n1025), .C(n1026) );
  CKBD0 U909 ( .CLK(n1026), .C(n1027) );
  CKBD0 U910 ( .CLK(n1027), .C(n1028) );
  CKBD0 U911 ( .CLK(n1028), .C(n1029) );
  CKBD0 U912 ( .CLK(n1029), .C(n1030) );
  BUFFD0 U913 ( .I(n1030), .Z(n1031) );
  CKBD0 U914 ( .CLK(n1031), .C(n1032) );
  CKBD0 U915 ( .CLK(n1032), .C(n1033) );
  CKBD0 U916 ( .CLK(n1033), .C(n1034) );
  CKBD0 U917 ( .CLK(n1034), .C(n1035) );
  CKBD0 U918 ( .CLK(n1035), .C(n1036) );
  CKBD0 U919 ( .CLK(n1036), .C(n1037) );
  CKBD0 U920 ( .CLK(n1037), .C(n1038) );
  CKBD0 U921 ( .CLK(n1038), .C(n1039) );
  CKBD0 U922 ( .CLK(n1039), .C(n1040) );
  CKBD0 U923 ( .CLK(n1040), .C(n1041) );
  BUFFD0 U924 ( .I(n1041), .Z(n1042) );
  CKBD0 U925 ( .CLK(n1042), .C(n1043) );
  CKBD0 U926 ( .CLK(n1043), .C(n1044) );
  CKBD0 U927 ( .CLK(n1044), .C(n1045) );
  CKBD0 U928 ( .CLK(n1045), .C(n1046) );
  CKBD0 U929 ( .CLK(n1046), .C(n1047) );
  CKBD0 U930 ( .CLK(n1047), .C(n1048) );
  CKBD0 U931 ( .CLK(n1048), .C(n1049) );
  BUFFD0 U932 ( .I(n5628), .Z(n1050) );
  CKBD0 U933 ( .CLK(FrameSR[24]), .C(n1051) );
  BUFFD0 U934 ( .I(n5491), .Z(n1052) );
  CKBD0 U935 ( .CLK(FrameSR[25]), .C(n1053) );
  BUFFD0 U936 ( .I(n5354), .Z(n1054) );
  CKBD0 U937 ( .CLK(FrameSR[26]), .C(n1055) );
  BUFFD0 U938 ( .I(n5218), .Z(n1056) );
  CKBD0 U939 ( .CLK(FrameSR[27]), .C(n1057) );
  BUFFD0 U940 ( .I(n5082), .Z(n1058) );
  CKBD0 U941 ( .CLK(FrameSR[28]), .C(n1059) );
  BUFFD0 U942 ( .I(n4946), .Z(n1060) );
  CKBD0 U943 ( .CLK(FrameSR[29]), .C(n1061) );
  BUFFD0 U944 ( .I(n4810), .Z(n1062) );
  CKBD0 U945 ( .CLK(FrameSR[30]), .C(n1063) );
  BUFFD0 U946 ( .I(n8342), .Z(n1064) );
  CKBD0 U947 ( .CLK(FrameSR[39]), .C(n1065) );
  CKBD0 U948 ( .CLK(n1065), .C(n1066) );
  CKBD0 U949 ( .CLK(n1066), .C(n1067) );
  CKBD0 U950 ( .CLK(n1067), .C(n1068) );
  CKBD0 U951 ( .CLK(n1068), .C(n1069) );
  CKBD0 U952 ( .CLK(n1069), .C(n1070) );
  CKBD0 U953 ( .CLK(n1070), .C(n1071) );
  BUFFD0 U954 ( .I(n1071), .Z(n1072) );
  CKBD0 U955 ( .CLK(n1072), .C(n1073) );
  CKBD0 U956 ( .CLK(n1073), .C(n1074) );
  CKBD0 U957 ( .CLK(n1074), .C(n1075) );
  CKBD0 U958 ( .CLK(n1075), .C(n1076) );
  CKBD0 U959 ( .CLK(n1076), .C(n1077) );
  CKBD0 U960 ( .CLK(n1077), .C(n1078) );
  CKBD0 U961 ( .CLK(n1078), .C(n1079) );
  CKBD0 U962 ( .CLK(n1079), .C(n1080) );
  CKBD0 U963 ( .CLK(n1080), .C(n1081) );
  CKBD0 U964 ( .CLK(n1081), .C(n1082) );
  BUFFD0 U965 ( .I(n1082), .Z(n1083) );
  CKBD0 U966 ( .CLK(n1083), .C(n1084) );
  CKBD0 U967 ( .CLK(n1084), .C(n1085) );
  CKBD0 U968 ( .CLK(n1085), .C(n1086) );
  CKBD0 U969 ( .CLK(n1086), .C(n1087) );
  CKBD0 U970 ( .CLK(n1087), .C(n1088) );
  CKBD0 U971 ( .CLK(n1088), .C(n1089) );
  CKBD0 U972 ( .CLK(n1089), .C(n1090) );
  CKBD0 U973 ( .CLK(n1090), .C(n1091) );
  CKBD0 U974 ( .CLK(n1091), .C(n1092) );
  CKBD0 U975 ( .CLK(n1092), .C(n1093) );
  BUFFD0 U976 ( .I(n1093), .Z(n1094) );
  CKBD0 U977 ( .CLK(n1094), .C(n1095) );
  CKBD0 U978 ( .CLK(n1095), .C(n1096) );
  CKBD0 U979 ( .CLK(n1096), .C(n1097) );
  CKBD0 U980 ( .CLK(n1097), .C(n1098) );
  CKBD0 U981 ( .CLK(n1098), .C(n1099) );
  CKBD0 U982 ( .CLK(n1099), .C(n1100) );
  CKBD0 U983 ( .CLK(n1100), .C(n1101) );
  CKBD0 U984 ( .CLK(n1101), .C(n1102) );
  CKBD0 U985 ( .CLK(n1102), .C(n1103) );
  BUFFD0 U986 ( .I(n1103), .Z(n1104) );
  CKBD0 U987 ( .CLK(n1104), .C(n1105) );
  CKBD0 U988 ( .CLK(n1105), .C(n1106) );
  CKBD0 U989 ( .CLK(n1106), .C(n1107) );
  CKBD0 U990 ( .CLK(n1107), .C(n1108) );
  CKBD0 U991 ( .CLK(n1108), .C(n1109) );
  CKBD0 U992 ( .CLK(n1109), .C(n1110) );
  CKBD0 U993 ( .CLK(n1110), .C(n1111) );
  CKBD0 U994 ( .CLK(n1111), .C(n1112) );
  CKBD0 U995 ( .CLK(n1112), .C(n1113) );
  CKBD0 U996 ( .CLK(n1113), .C(n1114) );
  BUFFD0 U997 ( .I(n1114), .Z(n1115) );
  CKBD0 U998 ( .CLK(n1115), .C(n1116) );
  CKBD0 U999 ( .CLK(n1116), .C(n1117) );
  CKBD0 U1000 ( .CLK(n1117), .C(n1118) );
  CKBD0 U1001 ( .CLK(n1118), .C(n1119) );
  CKBD0 U1002 ( .CLK(n1119), .C(n1120) );
  CKBD0 U1003 ( .CLK(n1120), .C(n1121) );
  CKBD0 U1004 ( .CLK(n1121), .C(n1122) );
  CKBD0 U1005 ( .CLK(n1122), .C(n1123) );
  CKBD0 U1006 ( .CLK(n1123), .C(n1124) );
  CKBD0 U1007 ( .CLK(n1124), .C(n1125) );
  BUFFD0 U1008 ( .I(n1125), .Z(n1126) );
  CKBD0 U1009 ( .CLK(n1126), .C(n1127) );
  CKBD0 U1010 ( .CLK(n1127), .C(n1128) );
  CKBD0 U1011 ( .CLK(n1128), .C(n1129) );
  CKBD0 U1012 ( .CLK(n1129), .C(n1130) );
  CKBD0 U1013 ( .CLK(n1130), .C(n1131) );
  CKBD0 U1014 ( .CLK(n1131), .C(n1132) );
  CKBD0 U1015 ( .CLK(n1132), .C(n1133) );
  CKBD0 U1016 ( .CLK(n1133), .C(n1134) );
  CKBD0 U1017 ( .CLK(n1134), .C(n1135) );
  CKBD0 U1018 ( .CLK(n1135), .C(n1136) );
  BUFFD0 U1019 ( .I(n1136), .Z(n1137) );
  CKBD0 U1020 ( .CLK(n1137), .C(n1138) );
  CKBD0 U1021 ( .CLK(n1138), .C(n1139) );
  CKBD0 U1022 ( .CLK(n1139), .C(n1140) );
  CKBD0 U1023 ( .CLK(n1140), .C(n1141) );
  CKBD0 U1024 ( .CLK(n1141), .C(n1142) );
  CKBD0 U1025 ( .CLK(n1142), .C(n1143) );
  CKBD0 U1026 ( .CLK(n1143), .C(n1144) );
  CKBD0 U1027 ( .CLK(n1144), .C(n1145) );
  CKBD0 U1028 ( .CLK(n1145), .C(n1146) );
  CKBD0 U1029 ( .CLK(n1146), .C(n1147) );
  BUFFD0 U1030 ( .I(n1147), .Z(n1148) );
  CKBD0 U1031 ( .CLK(n1148), .C(n1149) );
  CKBD0 U1032 ( .CLK(n1149), .C(n1150) );
  CKBD0 U1033 ( .CLK(n1150), .C(n1151) );
  CKBD0 U1034 ( .CLK(n1151), .C(n1152) );
  CKBD0 U1035 ( .CLK(n1152), .C(n1153) );
  BUFFD0 U1036 ( .I(n4538), .Z(n1154) );
  CKBD0 U1037 ( .CLK(FrameSR[40]), .C(n1155) );
  BUFFD0 U1038 ( .I(n4402), .Z(n1156) );
  CKBD0 U1039 ( .CLK(FrameSR[41]), .C(n1157) );
  BUFFD0 U1040 ( .I(n4266), .Z(n1158) );
  CKBD0 U1041 ( .CLK(FrameSR[42]), .C(n1159) );
  BUFFD0 U1042 ( .I(n4130), .Z(n1160) );
  CKBD0 U1043 ( .CLK(FrameSR[43]), .C(n1161) );
  BUFFD0 U1044 ( .I(n3994), .Z(n1162) );
  CKBD0 U1045 ( .CLK(FrameSR[44]), .C(n1163) );
  BUFFD0 U1046 ( .I(n3858), .Z(n1164) );
  CKBD0 U1047 ( .CLK(FrameSR[45]), .C(n1165) );
  BUFFD0 U1048 ( .I(n3722), .Z(n1166) );
  CKBD0 U1049 ( .CLK(FrameSR[46]), .C(n1167) );
  BUFFD0 U1050 ( .I(n8214), .Z(n1168) );
  CKBD0 U1051 ( .CLK(FrameSR[55]), .C(n1169) );
  CKBD0 U1052 ( .CLK(n1169), .C(n1170) );
  CKBD0 U1053 ( .CLK(n1170), .C(n1171) );
  CKBD0 U1054 ( .CLK(n1171), .C(n1172) );
  CKBD0 U1055 ( .CLK(n1172), .C(n1173) );
  CKBD0 U1056 ( .CLK(n1173), .C(n1174) );
  CKBD0 U1057 ( .CLK(n1174), .C(n1175) );
  BUFFD0 U1058 ( .I(n1175), .Z(n1176) );
  CKBD0 U1059 ( .CLK(n1176), .C(n1177) );
  CKBD0 U1060 ( .CLK(n1177), .C(n1178) );
  CKBD0 U1061 ( .CLK(n1178), .C(n1179) );
  CKBD0 U1062 ( .CLK(n1179), .C(n1180) );
  CKBD0 U1063 ( .CLK(n1180), .C(n1181) );
  CKBD0 U1064 ( .CLK(n1181), .C(n1182) );
  CKBD0 U1065 ( .CLK(n1182), .C(n1183) );
  CKBD0 U1066 ( .CLK(n1183), .C(n1184) );
  CKBD0 U1067 ( .CLK(n1184), .C(n1185) );
  CKBD0 U1068 ( .CLK(n1185), .C(n1186) );
  BUFFD0 U1069 ( .I(n1186), .Z(n1187) );
  CKBD0 U1070 ( .CLK(n1187), .C(n1188) );
  CKBD0 U1071 ( .CLK(n1188), .C(n1189) );
  CKBD0 U1072 ( .CLK(n1189), .C(n1190) );
  CKBD0 U1073 ( .CLK(n1190), .C(n1191) );
  CKBD0 U1074 ( .CLK(n1191), .C(n1192) );
  CKBD0 U1075 ( .CLK(n1192), .C(n1193) );
  CKBD0 U1076 ( .CLK(n1193), .C(n1194) );
  CKBD0 U1077 ( .CLK(n1194), .C(n1195) );
  CKBD0 U1078 ( .CLK(n1195), .C(n1196) );
  CKBD0 U1079 ( .CLK(n1196), .C(n1197) );
  BUFFD0 U1080 ( .I(n1197), .Z(n1198) );
  CKBD0 U1081 ( .CLK(n1198), .C(n1199) );
  CKBD0 U1082 ( .CLK(n1199), .C(n1200) );
  CKBD0 U1083 ( .CLK(n1200), .C(n1201) );
  CKBD0 U1084 ( .CLK(n1201), .C(n1202) );
  CKBD0 U1085 ( .CLK(n1202), .C(n1203) );
  CKBD0 U1086 ( .CLK(n1203), .C(n1204) );
  CKBD0 U1087 ( .CLK(n1204), .C(n1205) );
  CKBD0 U1088 ( .CLK(n1205), .C(n1206) );
  CKBD0 U1089 ( .CLK(n1206), .C(n1207) );
  BUFFD0 U1090 ( .I(n1207), .Z(n1208) );
  CKBD0 U1091 ( .CLK(n1208), .C(n1209) );
  CKBD0 U1092 ( .CLK(n1209), .C(n1210) );
  CKBD0 U1093 ( .CLK(n1210), .C(n1211) );
  CKBD0 U1094 ( .CLK(n1211), .C(n1212) );
  CKBD0 U1095 ( .CLK(n1212), .C(n1213) );
  CKBD0 U1096 ( .CLK(n1213), .C(n1214) );
  CKBD0 U1097 ( .CLK(n1214), .C(n1215) );
  CKBD0 U1098 ( .CLK(n1215), .C(n1216) );
  CKBD0 U1099 ( .CLK(n1216), .C(n1217) );
  CKBD0 U1100 ( .CLK(n1217), .C(n1218) );
  BUFFD0 U1101 ( .I(n1218), .Z(n1219) );
  CKBD0 U1102 ( .CLK(n1219), .C(n1220) );
  CKBD0 U1103 ( .CLK(n1220), .C(n1221) );
  CKBD0 U1104 ( .CLK(n1221), .C(n1222) );
  CKBD0 U1105 ( .CLK(n1222), .C(n1223) );
  CKBD0 U1106 ( .CLK(n1223), .C(n1224) );
  CKBD0 U1107 ( .CLK(n1224), .C(n1225) );
  CKBD0 U1108 ( .CLK(n1225), .C(n1226) );
  CKBD0 U1109 ( .CLK(n1226), .C(n1227) );
  CKBD0 U1110 ( .CLK(n1227), .C(n1228) );
  CKBD0 U1111 ( .CLK(n1228), .C(n1229) );
  BUFFD0 U1112 ( .I(n1229), .Z(n1230) );
  CKBD0 U1113 ( .CLK(n1230), .C(n1231) );
  CKBD0 U1114 ( .CLK(n1231), .C(n1232) );
  CKBD0 U1115 ( .CLK(n1232), .C(n1233) );
  CKBD0 U1116 ( .CLK(n1233), .C(n1234) );
  CKBD0 U1117 ( .CLK(n1234), .C(n1235) );
  CKBD0 U1118 ( .CLK(n1235), .C(n1236) );
  CKBD0 U1119 ( .CLK(n1236), .C(n1237) );
  CKBD0 U1120 ( .CLK(n1237), .C(n1238) );
  CKBD0 U1121 ( .CLK(n1238), .C(n1239) );
  CKBD0 U1122 ( .CLK(n1239), .C(n1240) );
  BUFFD0 U1123 ( .I(n1240), .Z(n1241) );
  CKBD0 U1124 ( .CLK(n1241), .C(n1242) );
  CKBD0 U1125 ( .CLK(n1242), .C(n1243) );
  CKBD0 U1126 ( .CLK(n1243), .C(n1244) );
  CKBD0 U1127 ( .CLK(n1244), .C(n1245) );
  CKBD0 U1128 ( .CLK(n1245), .C(n1246) );
  CKBD0 U1129 ( .CLK(n1246), .C(n1247) );
  CKBD0 U1130 ( .CLK(n1247), .C(n1248) );
  CKBD0 U1131 ( .CLK(n1248), .C(n1249) );
  CKBD0 U1132 ( .CLK(n1249), .C(n1250) );
  CKBD0 U1133 ( .CLK(n1250), .C(n1251) );
  BUFFD0 U1134 ( .I(n1251), .Z(n1252) );
  CKBD0 U1135 ( .CLK(n1252), .C(n1253) );
  CKBD0 U1136 ( .CLK(n1253), .C(n1254) );
  CKBD0 U1137 ( .CLK(n1254), .C(n1255) );
  CKBD0 U1138 ( .CLK(n1255), .C(n1256) );
  CKBD0 U1139 ( .CLK(n1256), .C(n1257) );
  BUFFD0 U1140 ( .I(n3450), .Z(n1258) );
  CKBD0 U1141 ( .CLK(FrameSR[56]), .C(n1259) );
  BUFFD0 U1142 ( .I(n3314), .Z(n1260) );
  CKBD0 U1143 ( .CLK(FrameSR[57]), .C(n1261) );
  BUFFD0 U1144 ( .I(n3178), .Z(n1262) );
  CKBD0 U1145 ( .CLK(FrameSR[58]), .C(n1263) );
  BUFFD0 U1146 ( .I(n3042), .Z(n1264) );
  CKBD0 U1147 ( .CLK(FrameSR[59]), .C(n1265) );
  BUFFD0 U1148 ( .I(n2906), .Z(n1266) );
  CKBD0 U1149 ( .CLK(FrameSR[60]), .C(n1267) );
  BUFFD0 U1150 ( .I(n2770), .Z(n1268) );
  CKBD0 U1151 ( .CLK(FrameSR[61]), .C(n1269) );
  BUFFD0 U1152 ( .I(n8916), .Z(n1270) );
  CKBD0 U1153 ( .CLK(FrameSR[3]), .C(n1271) );
  CKBD0 U1154 ( .CLK(n1271), .C(n1272) );
  BUFFD0 U1155 ( .I(n8383), .Z(n1273) );
  CKBD0 U1156 ( .CLK(FrameSR[19]), .C(n1274) );
  CKBD0 U1157 ( .CLK(n1274), .C(n1275) );
  CKBD0 U1158 ( .CLK(n1275), .C(n1276) );
  CKBD0 U1159 ( .CLK(n1276), .C(n1277) );
  BUFFD0 U1160 ( .I(n1277), .Z(n1278) );
  CKBD0 U1161 ( .CLK(n1278), .C(n1279) );
  CKBD0 U1162 ( .CLK(n1279), .C(n1280) );
  CKBD0 U1163 ( .CLK(n1280), .C(n1281) );
  CKBD0 U1164 ( .CLK(n1281), .C(n1282) );
  CKBD0 U1165 ( .CLK(n1282), .C(n1283) );
  CKBD0 U1166 ( .CLK(n1283), .C(n1284) );
  CKBD0 U1167 ( .CLK(n1284), .C(n1285) );
  CKBD0 U1168 ( .CLK(n1285), .C(n1286) );
  CKBD0 U1169 ( .CLK(n1286), .C(n1287) );
  CKBD0 U1170 ( .CLK(n1287), .C(n1288) );
  BUFFD0 U1171 ( .I(n1288), .Z(n1289) );
  CKBD0 U1172 ( .CLK(n1289), .C(n1290) );
  CKBD0 U1173 ( .CLK(n1290), .C(n1291) );
  CKBD0 U1174 ( .CLK(n1291), .C(n1292) );
  CKBD0 U1175 ( .CLK(n1292), .C(n1293) );
  CKBD0 U1176 ( .CLK(n1293), .C(n1294) );
  CKBD0 U1177 ( .CLK(n1294), .C(n1295) );
  CKBD0 U1178 ( .CLK(n1295), .C(n1296) );
  CKBD0 U1179 ( .CLK(n1296), .C(n1297) );
  CKBD0 U1180 ( .CLK(n1297), .C(n1298) );
  CKBD0 U1181 ( .CLK(n1298), .C(n1299) );
  BUFFD0 U1182 ( .I(n1299), .Z(n1300) );
  CKBD0 U1183 ( .CLK(n1300), .C(n1301) );
  CKBD0 U1184 ( .CLK(n1301), .C(n1302) );
  CKBD0 U1185 ( .CLK(n1302), .C(n1303) );
  CKBD0 U1186 ( .CLK(n1303), .C(n1304) );
  CKBD0 U1187 ( .CLK(n1304), .C(n1305) );
  CKBD0 U1188 ( .CLK(n1305), .C(n1306) );
  CKBD0 U1189 ( .CLK(n1306), .C(n1307) );
  CKBD0 U1190 ( .CLK(n1307), .C(n1308) );
  CKBD0 U1191 ( .CLK(n1308), .C(n1309) );
  CKBD0 U1192 ( .CLK(n1309), .C(n1310) );
  BUFFD0 U1193 ( .I(n1310), .Z(n1311) );
  CKBD0 U1194 ( .CLK(n1311), .C(n1312) );
  CKBD0 U1195 ( .CLK(n1312), .C(n1313) );
  CKBD0 U1196 ( .CLK(n1313), .C(n1314) );
  CKBD0 U1197 ( .CLK(n1314), .C(n1315) );
  CKBD0 U1198 ( .CLK(n1315), .C(n1316) );
  CKBD0 U1199 ( .CLK(n1316), .C(n1317) );
  CKBD0 U1200 ( .CLK(n1317), .C(n1318) );
  CKBD0 U1201 ( .CLK(n1318), .C(n1319) );
  CKBD0 U1202 ( .CLK(n1319), .C(n1320) );
  BUFFD0 U1203 ( .I(n1320), .Z(n1321) );
  CKBD0 U1204 ( .CLK(n1321), .C(n1322) );
  CKBD0 U1205 ( .CLK(n1322), .C(n1323) );
  CKBD0 U1206 ( .CLK(n1323), .C(n1324) );
  CKBD0 U1207 ( .CLK(n1324), .C(n1325) );
  CKBD0 U1208 ( .CLK(n1325), .C(n1326) );
  CKBD0 U1209 ( .CLK(n1326), .C(n1327) );
  CKBD0 U1210 ( .CLK(n1327), .C(n1328) );
  CKBD0 U1211 ( .CLK(n1328), .C(n1329) );
  CKBD0 U1212 ( .CLK(n1329), .C(n1330) );
  CKBD0 U1213 ( .CLK(n1330), .C(n1331) );
  BUFFD0 U1214 ( .I(n1331), .Z(n1332) );
  CKBD0 U1215 ( .CLK(n1332), .C(n1333) );
  CKBD0 U1216 ( .CLK(n1333), .C(n1334) );
  CKBD0 U1217 ( .CLK(n1334), .C(n1335) );
  CKBD0 U1218 ( .CLK(n1335), .C(n1336) );
  CKBD0 U1219 ( .CLK(n1336), .C(n1337) );
  CKBD0 U1220 ( .CLK(n1337), .C(n1338) );
  CKBD0 U1221 ( .CLK(n1338), .C(n1339) );
  CKBD0 U1222 ( .CLK(n1339), .C(n1340) );
  CKBD0 U1223 ( .CLK(n1340), .C(n1341) );
  CKBD0 U1224 ( .CLK(n1341), .C(n1342) );
  BUFFD0 U1225 ( .I(n1342), .Z(n1343) );
  CKBD0 U1226 ( .CLK(n1343), .C(n1344) );
  CKBD0 U1227 ( .CLK(n1344), .C(n1345) );
  CKBD0 U1228 ( .CLK(n1345), .C(n1346) );
  CKBD0 U1229 ( .CLK(n1346), .C(n1347) );
  CKBD0 U1230 ( .CLK(n1347), .C(n1348) );
  CKBD0 U1231 ( .CLK(n1348), .C(n1349) );
  CKBD0 U1232 ( .CLK(n1349), .C(n1350) );
  CKBD0 U1233 ( .CLK(n1350), .C(n1351) );
  CKBD0 U1234 ( .CLK(n1351), .C(n1352) );
  CKBD0 U1235 ( .CLK(n1352), .C(n1353) );
  BUFFD0 U1236 ( .I(n1353), .Z(n1354) );
  CKBD0 U1237 ( .CLK(n1354), .C(n1355) );
  CKBD0 U1238 ( .CLK(n1355), .C(n1356) );
  CKBD0 U1239 ( .CLK(n1356), .C(n1357) );
  CKBD0 U1240 ( .CLK(n1357), .C(n1358) );
  CKBD0 U1241 ( .CLK(n1358), .C(n1359) );
  CKBD0 U1242 ( .CLK(n1359), .C(n1360) );
  BUFFD0 U1243 ( .I(n8343), .Z(n1361) );
  CKBD0 U1244 ( .CLK(FrameSR[33]), .C(n1362) );
  CKBD0 U1245 ( .CLK(n1362), .C(n1363) );
  CKBD0 U1246 ( .CLK(n1363), .C(n1364) );
  CKBD0 U1247 ( .CLK(n1364), .C(n1365) );
  CKBD0 U1248 ( .CLK(n1365), .C(n1366) );
  CKBD0 U1249 ( .CLK(n1366), .C(n1367) );
  CKBD0 U1250 ( .CLK(n1367), .C(n1368) );
  CKBD0 U1251 ( .CLK(n1368), .C(n1369) );
  CKBD0 U1252 ( .CLK(n1369), .C(n1370) );
  CKBD0 U1253 ( .CLK(n1370), .C(n1371) );
  BUFFD0 U1254 ( .I(n1371), .Z(n1372) );
  CKBD0 U1255 ( .CLK(n1372), .C(n1373) );
  CKBD0 U1256 ( .CLK(n1373), .C(n1374) );
  CKBD0 U1257 ( .CLK(n1374), .C(n1375) );
  CKBD0 U1258 ( .CLK(n1375), .C(n1376) );
  CKBD0 U1259 ( .CLK(n1376), .C(n1377) );
  CKBD0 U1260 ( .CLK(n1377), .C(n1378) );
  CKBD0 U1261 ( .CLK(n1378), .C(n1379) );
  CKBD0 U1262 ( .CLK(n1379), .C(n1380) );
  CKBD0 U1263 ( .CLK(n1380), .C(n1381) );
  CKBD0 U1264 ( .CLK(n1381), .C(n1382) );
  BUFFD0 U1265 ( .I(n1382), .Z(n1383) );
  CKBD0 U1266 ( .CLK(n1383), .C(n1384) );
  CKBD0 U1267 ( .CLK(n1384), .C(n1385) );
  CKBD0 U1268 ( .CLK(n1385), .C(n1386) );
  CKBD0 U1269 ( .CLK(n1386), .C(n1387) );
  CKBD0 U1270 ( .CLK(n1387), .C(n1388) );
  CKBD0 U1271 ( .CLK(n1388), .C(n1389) );
  CKBD0 U1272 ( .CLK(n1389), .C(n1390) );
  CKBD0 U1273 ( .CLK(n1390), .C(n1391) );
  CKBD0 U1274 ( .CLK(n1391), .C(n1392) );
  CKBD0 U1275 ( .CLK(n1392), .C(n1393) );
  BUFFD0 U1276 ( .I(n1393), .Z(n1394) );
  CKBD0 U1277 ( .CLK(n1394), .C(n1395) );
  CKBD0 U1278 ( .CLK(n1395), .C(n1396) );
  CKBD0 U1279 ( .CLK(n1396), .C(n1397) );
  CKBD0 U1280 ( .CLK(n1397), .C(n1398) );
  CKBD0 U1281 ( .CLK(n1398), .C(n1399) );
  CKBD0 U1282 ( .CLK(n1399), .C(n1400) );
  CKBD0 U1283 ( .CLK(n1400), .C(n1401) );
  CKBD0 U1284 ( .CLK(n1401), .C(n1402) );
  CKBD0 U1285 ( .CLK(n1402), .C(n1403) );
  CKBD0 U1286 ( .CLK(n1403), .C(n1404) );
  BUFFD0 U1287 ( .I(n1404), .Z(n1405) );
  CKBD0 U1288 ( .CLK(n1405), .C(n1406) );
  CKBD0 U1289 ( .CLK(n1406), .C(n1407) );
  CKBD0 U1290 ( .CLK(n1407), .C(n1408) );
  CKBD0 U1291 ( .CLK(n1408), .C(n1409) );
  CKBD0 U1292 ( .CLK(n1409), .C(n1410) );
  CKBD0 U1293 ( .CLK(n1410), .C(n1411) );
  CKBD0 U1294 ( .CLK(n1411), .C(n1412) );
  CKBD0 U1295 ( .CLK(n1412), .C(n1413) );
  CKBD0 U1296 ( .CLK(n1413), .C(n1414) );
  CKBD0 U1297 ( .CLK(n1414), .C(n1415) );
  BUFFD0 U1298 ( .I(n1415), .Z(n1416) );
  CKBD0 U1299 ( .CLK(n1416), .C(n1417) );
  CKBD0 U1300 ( .CLK(n1417), .C(n1418) );
  CKBD0 U1301 ( .CLK(n1418), .C(n1419) );
  CKBD0 U1302 ( .CLK(n1419), .C(n1420) );
  CKBD0 U1303 ( .CLK(n1420), .C(n1421) );
  CKBD0 U1304 ( .CLK(n1421), .C(n1422) );
  CKBD0 U1305 ( .CLK(n1422), .C(n1423) );
  CKBD0 U1306 ( .CLK(n1423), .C(n1424) );
  CKBD0 U1307 ( .CLK(n1424), .C(n1425) );
  BUFFD0 U1308 ( .I(n1425), .Z(n1426) );
  CKBD0 U1309 ( .CLK(n1426), .C(n1427) );
  CKBD0 U1310 ( .CLK(n1427), .C(n1428) );
  CKBD0 U1311 ( .CLK(n1428), .C(n1429) );
  CKBD0 U1312 ( .CLK(n1429), .C(n1430) );
  CKBD0 U1313 ( .CLK(n1430), .C(n1431) );
  CKBD0 U1314 ( .CLK(n1431), .C(n1432) );
  CKBD0 U1315 ( .CLK(n1432), .C(n1433) );
  CKBD0 U1316 ( .CLK(n1433), .C(n1434) );
  CKBD0 U1317 ( .CLK(n1434), .C(n1435) );
  CKBD0 U1318 ( .CLK(n1435), .C(n1436) );
  BUFFD0 U1319 ( .I(n1436), .Z(n1437) );
  CKBD0 U1320 ( .CLK(n1437), .C(n1438) );
  CKBD0 U1321 ( .CLK(n1438), .C(n1439) );
  CKBD0 U1322 ( .CLK(n1439), .C(n1440) );
  CKBD0 U1323 ( .CLK(n1440), .C(n1441) );
  CKBD0 U1324 ( .CLK(n1441), .C(n1442) );
  CKBD0 U1325 ( .CLK(n1442), .C(n1443) );
  CKBD0 U1326 ( .CLK(n1443), .C(n1444) );
  CKBD0 U1327 ( .CLK(n1444), .C(n1445) );
  CKBD0 U1328 ( .CLK(n1445), .C(n1446) );
  CKBD0 U1329 ( .CLK(n1446), .C(n1447) );
  BUFFD0 U1330 ( .I(n1447), .Z(n1448) );
  CKBD0 U1331 ( .CLK(n1448), .C(n1449) );
  BUFFD0 U1332 ( .I(n8286), .Z(n1450) );
  CKBD0 U1333 ( .CLK(FrameSR[48]), .C(n1451) );
  CKBD0 U1334 ( .CLK(n1451), .C(n1452) );
  CKBD0 U1335 ( .CLK(n1452), .C(n1453) );
  CKBD0 U1336 ( .CLK(n1453), .C(n1454) );
  CKBD0 U1337 ( .CLK(n1454), .C(n1455) );
  CKBD0 U1338 ( .CLK(n1455), .C(n1456) );
  CKBD0 U1339 ( .CLK(n1456), .C(n1457) );
  CKBD0 U1340 ( .CLK(n1457), .C(n1458) );
  BUFFD0 U1341 ( .I(n1458), .Z(n1459) );
  CKBD0 U1342 ( .CLK(n1459), .C(n1460) );
  CKBD0 U1343 ( .CLK(n1460), .C(n1461) );
  CKBD0 U1344 ( .CLK(n1461), .C(n1462) );
  CKBD0 U1345 ( .CLK(n1462), .C(n1463) );
  CKBD0 U1346 ( .CLK(n1463), .C(n1464) );
  CKBD0 U1347 ( .CLK(n1464), .C(n1465) );
  CKBD0 U1348 ( .CLK(n1465), .C(n1466) );
  CKBD0 U1349 ( .CLK(n1466), .C(n1467) );
  CKBD0 U1350 ( .CLK(n1467), .C(n1468) );
  CKBD0 U1351 ( .CLK(n1468), .C(n1469) );
  BUFFD0 U1352 ( .I(n1469), .Z(n1470) );
  CKBD0 U1353 ( .CLK(n1470), .C(n1471) );
  CKBD0 U1354 ( .CLK(n1471), .C(n1472) );
  CKBD0 U1355 ( .CLK(n1472), .C(n1473) );
  CKBD0 U1356 ( .CLK(n1473), .C(n1474) );
  CKBD0 U1357 ( .CLK(n1474), .C(n1475) );
  CKBD0 U1358 ( .CLK(n1475), .C(n1476) );
  CKBD0 U1359 ( .CLK(n1476), .C(n1477) );
  CKBD0 U1360 ( .CLK(n1477), .C(n1478) );
  CKBD0 U1361 ( .CLK(n1478), .C(n1479) );
  CKBD0 U1362 ( .CLK(n1479), .C(n1480) );
  BUFFD0 U1363 ( .I(n1480), .Z(n1481) );
  CKBD0 U1364 ( .CLK(n1481), .C(n1482) );
  CKBD0 U1365 ( .CLK(n1482), .C(n1483) );
  CKBD0 U1366 ( .CLK(n1483), .C(n1484) );
  CKBD0 U1367 ( .CLK(n1484), .C(n1485) );
  CKBD0 U1368 ( .CLK(n1485), .C(n1486) );
  CKBD0 U1369 ( .CLK(n1486), .C(n1487) );
  CKBD0 U1370 ( .CLK(n1487), .C(n1488) );
  CKBD0 U1371 ( .CLK(n1488), .C(n1489) );
  CKBD0 U1372 ( .CLK(n1489), .C(n1490) );
  CKBD0 U1373 ( .CLK(n1490), .C(n1491) );
  BUFFD0 U1374 ( .I(n1491), .Z(n1492) );
  CKBD0 U1375 ( .CLK(n1492), .C(n1493) );
  CKBD0 U1376 ( .CLK(n1493), .C(n1494) );
  CKBD0 U1377 ( .CLK(n1494), .C(n1495) );
  CKBD0 U1378 ( .CLK(n1495), .C(n1496) );
  CKBD0 U1379 ( .CLK(n1496), .C(n1497) );
  CKBD0 U1380 ( .CLK(n1497), .C(n1498) );
  CKBD0 U1381 ( .CLK(n1498), .C(n1499) );
  CKBD0 U1382 ( .CLK(n1499), .C(n1500) );
  CKBD0 U1383 ( .CLK(n1500), .C(n1501) );
  BUFFD0 U1384 ( .I(n1501), .Z(n1502) );
  CKBD0 U1385 ( .CLK(n1502), .C(n1503) );
  CKBD0 U1386 ( .CLK(n1503), .C(n1504) );
  CKBD0 U1387 ( .CLK(n1504), .C(n1505) );
  CKBD0 U1388 ( .CLK(n1505), .C(n1506) );
  CKBD0 U1389 ( .CLK(n1506), .C(n1507) );
  CKBD0 U1390 ( .CLK(n1507), .C(n1508) );
  CKBD0 U1391 ( .CLK(n1508), .C(n1509) );
  CKBD0 U1392 ( .CLK(n1509), .C(n1510) );
  CKBD0 U1393 ( .CLK(n1510), .C(n1511) );
  CKBD0 U1394 ( .CLK(n1511), .C(n1512) );
  BUFFD0 U1395 ( .I(n1512), .Z(n1513) );
  CKBD0 U1396 ( .CLK(n1513), .C(n1514) );
  CKBD0 U1397 ( .CLK(n1514), .C(n1515) );
  CKBD0 U1398 ( .CLK(n1515), .C(n1516) );
  CKBD0 U1399 ( .CLK(n1516), .C(n1517) );
  CKBD0 U1400 ( .CLK(n1517), .C(n1518) );
  CKBD0 U1401 ( .CLK(n1518), .C(n1519) );
  CKBD0 U1402 ( .CLK(n1519), .C(n1520) );
  CKBD0 U1403 ( .CLK(n1520), .C(n1521) );
  CKBD0 U1404 ( .CLK(n1521), .C(n1522) );
  CKBD0 U1405 ( .CLK(n1522), .C(n1523) );
  BUFFD0 U1406 ( .I(n1523), .Z(n1524) );
  CKBD0 U1407 ( .CLK(n1524), .C(n1525) );
  CKBD0 U1408 ( .CLK(n1525), .C(n1526) );
  CKBD0 U1409 ( .CLK(n1526), .C(n1527) );
  CKBD0 U1410 ( .CLK(n1527), .C(n1528) );
  CKBD0 U1411 ( .CLK(n1528), .C(n1529) );
  CKBD0 U1412 ( .CLK(n1529), .C(n1530) );
  CKBD0 U1413 ( .CLK(n1530), .C(n1531) );
  CKBD0 U1414 ( .CLK(n1531), .C(n1532) );
  CKBD0 U1415 ( .CLK(n1532), .C(n1533) );
  CKBD0 U1416 ( .CLK(n1533), .C(n1534) );
  BUFFD0 U1417 ( .I(n1534), .Z(n1535) );
  CKBD0 U1418 ( .CLK(n1535), .C(n1536) );
  CKBD0 U1419 ( .CLK(n1536), .C(n1537) );
  CKBD0 U1420 ( .CLK(n1537), .C(n1538) );
  BUFFD0 U1421 ( .I(n8913), .Z(n1539) );
  CKBD0 U1422 ( .CLK(FrameSR[1]), .C(n1540) );
  CKBD0 U1423 ( .CLK(n1540), .C(n1541) );
  BUFFD0 U1424 ( .I(n8875), .Z(n1542) );
  CKBD0 U1425 ( .CLK(FrameSR[5]), .C(n1543) );
  CKBD0 U1426 ( .CLK(n1543), .C(n1544) );
  CKBD0 U1427 ( .CLK(n1544), .C(n1545) );
  BUFFD0 U1428 ( .I(n8553), .Z(n1546) );
  CKBD0 U1429 ( .CLK(FrameSR[17]), .C(n1547) );
  BUFFD0 U1430 ( .I(n1547), .Z(n1548) );
  CKBD0 U1431 ( .CLK(n1548), .C(n1549) );
  CKBD0 U1432 ( .CLK(n1549), .C(n1550) );
  CKBD0 U1433 ( .CLK(n1550), .C(n1551) );
  CKBD0 U1434 ( .CLK(n1551), .C(n1552) );
  CKBD0 U1435 ( .CLK(n1552), .C(n1553) );
  CKBD0 U1436 ( .CLK(n1553), .C(n1554) );
  CKBD0 U1437 ( .CLK(n1554), .C(n1555) );
  CKBD0 U1438 ( .CLK(n1555), .C(n1556) );
  CKBD0 U1439 ( .CLK(n1556), .C(n1557) );
  CKBD0 U1440 ( .CLK(n1557), .C(n1558) );
  BUFFD0 U1441 ( .I(n1558), .Z(n1559) );
  CKBD0 U1442 ( .CLK(n1559), .C(n1560) );
  CKBD0 U1443 ( .CLK(n1560), .C(n1561) );
  CKBD0 U1444 ( .CLK(n1561), .C(n1562) );
  CKBD0 U1445 ( .CLK(n1562), .C(n1563) );
  CKBD0 U1446 ( .CLK(n1563), .C(n1564) );
  CKBD0 U1447 ( .CLK(n1564), .C(n1565) );
  CKBD0 U1448 ( .CLK(n1565), .C(n1566) );
  CKBD0 U1449 ( .CLK(n1566), .C(n1567) );
  CKBD0 U1450 ( .CLK(n1567), .C(n1568) );
  CKBD0 U1451 ( .CLK(n1568), .C(n1569) );
  BUFFD0 U1452 ( .I(n1569), .Z(n1570) );
  CKBD0 U1453 ( .CLK(n1570), .C(n1571) );
  CKBD0 U1454 ( .CLK(n1571), .C(n1572) );
  CKBD0 U1455 ( .CLK(n1572), .C(n1573) );
  CKBD0 U1456 ( .CLK(n1573), .C(n1574) );
  CKBD0 U1457 ( .CLK(n1574), .C(n1575) );
  CKBD0 U1458 ( .CLK(n1575), .C(n1576) );
  CKBD0 U1459 ( .CLK(n1576), .C(n1577) );
  CKBD0 U1460 ( .CLK(n1577), .C(n1578) );
  CKBD0 U1461 ( .CLK(n1578), .C(n1579) );
  BUFFD0 U1462 ( .I(n1579), .Z(n1580) );
  CKBD0 U1463 ( .CLK(n1580), .C(n1581) );
  CKBD0 U1464 ( .CLK(n1581), .C(n1582) );
  CKBD0 U1465 ( .CLK(n1582), .C(n1583) );
  CKBD0 U1466 ( .CLK(n1583), .C(n1584) );
  CKBD0 U1467 ( .CLK(n1584), .C(n1585) );
  CKBD0 U1468 ( .CLK(n1585), .C(n1586) );
  CKBD0 U1469 ( .CLK(n1586), .C(n1587) );
  CKBD0 U1470 ( .CLK(n1587), .C(n1588) );
  CKBD0 U1471 ( .CLK(n1588), .C(n1589) );
  CKBD0 U1472 ( .CLK(n1589), .C(n1590) );
  BUFFD0 U1473 ( .I(n1590), .Z(n1591) );
  CKBD0 U1474 ( .CLK(n1591), .C(n1592) );
  CKBD0 U1475 ( .CLK(n1592), .C(n1593) );
  CKBD0 U1476 ( .CLK(n1593), .C(n1594) );
  CKBD0 U1477 ( .CLK(n1594), .C(n1595) );
  CKBD0 U1478 ( .CLK(n1595), .C(n1596) );
  CKBD0 U1479 ( .CLK(n1596), .C(n1597) );
  CKBD0 U1480 ( .CLK(n1597), .C(n1598) );
  CKBD0 U1481 ( .CLK(n1598), .C(n1599) );
  CKBD0 U1482 ( .CLK(n1599), .C(n1600) );
  CKBD0 U1483 ( .CLK(n1600), .C(n1601) );
  BUFFD0 U1484 ( .I(n1601), .Z(n1602) );
  CKBD0 U1485 ( .CLK(n1602), .C(n1603) );
  CKBD0 U1486 ( .CLK(n1603), .C(n1604) );
  CKBD0 U1487 ( .CLK(n1604), .C(n1605) );
  CKBD0 U1488 ( .CLK(n1605), .C(n1606) );
  CKBD0 U1489 ( .CLK(n1606), .C(n1607) );
  CKBD0 U1490 ( .CLK(n1607), .C(n1608) );
  CKBD0 U1491 ( .CLK(n1608), .C(n1609) );
  CKBD0 U1492 ( .CLK(n1609), .C(n1610) );
  CKBD0 U1493 ( .CLK(n1610), .C(n1611) );
  CKBD0 U1494 ( .CLK(n1611), .C(n1612) );
  BUFFD0 U1495 ( .I(n1612), .Z(n1613) );
  CKBD0 U1496 ( .CLK(n1613), .C(n1614) );
  CKBD0 U1497 ( .CLK(n1614), .C(n1615) );
  CKBD0 U1498 ( .CLK(n1615), .C(n1616) );
  CKBD0 U1499 ( .CLK(n1616), .C(n1617) );
  CKBD0 U1500 ( .CLK(n1617), .C(n1618) );
  CKBD0 U1501 ( .CLK(n1618), .C(n1619) );
  CKBD0 U1502 ( .CLK(n1619), .C(n1620) );
  CKBD0 U1503 ( .CLK(n1620), .C(n1621) );
  CKBD0 U1504 ( .CLK(n1621), .C(n1622) );
  CKBD0 U1505 ( .CLK(n1622), .C(n1623) );
  BUFFD0 U1506 ( .I(n1623), .Z(n1624) );
  CKBD0 U1507 ( .CLK(n1624), .C(n1625) );
  CKBD0 U1508 ( .CLK(n1625), .C(n1626) );
  CKBD0 U1509 ( .CLK(n1626), .C(n1627) );
  CKBD0 U1510 ( .CLK(n1627), .C(n1628) );
  CKBD0 U1511 ( .CLK(n1628), .C(n1629) );
  CKBD0 U1512 ( .CLK(n1629), .C(n1630) );
  CKBD0 U1513 ( .CLK(n1630), .C(n1631) );
  CKBD0 U1514 ( .CLK(n1631), .C(n1632) );
  CKBD0 U1515 ( .CLK(n1632), .C(n1633) );
  CKBD0 U1516 ( .CLK(n1633), .C(n1634) );
  BUFFD0 U1517 ( .I(n8539), .Z(n1635) );
  CKBD0 U1518 ( .CLK(FrameSR[32]), .C(n1636) );
  CKBD0 U1519 ( .CLK(n1636), .C(n1637) );
  CKBD0 U1520 ( .CLK(n1637), .C(n1638) );
  CKBD0 U1521 ( .CLK(n1638), .C(n1639) );
  CKBD0 U1522 ( .CLK(n1639), .C(n1640) );
  CKBD0 U1523 ( .CLK(n1640), .C(n1641) );
  CKBD0 U1524 ( .CLK(n1641), .C(n1642) );
  CKBD0 U1525 ( .CLK(n1642), .C(n1643) );
  CKBD0 U1526 ( .CLK(n1643), .C(n1644) );
  BUFFD0 U1527 ( .I(n1644), .Z(n1645) );
  CKBD0 U1528 ( .CLK(n1645), .C(n1646) );
  CKBD0 U1529 ( .CLK(n1646), .C(n1647) );
  CKBD0 U1530 ( .CLK(n1647), .C(n1648) );
  CKBD0 U1531 ( .CLK(n1648), .C(n1649) );
  CKBD0 U1532 ( .CLK(n1649), .C(n1650) );
  CKBD0 U1533 ( .CLK(n1650), .C(n1651) );
  CKBD0 U1534 ( .CLK(n1651), .C(n1652) );
  CKBD0 U1535 ( .CLK(n1652), .C(n1653) );
  CKBD0 U1536 ( .CLK(n1653), .C(n1654) );
  CKBD0 U1537 ( .CLK(n1654), .C(n1655) );
  BUFFD0 U1538 ( .I(n1655), .Z(n1656) );
  CKBD0 U1539 ( .CLK(n1656), .C(n1657) );
  CKBD0 U1540 ( .CLK(n1657), .C(n1658) );
  CKBD0 U1541 ( .CLK(n1658), .C(n1659) );
  CKBD0 U1542 ( .CLK(n1659), .C(n1660) );
  CKBD0 U1543 ( .CLK(n1660), .C(n1661) );
  CKBD0 U1544 ( .CLK(n1661), .C(n1662) );
  CKBD0 U1545 ( .CLK(n1662), .C(n1663) );
  CKBD0 U1546 ( .CLK(n1663), .C(n1664) );
  CKBD0 U1547 ( .CLK(n1664), .C(n1665) );
  CKBD0 U1548 ( .CLK(n1665), .C(n1666) );
  BUFFD0 U1549 ( .I(n1666), .Z(n1667) );
  CKBD0 U1550 ( .CLK(n1667), .C(n1668) );
  CKBD0 U1551 ( .CLK(n1668), .C(n1669) );
  CKBD0 U1552 ( .CLK(n1669), .C(n1670) );
  CKBD0 U1553 ( .CLK(n1670), .C(n1671) );
  CKBD0 U1554 ( .CLK(n1671), .C(n1672) );
  CKBD0 U1555 ( .CLK(n1672), .C(n1673) );
  CKBD0 U1556 ( .CLK(n1673), .C(n1674) );
  CKBD0 U1557 ( .CLK(n1674), .C(n1675) );
  CKBD0 U1558 ( .CLK(n1675), .C(n1676) );
  CKBD0 U1559 ( .CLK(n1676), .C(n1677) );
  BUFFD0 U1560 ( .I(n1677), .Z(n1678) );
  CKBD0 U1561 ( .CLK(n1678), .C(n1679) );
  CKBD0 U1562 ( .CLK(n1679), .C(n1680) );
  CKBD0 U1563 ( .CLK(n1680), .C(n1681) );
  CKBD0 U1564 ( .CLK(n1681), .C(n1682) );
  CKBD0 U1565 ( .CLK(n1682), .C(n1683) );
  CKBD0 U1566 ( .CLK(n1683), .C(n1684) );
  CKBD0 U1567 ( .CLK(n1684), .C(n1685) );
  CKBD0 U1568 ( .CLK(n1685), .C(n1686) );
  CKBD0 U1569 ( .CLK(n1686), .C(n1687) );
  BUFFD0 U1570 ( .I(n1687), .Z(n1688) );
  CKBD0 U1571 ( .CLK(n1688), .C(n1689) );
  CKBD0 U1572 ( .CLK(n1689), .C(n1690) );
  CKBD0 U1573 ( .CLK(n1690), .C(n1691) );
  CKBD0 U1574 ( .CLK(n1691), .C(n1692) );
  CKBD0 U1575 ( .CLK(n1692), .C(n1693) );
  CKBD0 U1576 ( .CLK(n1693), .C(n1694) );
  CKBD0 U1577 ( .CLK(n1694), .C(n1695) );
  CKBD0 U1578 ( .CLK(n1695), .C(n1696) );
  CKBD0 U1579 ( .CLK(n1696), .C(n1697) );
  CKBD0 U1580 ( .CLK(n1697), .C(n1698) );
  BUFFD0 U1581 ( .I(n1698), .Z(n1699) );
  CKBD0 U1582 ( .CLK(n1699), .C(n1700) );
  CKBD0 U1583 ( .CLK(n1700), .C(n1701) );
  CKBD0 U1584 ( .CLK(n1701), .C(n1702) );
  CKBD0 U1585 ( .CLK(n1702), .C(n1703) );
  CKBD0 U1586 ( .CLK(n1703), .C(n1704) );
  CKBD0 U1587 ( .CLK(n1704), .C(n1705) );
  CKBD0 U1588 ( .CLK(n1705), .C(n1706) );
  CKBD0 U1589 ( .CLK(n1706), .C(n1707) );
  CKBD0 U1590 ( .CLK(n1707), .C(n1708) );
  CKBD0 U1591 ( .CLK(n1708), .C(n1709) );
  BUFFD0 U1592 ( .I(n1709), .Z(n1710) );
  CKBD0 U1593 ( .CLK(n1710), .C(n1711) );
  CKBD0 U1594 ( .CLK(n1711), .C(n1712) );
  CKBD0 U1595 ( .CLK(n1712), .C(n1713) );
  CKBD0 U1596 ( .CLK(n1713), .C(n1714) );
  CKBD0 U1597 ( .CLK(n1714), .C(n1715) );
  CKBD0 U1598 ( .CLK(n1715), .C(n1716) );
  CKBD0 U1599 ( .CLK(n1716), .C(n1717) );
  CKBD0 U1600 ( .CLK(n1717), .C(n1718) );
  CKBD0 U1601 ( .CLK(n1718), .C(n1719) );
  CKBD0 U1602 ( .CLK(n1719), .C(n1720) );
  BUFFD0 U1603 ( .I(n1720), .Z(n1721) );
  CKBD0 U1604 ( .CLK(n1721), .C(n1722) );
  CKBD0 U1605 ( .CLK(n1722), .C(n1723) );
  CKBD0 U1606 ( .CLK(n1723), .C(n1724) );
  BUFFD0 U1607 ( .I(n3586), .Z(n1725) );
  CKBD0 U1608 ( .CLK(FrameSR[47]), .C(n1726) );
  BUFFD0 U1609 ( .I(n8910), .Z(n1727) );
  CKBD0 U1610 ( .CLK(FrameSR[0]), .C(n1728) );
  CKBD0 U1611 ( .CLK(n1728), .C(n1729) );
  BUFFD0 U1612 ( .I(n8906), .Z(n1730) );
  CKBD0 U1613 ( .CLK(FrameSR[2]), .C(n1731) );
  CKBD0 U1614 ( .CLK(n1731), .C(n1732) );
  BUFFD0 U1615 ( .I(n8919), .Z(n1733) );
  CKBD0 U1616 ( .CLK(FrameSR[4]), .C(n1734) );
  CKBD0 U1617 ( .CLK(n1734), .C(n1735) );
  BUFFD0 U1618 ( .I(n8882), .Z(n1736) );
  CKBD0 U1619 ( .CLK(FrameSR[6]), .C(n1737) );
  CKBD0 U1620 ( .CLK(n1737), .C(n1738) );
  CKBD0 U1621 ( .CLK(n1738), .C(n1739) );
  BUFFD0 U1622 ( .I(n8530), .Z(n1740) );
  CKBD0 U1623 ( .CLK(FrameSR[20]), .C(n1741) );
  CKBD0 U1624 ( .CLK(n1741), .C(n1742) );
  CKBD0 U1625 ( .CLK(n1742), .C(n1743) );
  CKBD0 U1626 ( .CLK(n1743), .C(n1744) );
  CKBD0 U1627 ( .CLK(n1744), .C(n1745) );
  CKBD0 U1628 ( .CLK(n1745), .C(n1746) );
  CKBD0 U1629 ( .CLK(n1746), .C(n1747) );
  CKBD0 U1630 ( .CLK(n1747), .C(n1748) );
  BUFFD0 U1631 ( .I(n1748), .Z(n1749) );
  CKBD0 U1632 ( .CLK(n1749), .C(n1750) );
  CKBD0 U1633 ( .CLK(n1750), .C(n1751) );
  CKBD0 U1634 ( .CLK(n1751), .C(n1752) );
  CKBD0 U1635 ( .CLK(n1752), .C(n1753) );
  CKBD0 U1636 ( .CLK(n1753), .C(n1754) );
  CKBD0 U1637 ( .CLK(n1754), .C(n1755) );
  CKBD0 U1638 ( .CLK(n1755), .C(n1756) );
  CKBD0 U1639 ( .CLK(n1756), .C(n1757) );
  CKBD0 U1640 ( .CLK(n1757), .C(n1758) );
  CKBD0 U1641 ( .CLK(n1758), .C(n1759) );
  BUFFD0 U1642 ( .I(n1759), .Z(n1760) );
  CKBD0 U1643 ( .CLK(n1760), .C(n1761) );
  CKBD0 U1644 ( .CLK(n1761), .C(n1762) );
  CKBD0 U1645 ( .CLK(n1762), .C(n1763) );
  CKBD0 U1646 ( .CLK(n1763), .C(n1764) );
  CKBD0 U1647 ( .CLK(n1764), .C(n1765) );
  CKBD0 U1648 ( .CLK(n1765), .C(n1766) );
  CKBD0 U1649 ( .CLK(n1766), .C(n1767) );
  CKBD0 U1650 ( .CLK(n1767), .C(n1768) );
  CKBD0 U1651 ( .CLK(n1768), .C(n1769) );
  CKBD0 U1652 ( .CLK(n1769), .C(n1770) );
  BUFFD0 U1653 ( .I(n1770), .Z(n1771) );
  CKBD0 U1654 ( .CLK(n1771), .C(n1772) );
  CKBD0 U1655 ( .CLK(n1772), .C(n1773) );
  CKBD0 U1656 ( .CLK(n1773), .C(n1774) );
  CKBD0 U1657 ( .CLK(n1774), .C(n1775) );
  CKBD0 U1658 ( .CLK(n1775), .C(n1776) );
  CKBD0 U1659 ( .CLK(n1776), .C(n1777) );
  CKBD0 U1660 ( .CLK(n1777), .C(n1778) );
  CKBD0 U1661 ( .CLK(n1778), .C(n1779) );
  CKBD0 U1662 ( .CLK(n1779), .C(n1780) );
  CKBD0 U1663 ( .CLK(n1780), .C(n1781) );
  BUFFD0 U1664 ( .I(n1781), .Z(n1782) );
  CKBD0 U1665 ( .CLK(n1782), .C(n1783) );
  CKBD0 U1666 ( .CLK(n1783), .C(n1784) );
  CKBD0 U1667 ( .CLK(n1784), .C(n1785) );
  CKBD0 U1668 ( .CLK(n1785), .C(n1786) );
  CKBD0 U1669 ( .CLK(n1786), .C(n1787) );
  CKBD0 U1670 ( .CLK(n1787), .C(n1788) );
  CKBD0 U1671 ( .CLK(n1788), .C(n1789) );
  CKBD0 U1672 ( .CLK(n1789), .C(n1790) );
  CKBD0 U1673 ( .CLK(n1790), .C(n1791) );
  BUFFD0 U1674 ( .I(n1791), .Z(n1792) );
  CKBD0 U1675 ( .CLK(n1792), .C(n1793) );
  CKBD0 U1676 ( .CLK(n1793), .C(n1794) );
  CKBD0 U1677 ( .CLK(n1794), .C(n1795) );
  CKBD0 U1678 ( .CLK(n1795), .C(n1796) );
  CKBD0 U1679 ( .CLK(n1796), .C(n1797) );
  CKBD0 U1680 ( .CLK(n1797), .C(n1798) );
  CKBD0 U1681 ( .CLK(n1798), .C(n1799) );
  CKBD0 U1682 ( .CLK(n1799), .C(n1800) );
  CKBD0 U1683 ( .CLK(n1800), .C(n1801) );
  CKBD0 U1684 ( .CLK(n1801), .C(n1802) );
  BUFFD0 U1685 ( .I(n1802), .Z(n1803) );
  CKBD0 U1686 ( .CLK(n1803), .C(n1804) );
  CKBD0 U1687 ( .CLK(n1804), .C(n1805) );
  CKBD0 U1688 ( .CLK(n1805), .C(n1806) );
  CKBD0 U1689 ( .CLK(n1806), .C(n1807) );
  CKBD0 U1690 ( .CLK(n1807), .C(n1808) );
  CKBD0 U1691 ( .CLK(n1808), .C(n1809) );
  CKBD0 U1692 ( .CLK(n1809), .C(n1810) );
  CKBD0 U1693 ( .CLK(n1810), .C(n1811) );
  CKBD0 U1694 ( .CLK(n1811), .C(n1812) );
  CKBD0 U1695 ( .CLK(n1812), .C(n1813) );
  BUFFD0 U1696 ( .I(n1813), .Z(n1814) );
  CKBD0 U1697 ( .CLK(n1814), .C(n1815) );
  CKBD0 U1698 ( .CLK(n1815), .C(n1816) );
  CKBD0 U1699 ( .CLK(n1816), .C(n1817) );
  CKBD0 U1700 ( .CLK(n1817), .C(n1818) );
  CKBD0 U1701 ( .CLK(n1818), .C(n1819) );
  CKBD0 U1702 ( .CLK(n1819), .C(n1820) );
  CKBD0 U1703 ( .CLK(n1820), .C(n1821) );
  CKBD0 U1704 ( .CLK(n1821), .C(n1822) );
  CKBD0 U1705 ( .CLK(n1822), .C(n1823) );
  CKBD0 U1706 ( .CLK(n1823), .C(n1824) );
  BUFFD0 U1707 ( .I(n1824), .Z(n1825) );
  CKBD0 U1708 ( .CLK(n1825), .C(n1826) );
  CKBD0 U1709 ( .CLK(n1826), .C(n1827) );
  CKBD0 U1710 ( .CLK(n1827), .C(n1828) );
  BUFFD0 U1711 ( .I(n8420), .Z(n1829) );
  CKBD0 U1712 ( .CLK(FrameSR[34]), .C(n1830) );
  CKBD0 U1713 ( .CLK(n1830), .C(n1831) );
  CKBD0 U1714 ( .CLK(n1831), .C(n1832) );
  CKBD0 U1715 ( .CLK(n1832), .C(n1833) );
  CKBD0 U1716 ( .CLK(n1833), .C(n1834) );
  CKBD0 U1717 ( .CLK(n1834), .C(n1835) );
  BUFFD0 U1718 ( .I(n1835), .Z(n1836) );
  CKBD0 U1719 ( .CLK(n1836), .C(n1837) );
  CKBD0 U1720 ( .CLK(n1837), .C(n1838) );
  CKBD0 U1721 ( .CLK(n1838), .C(n1839) );
  CKBD0 U1722 ( .CLK(n1839), .C(n1840) );
  CKBD0 U1723 ( .CLK(n1840), .C(n1841) );
  CKBD0 U1724 ( .CLK(n1841), .C(n1842) );
  CKBD0 U1725 ( .CLK(n1842), .C(n1843) );
  CKBD0 U1726 ( .CLK(n1843), .C(n1844) );
  CKBD0 U1727 ( .CLK(n1844), .C(n1845) );
  CKBD0 U1728 ( .CLK(n1845), .C(n1846) );
  BUFFD0 U1729 ( .I(n1846), .Z(n1847) );
  CKBD0 U1730 ( .CLK(n1847), .C(n1848) );
  CKBD0 U1731 ( .CLK(n1848), .C(n1849) );
  CKBD0 U1732 ( .CLK(n1849), .C(n1850) );
  CKBD0 U1733 ( .CLK(n1850), .C(n1851) );
  CKBD0 U1734 ( .CLK(n1851), .C(n1852) );
  CKBD0 U1735 ( .CLK(n1852), .C(n1853) );
  CKBD0 U1736 ( .CLK(n1853), .C(n1854) );
  CKBD0 U1737 ( .CLK(n1854), .C(n1855) );
  CKBD0 U1738 ( .CLK(n1855), .C(n1856) );
  CKBD0 U1739 ( .CLK(n1856), .C(n1857) );
  BUFFD0 U1740 ( .I(n1857), .Z(n1858) );
  CKBD0 U1741 ( .CLK(n1858), .C(n1859) );
  CKBD0 U1742 ( .CLK(n1859), .C(n1860) );
  CKBD0 U1743 ( .CLK(n1860), .C(n1861) );
  CKBD0 U1744 ( .CLK(n1861), .C(n1862) );
  CKBD0 U1745 ( .CLK(n1862), .C(n1863) );
  CKBD0 U1746 ( .CLK(n1863), .C(n1864) );
  CKBD0 U1747 ( .CLK(n1864), .C(n1865) );
  CKBD0 U1748 ( .CLK(n1865), .C(n1866) );
  CKBD0 U1749 ( .CLK(n1866), .C(n1867) );
  CKBD0 U1750 ( .CLK(n1867), .C(n1868) );
  BUFFD0 U1751 ( .I(n1868), .Z(n1869) );
  CKBD0 U1752 ( .CLK(n1869), .C(n1870) );
  CKBD0 U1753 ( .CLK(n1870), .C(n1871) );
  CKBD0 U1754 ( .CLK(n1871), .C(n1872) );
  CKBD0 U1755 ( .CLK(n1872), .C(n1873) );
  CKBD0 U1756 ( .CLK(n1873), .C(n1874) );
  CKBD0 U1757 ( .CLK(n1874), .C(n1875) );
  CKBD0 U1758 ( .CLK(n1875), .C(n1876) );
  CKBD0 U1759 ( .CLK(n1876), .C(n1877) );
  CKBD0 U1760 ( .CLK(n1877), .C(n1878) );
  BUFFD0 U1761 ( .I(n1878), .Z(n1879) );
  CKBD0 U1762 ( .CLK(n1879), .C(n1880) );
  CKBD0 U1763 ( .CLK(n1880), .C(n1881) );
  CKBD0 U1764 ( .CLK(n1881), .C(n1882) );
  CKBD0 U1765 ( .CLK(n1882), .C(n1883) );
  CKBD0 U1766 ( .CLK(n1883), .C(n1884) );
  CKBD0 U1767 ( .CLK(n1884), .C(n1885) );
  CKBD0 U1768 ( .CLK(n1885), .C(n1886) );
  CKBD0 U1769 ( .CLK(n1886), .C(n1887) );
  CKBD0 U1770 ( .CLK(n1887), .C(n1888) );
  CKBD0 U1771 ( .CLK(n1888), .C(n1889) );
  BUFFD0 U1772 ( .I(n1889), .Z(n1890) );
  CKBD0 U1773 ( .CLK(n1890), .C(n1891) );
  CKBD0 U1774 ( .CLK(n1891), .C(n1892) );
  CKBD0 U1775 ( .CLK(n1892), .C(n1893) );
  CKBD0 U1776 ( .CLK(n1893), .C(n1894) );
  CKBD0 U1777 ( .CLK(n1894), .C(n1895) );
  CKBD0 U1778 ( .CLK(n1895), .C(n1896) );
  CKBD0 U1779 ( .CLK(n1896), .C(n1897) );
  CKBD0 U1780 ( .CLK(n1897), .C(n1898) );
  CKBD0 U1781 ( .CLK(n1898), .C(n1899) );
  CKBD0 U1782 ( .CLK(n1899), .C(n1900) );
  BUFFD0 U1783 ( .I(n1900), .Z(n1901) );
  CKBD0 U1784 ( .CLK(n1901), .C(n1902) );
  CKBD0 U1785 ( .CLK(n1902), .C(n1903) );
  CKBD0 U1786 ( .CLK(n1903), .C(n1904) );
  CKBD0 U1787 ( .CLK(n1904), .C(n1905) );
  CKBD0 U1788 ( .CLK(n1905), .C(n1906) );
  CKBD0 U1789 ( .CLK(n1906), .C(n1907) );
  CKBD0 U1790 ( .CLK(n1907), .C(n1908) );
  CKBD0 U1791 ( .CLK(n1908), .C(n1909) );
  CKBD0 U1792 ( .CLK(n1909), .C(n1910) );
  CKBD0 U1793 ( .CLK(n1910), .C(n1911) );
  BUFFD0 U1794 ( .I(n1911), .Z(n1912) );
  CKBD0 U1795 ( .CLK(n1912), .C(n1913) );
  CKBD0 U1796 ( .CLK(n1913), .C(n1914) );
  CKBD0 U1797 ( .CLK(n1914), .C(n1915) );
  CKBD0 U1798 ( .CLK(n1915), .C(n1916) );
  CKBD0 U1799 ( .CLK(n1916), .C(n1917) );
  BUFFD0 U1800 ( .I(n8333), .Z(n1918) );
  CKBD0 U1801 ( .CLK(FrameSR[49]), .C(n1919) );
  CKBD0 U1802 ( .CLK(n1919), .C(n1920) );
  CKBD0 U1803 ( .CLK(n1920), .C(n1921) );
  CKBD0 U1804 ( .CLK(n1921), .C(n1922) );
  CKBD0 U1805 ( .CLK(n1922), .C(n1923) );
  CKBD0 U1806 ( .CLK(n1923), .C(n1924) );
  CKBD0 U1807 ( .CLK(n1924), .C(n1925) );
  CKBD0 U1808 ( .CLK(n1925), .C(n1926) );
  CKBD0 U1809 ( .CLK(n1926), .C(n1927) );
  CKBD0 U1810 ( .CLK(n1927), .C(n1928) );
  BUFFD0 U1811 ( .I(n1928), .Z(n1929) );
  CKBD0 U1812 ( .CLK(n1929), .C(n1930) );
  CKBD0 U1813 ( .CLK(n1930), .C(n1931) );
  CKBD0 U1814 ( .CLK(n1931), .C(n1932) );
  CKBD0 U1815 ( .CLK(n1932), .C(n1933) );
  CKBD0 U1816 ( .CLK(n1933), .C(n1934) );
  CKBD0 U1817 ( .CLK(n1934), .C(n1935) );
  CKBD0 U1818 ( .CLK(n1935), .C(n1936) );
  CKBD0 U1819 ( .CLK(n1936), .C(n1937) );
  CKBD0 U1820 ( .CLK(n1937), .C(n1938) );
  CKBD0 U1821 ( .CLK(n1938), .C(n1939) );
  BUFFD0 U1822 ( .I(n1939), .Z(n1940) );
  CKBD0 U1823 ( .CLK(n1940), .C(n1941) );
  CKBD0 U1824 ( .CLK(n1941), .C(n1942) );
  CKBD0 U1825 ( .CLK(n1942), .C(n1943) );
  CKBD0 U1826 ( .CLK(n1943), .C(n1944) );
  CKBD0 U1827 ( .CLK(n1944), .C(n1945) );
  CKBD0 U1828 ( .CLK(n1945), .C(n1946) );
  CKBD0 U1829 ( .CLK(n1946), .C(n1947) );
  CKBD0 U1830 ( .CLK(n1947), .C(n1948) );
  CKBD0 U1831 ( .CLK(n1948), .C(n1949) );
  CKBD0 U1832 ( .CLK(n1949), .C(n1950) );
  BUFFD0 U1833 ( .I(n1950), .Z(n1951) );
  CKBD0 U1834 ( .CLK(n1951), .C(n1952) );
  CKBD0 U1835 ( .CLK(n1952), .C(n1953) );
  CKBD0 U1836 ( .CLK(n1953), .C(n1954) );
  CKBD0 U1837 ( .CLK(n1954), .C(n1955) );
  CKBD0 U1838 ( .CLK(n1955), .C(n1956) );
  CKBD0 U1839 ( .CLK(n1956), .C(n1957) );
  CKBD0 U1840 ( .CLK(n1957), .C(n1958) );
  CKBD0 U1841 ( .CLK(n1958), .C(n1959) );
  CKBD0 U1842 ( .CLK(n1959), .C(n1960) );
  CKBD0 U1843 ( .CLK(n1960), .C(n1961) );
  BUFFD0 U1844 ( .I(n1961), .Z(n1962) );
  CKBD0 U1845 ( .CLK(n1962), .C(n1963) );
  CKBD0 U1846 ( .CLK(n1963), .C(n1964) );
  CKBD0 U1847 ( .CLK(n1964), .C(n1965) );
  CKBD0 U1848 ( .CLK(n1965), .C(n1966) );
  CKBD0 U1849 ( .CLK(n1966), .C(n1967) );
  CKBD0 U1850 ( .CLK(n1967), .C(n1968) );
  CKBD0 U1851 ( .CLK(n1968), .C(n1969) );
  CKBD0 U1852 ( .CLK(n1969), .C(n1970) );
  CKBD0 U1853 ( .CLK(n1970), .C(n1971) );
  CKBD0 U1854 ( .CLK(n1971), .C(n1972) );
  BUFFD0 U1855 ( .I(n1972), .Z(n1973) );
  CKBD0 U1856 ( .CLK(n1973), .C(n1974) );
  CKBD0 U1857 ( .CLK(n1974), .C(n1975) );
  CKBD0 U1858 ( .CLK(n1975), .C(n1976) );
  CKBD0 U1859 ( .CLK(n1976), .C(n1977) );
  CKBD0 U1860 ( .CLK(n1977), .C(n1978) );
  CKBD0 U1861 ( .CLK(n1978), .C(n1979) );
  CKBD0 U1862 ( .CLK(n1979), .C(n1980) );
  CKBD0 U1863 ( .CLK(n1980), .C(n1981) );
  CKBD0 U1864 ( .CLK(n1981), .C(n1982) );
  BUFFD0 U1865 ( .I(n1982), .Z(n1983) );
  CKBD0 U1866 ( .CLK(n1983), .C(n1984) );
  CKBD0 U1867 ( .CLK(n1984), .C(n1985) );
  CKBD0 U1868 ( .CLK(n1985), .C(n1986) );
  CKBD0 U1869 ( .CLK(n1986), .C(n1987) );
  CKBD0 U1870 ( .CLK(n1987), .C(n1988) );
  CKBD0 U1871 ( .CLK(n1988), .C(n1989) );
  CKBD0 U1872 ( .CLK(n1989), .C(n1990) );
  CKBD0 U1873 ( .CLK(n1990), .C(n1991) );
  CKBD0 U1874 ( .CLK(n1991), .C(n1992) );
  CKBD0 U1875 ( .CLK(n1992), .C(n1993) );
  BUFFD0 U1876 ( .I(n1993), .Z(n1994) );
  CKBD0 U1877 ( .CLK(n1994), .C(n1995) );
  CKBD0 U1878 ( .CLK(n1995), .C(n1996) );
  CKBD0 U1879 ( .CLK(n1996), .C(n1997) );
  CKBD0 U1880 ( .CLK(n1997), .C(n1998) );
  CKBD0 U1881 ( .CLK(n1998), .C(n1999) );
  CKBD0 U1882 ( .CLK(n1999), .C(n2000) );
  CKBD0 U1883 ( .CLK(n2000), .C(n2001) );
  CKBD0 U1884 ( .CLK(n2001), .C(n2002) );
  CKBD0 U1885 ( .CLK(n2002), .C(n2003) );
  CKBD0 U1886 ( .CLK(n2003), .C(n2004) );
  BUFFD0 U1887 ( .I(n2004), .Z(n2005) );
  CKBD0 U1888 ( .CLK(n2005), .C(n2006) );
  BUFFD0 U1889 ( .I(n8275), .Z(n2007) );
  CKBD0 U1890 ( .CLK(FrameSR[50]), .C(n2008) );
  CKBD0 U1891 ( .CLK(n2008), .C(n2009) );
  CKBD0 U1892 ( .CLK(n2009), .C(n2010) );
  CKBD0 U1893 ( .CLK(n2010), .C(n2011) );
  CKBD0 U1894 ( .CLK(n2011), .C(n2012) );
  CKBD0 U1895 ( .CLK(n2012), .C(n2013) );
  CKBD0 U1896 ( .CLK(n2013), .C(n2014) );
  CKBD0 U1897 ( .CLK(n2014), .C(n2015) );
  BUFFD0 U1898 ( .I(n2015), .Z(n2016) );
  CKBD0 U1899 ( .CLK(n2016), .C(n2017) );
  CKBD0 U1900 ( .CLK(n2017), .C(n2018) );
  CKBD0 U1901 ( .CLK(n2018), .C(n2019) );
  CKBD0 U1902 ( .CLK(n2019), .C(n2020) );
  CKBD0 U1903 ( .CLK(n2020), .C(n2021) );
  CKBD0 U1904 ( .CLK(n2021), .C(n2022) );
  CKBD0 U1905 ( .CLK(n2022), .C(n2023) );
  CKBD0 U1906 ( .CLK(n2023), .C(n2024) );
  CKBD0 U1907 ( .CLK(n2024), .C(n2025) );
  CKBD0 U1908 ( .CLK(n2025), .C(n2026) );
  BUFFD0 U1909 ( .I(n2026), .Z(n2027) );
  CKBD0 U1910 ( .CLK(n2027), .C(n2028) );
  CKBD0 U1911 ( .CLK(n2028), .C(n2029) );
  CKBD0 U1912 ( .CLK(n2029), .C(n2030) );
  CKBD0 U1913 ( .CLK(n2030), .C(n2031) );
  CKBD0 U1914 ( .CLK(n2031), .C(n2032) );
  CKBD0 U1915 ( .CLK(n2032), .C(n2033) );
  CKBD0 U1916 ( .CLK(n2033), .C(n2034) );
  CKBD0 U1917 ( .CLK(n2034), .C(n2035) );
  CKBD0 U1918 ( .CLK(n2035), .C(n2036) );
  CKBD0 U1919 ( .CLK(n2036), .C(n2037) );
  BUFFD0 U1920 ( .I(n2037), .Z(n2038) );
  CKBD0 U1921 ( .CLK(n2038), .C(n2039) );
  CKBD0 U1922 ( .CLK(n2039), .C(n2040) );
  CKBD0 U1923 ( .CLK(n2040), .C(n2041) );
  CKBD0 U1924 ( .CLK(n2041), .C(n2042) );
  CKBD0 U1925 ( .CLK(n2042), .C(n2043) );
  CKBD0 U1926 ( .CLK(n2043), .C(n2044) );
  CKBD0 U1927 ( .CLK(n2044), .C(n2045) );
  CKBD0 U1928 ( .CLK(n2045), .C(n2046) );
  CKBD0 U1929 ( .CLK(n2046), .C(n2047) );
  CKBD0 U1930 ( .CLK(n2047), .C(n2048) );
  BUFFD0 U1931 ( .I(n2048), .Z(n2049) );
  CKBD0 U1932 ( .CLK(n2049), .C(n2050) );
  CKBD0 U1933 ( .CLK(n2050), .C(n2051) );
  CKBD0 U1934 ( .CLK(n2051), .C(n2052) );
  CKBD0 U1935 ( .CLK(n2052), .C(n2053) );
  CKBD0 U1936 ( .CLK(n2053), .C(n2054) );
  CKBD0 U1937 ( .CLK(n2054), .C(n2055) );
  CKBD0 U1938 ( .CLK(n2055), .C(n2056) );
  CKBD0 U1939 ( .CLK(n2056), .C(n2057) );
  CKBD0 U1940 ( .CLK(n2057), .C(n2058) );
  BUFFD0 U1941 ( .I(n2058), .Z(n2059) );
  CKBD0 U1942 ( .CLK(n2059), .C(n2060) );
  CKBD0 U1943 ( .CLK(n2060), .C(n2061) );
  CKBD0 U1944 ( .CLK(n2061), .C(n2062) );
  CKBD0 U1945 ( .CLK(n2062), .C(n2063) );
  CKBD0 U1946 ( .CLK(n2063), .C(n2064) );
  CKBD0 U1947 ( .CLK(n2064), .C(n2065) );
  CKBD0 U1948 ( .CLK(n2065), .C(n2066) );
  CKBD0 U1949 ( .CLK(n2066), .C(n2067) );
  CKBD0 U1950 ( .CLK(n2067), .C(n2068) );
  CKBD0 U1951 ( .CLK(n2068), .C(n2069) );
  BUFFD0 U1952 ( .I(n2069), .Z(n2070) );
  CKBD0 U1953 ( .CLK(n2070), .C(n2071) );
  CKBD0 U1954 ( .CLK(n2071), .C(n2072) );
  CKBD0 U1955 ( .CLK(n2072), .C(n2073) );
  CKBD0 U1956 ( .CLK(n2073), .C(n2074) );
  CKBD0 U1957 ( .CLK(n2074), .C(n2075) );
  CKBD0 U1958 ( .CLK(n2075), .C(n2076) );
  CKBD0 U1959 ( .CLK(n2076), .C(n2077) );
  CKBD0 U1960 ( .CLK(n2077), .C(n2078) );
  CKBD0 U1961 ( .CLK(n2078), .C(n2079) );
  CKBD0 U1962 ( .CLK(n2079), .C(n2080) );
  BUFFD0 U1963 ( .I(n2080), .Z(n2081) );
  CKBD0 U1964 ( .CLK(n2081), .C(n2082) );
  CKBD0 U1965 ( .CLK(n2082), .C(n2083) );
  CKBD0 U1966 ( .CLK(n2083), .C(n2084) );
  CKBD0 U1967 ( .CLK(n2084), .C(n2085) );
  CKBD0 U1968 ( .CLK(n2085), .C(n2086) );
  CKBD0 U1969 ( .CLK(n2086), .C(n2087) );
  CKBD0 U1970 ( .CLK(n2087), .C(n2088) );
  CKBD0 U1971 ( .CLK(n2088), .C(n2089) );
  CKBD0 U1972 ( .CLK(n2089), .C(n2090) );
  CKBD0 U1973 ( .CLK(n2090), .C(n2091) );
  BUFFD0 U1974 ( .I(n2091), .Z(n2092) );
  CKBD0 U1975 ( .CLK(n2092), .C(n2093) );
  CKBD0 U1976 ( .CLK(n2093), .C(n2094) );
  CKBD0 U1977 ( .CLK(n2094), .C(n2095) );
  BUFFD0 U1978 ( .I(n8215), .Z(n2096) );
  CKBD0 U1979 ( .CLK(FrameSR[35]), .C(n2097) );
  CKBD0 U1980 ( .CLK(n2097), .C(n2098) );
  CKBD0 U1981 ( .CLK(n2098), .C(n2099) );
  CKBD0 U1982 ( .CLK(n2099), .C(n2100) );
  CKBD0 U1983 ( .CLK(n2100), .C(n2101) );
  CKBD0 U1984 ( .CLK(n2101), .C(n2102) );
  BUFFD0 U1985 ( .I(n2102), .Z(n2103) );
  CKBD0 U1986 ( .CLK(n2103), .C(n2104) );
  CKBD0 U1987 ( .CLK(n2104), .C(n2105) );
  CKBD0 U1988 ( .CLK(n2105), .C(n2106) );
  CKBD0 U1989 ( .CLK(n2106), .C(n2107) );
  CKBD0 U1990 ( .CLK(n2107), .C(n2108) );
  CKBD0 U1991 ( .CLK(n2108), .C(n2109) );
  CKBD0 U1992 ( .CLK(n2109), .C(n2110) );
  CKBD0 U1993 ( .CLK(n2110), .C(n2111) );
  CKBD0 U1994 ( .CLK(n2111), .C(n2112) );
  CKBD0 U1995 ( .CLK(n2112), .C(n2113) );
  BUFFD0 U1996 ( .I(n2113), .Z(n2114) );
  CKBD0 U1997 ( .CLK(n2114), .C(n2115) );
  CKBD0 U1998 ( .CLK(n2115), .C(n2116) );
  CKBD0 U1999 ( .CLK(n2116), .C(n2117) );
  CKBD0 U2000 ( .CLK(n2117), .C(n2118) );
  CKBD0 U2001 ( .CLK(n2118), .C(n2119) );
  CKBD0 U2002 ( .CLK(n2119), .C(n2120) );
  CKBD0 U2003 ( .CLK(n2120), .C(n2121) );
  CKBD0 U2004 ( .CLK(n2121), .C(n2122) );
  CKBD0 U2005 ( .CLK(n2122), .C(n2123) );
  CKBD0 U2006 ( .CLK(n2123), .C(n2124) );
  BUFFD0 U2007 ( .I(n2124), .Z(n2125) );
  CKBD0 U2008 ( .CLK(n2125), .C(n2126) );
  CKBD0 U2009 ( .CLK(n2126), .C(n2127) );
  CKBD0 U2010 ( .CLK(n2127), .C(n2128) );
  CKBD0 U2011 ( .CLK(n2128), .C(n2129) );
  CKBD0 U2012 ( .CLK(n2129), .C(n2130) );
  CKBD0 U2013 ( .CLK(n2130), .C(n2131) );
  CKBD0 U2014 ( .CLK(n2131), .C(n2132) );
  CKBD0 U2015 ( .CLK(n2132), .C(n2133) );
  CKBD0 U2016 ( .CLK(n2133), .C(n2134) );
  CKBD0 U2017 ( .CLK(n2134), .C(n2135) );
  BUFFD0 U2018 ( .I(n2135), .Z(n2136) );
  CKBD0 U2019 ( .CLK(n2136), .C(n2137) );
  CKBD0 U2020 ( .CLK(n2137), .C(n2138) );
  CKBD0 U2021 ( .CLK(n2138), .C(n2139) );
  CKBD0 U2022 ( .CLK(n2139), .C(n2140) );
  CKBD0 U2023 ( .CLK(n2140), .C(n2141) );
  CKBD0 U2024 ( .CLK(n2141), .C(n2142) );
  CKBD0 U2025 ( .CLK(n2142), .C(n2143) );
  CKBD0 U2026 ( .CLK(n2143), .C(n2144) );
  CKBD0 U2027 ( .CLK(n2144), .C(n2145) );
  BUFFD0 U2028 ( .I(n2145), .Z(n2146) );
  CKBD0 U2029 ( .CLK(n2146), .C(n2147) );
  CKBD0 U2030 ( .CLK(n2147), .C(n2148) );
  CKBD0 U2031 ( .CLK(n2148), .C(n2149) );
  CKBD0 U2032 ( .CLK(n2149), .C(n2150) );
  CKBD0 U2033 ( .CLK(n2150), .C(n2151) );
  CKBD0 U2034 ( .CLK(n2151), .C(n2152) );
  CKBD0 U2035 ( .CLK(n2152), .C(n2153) );
  CKBD0 U2036 ( .CLK(n2153), .C(n2154) );
  CKBD0 U2037 ( .CLK(n2154), .C(n2155) );
  CKBD0 U2038 ( .CLK(n2155), .C(n2156) );
  BUFFD0 U2039 ( .I(n2156), .Z(n2157) );
  CKBD0 U2040 ( .CLK(n2157), .C(n2158) );
  CKBD0 U2041 ( .CLK(n2158), .C(n2159) );
  CKBD0 U2042 ( .CLK(n2159), .C(n2160) );
  CKBD0 U2043 ( .CLK(n2160), .C(n2161) );
  CKBD0 U2044 ( .CLK(n2161), .C(n2162) );
  CKBD0 U2045 ( .CLK(n2162), .C(n2163) );
  CKBD0 U2046 ( .CLK(n2163), .C(n2164) );
  CKBD0 U2047 ( .CLK(n2164), .C(n2165) );
  CKBD0 U2048 ( .CLK(n2165), .C(n2166) );
  CKBD0 U2049 ( .CLK(n2166), .C(n2167) );
  BUFFD0 U2050 ( .I(n2167), .Z(n2168) );
  CKBD0 U2051 ( .CLK(n2168), .C(n2169) );
  CKBD0 U2052 ( .CLK(n2169), .C(n2170) );
  CKBD0 U2053 ( .CLK(n2170), .C(n2171) );
  CKBD0 U2054 ( .CLK(n2171), .C(n2172) );
  CKBD0 U2055 ( .CLK(n2172), .C(n2173) );
  CKBD0 U2056 ( .CLK(n2173), .C(n2174) );
  CKBD0 U2057 ( .CLK(n2174), .C(n2175) );
  CKBD0 U2058 ( .CLK(n2175), .C(n2176) );
  CKBD0 U2059 ( .CLK(n2176), .C(n2177) );
  CKBD0 U2060 ( .CLK(n2177), .C(n2178) );
  BUFFD0 U2061 ( .I(n2178), .Z(n2179) );
  CKBD0 U2062 ( .CLK(n2179), .C(n2180) );
  CKBD0 U2063 ( .CLK(n2180), .C(n2181) );
  CKBD0 U2064 ( .CLK(n2181), .C(n2182) );
  CKBD0 U2065 ( .CLK(n2182), .C(n2183) );
  CKBD0 U2066 ( .CLK(n2183), .C(n2184) );
  BUFFD0 U2067 ( .I(n8518), .Z(n2185) );
  CKBD0 U2068 ( .CLK(FrameSR[51]), .C(n2186) );
  CKBD0 U2069 ( .CLK(n2186), .C(n2187) );
  CKBD0 U2070 ( .CLK(n2187), .C(n2188) );
  CKBD0 U2071 ( .CLK(n2188), .C(n2189) );
  CKBD0 U2072 ( .CLK(n2189), .C(n2190) );
  CKBD0 U2073 ( .CLK(n2190), .C(n2191) );
  CKBD0 U2074 ( .CLK(n2191), .C(n2192) );
  BUFFD0 U2075 ( .I(n2192), .Z(n2193) );
  CKBD0 U2076 ( .CLK(n2193), .C(n2194) );
  CKBD0 U2077 ( .CLK(n2194), .C(n2195) );
  CKBD0 U2078 ( .CLK(n2195), .C(n2196) );
  CKBD0 U2079 ( .CLK(n2196), .C(n2197) );
  CKBD0 U2080 ( .CLK(n2197), .C(n2198) );
  CKBD0 U2081 ( .CLK(n2198), .C(n2199) );
  CKBD0 U2082 ( .CLK(n2199), .C(n2200) );
  CKBD0 U2083 ( .CLK(n2200), .C(n2201) );
  CKBD0 U2084 ( .CLK(n2201), .C(n2202) );
  CKBD0 U2085 ( .CLK(n2202), .C(n2203) );
  BUFFD0 U2086 ( .I(n2203), .Z(n2204) );
  CKBD0 U2087 ( .CLK(n2204), .C(n2205) );
  CKBD0 U2088 ( .CLK(n2205), .C(n2206) );
  CKBD0 U2089 ( .CLK(n2206), .C(n2207) );
  CKBD0 U2090 ( .CLK(n2207), .C(n2208) );
  CKBD0 U2091 ( .CLK(n2208), .C(n2209) );
  CKBD0 U2092 ( .CLK(n2209), .C(n2210) );
  CKBD0 U2093 ( .CLK(n2210), .C(n2211) );
  CKBD0 U2094 ( .CLK(n2211), .C(n2212) );
  CKBD0 U2095 ( .CLK(n2212), .C(n2213) );
  CKBD0 U2096 ( .CLK(n2213), .C(n2214) );
  BUFFD0 U2097 ( .I(n2214), .Z(n2215) );
  CKBD0 U2098 ( .CLK(n2215), .C(n2216) );
  CKBD0 U2099 ( .CLK(n2216), .C(n2217) );
  CKBD0 U2100 ( .CLK(n2217), .C(n2218) );
  CKBD0 U2101 ( .CLK(n2218), .C(n2219) );
  CKBD0 U2102 ( .CLK(n2219), .C(n2220) );
  CKBD0 U2103 ( .CLK(n2220), .C(n2221) );
  CKBD0 U2104 ( .CLK(n2221), .C(n2222) );
  CKBD0 U2105 ( .CLK(n2222), .C(n2223) );
  CKBD0 U2106 ( .CLK(n2223), .C(n2224) );
  CKBD0 U2107 ( .CLK(n2224), .C(n2225) );
  BUFFD0 U2108 ( .I(n2225), .Z(n2226) );
  CKBD0 U2109 ( .CLK(n2226), .C(n2227) );
  CKBD0 U2110 ( .CLK(n2227), .C(n2228) );
  CKBD0 U2111 ( .CLK(n2228), .C(n2229) );
  CKBD0 U2112 ( .CLK(n2229), .C(n2230) );
  CKBD0 U2113 ( .CLK(n2230), .C(n2231) );
  CKBD0 U2114 ( .CLK(n2231), .C(n2232) );
  CKBD0 U2115 ( .CLK(n2232), .C(n2233) );
  CKBD0 U2116 ( .CLK(n2233), .C(n2234) );
  CKBD0 U2117 ( .CLK(n2234), .C(n2235) );
  BUFFD0 U2118 ( .I(n2235), .Z(n2236) );
  CKBD0 U2119 ( .CLK(n2236), .C(n2237) );
  CKBD0 U2120 ( .CLK(n2237), .C(n2238) );
  CKBD0 U2121 ( .CLK(n2238), .C(n2239) );
  CKBD0 U2122 ( .CLK(n2239), .C(n2240) );
  CKBD0 U2123 ( .CLK(n2240), .C(n2241) );
  CKBD0 U2124 ( .CLK(n2241), .C(n2242) );
  CKBD0 U2125 ( .CLK(n2242), .C(n2243) );
  CKBD0 U2126 ( .CLK(n2243), .C(n2244) );
  CKBD0 U2127 ( .CLK(n2244), .C(n2245) );
  CKBD0 U2128 ( .CLK(n2245), .C(n2246) );
  BUFFD0 U2129 ( .I(n2246), .Z(n2247) );
  CKBD0 U2130 ( .CLK(n2247), .C(n2248) );
  CKBD0 U2131 ( .CLK(n2248), .C(n2249) );
  CKBD0 U2132 ( .CLK(n2249), .C(n2250) );
  CKBD0 U2133 ( .CLK(n2250), .C(n2251) );
  CKBD0 U2134 ( .CLK(n2251), .C(n2252) );
  CKBD0 U2135 ( .CLK(n2252), .C(n2253) );
  CKBD0 U2136 ( .CLK(n2253), .C(n2254) );
  CKBD0 U2137 ( .CLK(n2254), .C(n2255) );
  CKBD0 U2138 ( .CLK(n2255), .C(n2256) );
  CKBD0 U2139 ( .CLK(n2256), .C(n2257) );
  BUFFD0 U2140 ( .I(n2257), .Z(n2258) );
  CKBD0 U2141 ( .CLK(n2258), .C(n2259) );
  CKBD0 U2142 ( .CLK(n2259), .C(n2260) );
  CKBD0 U2143 ( .CLK(n2260), .C(n2261) );
  CKBD0 U2144 ( .CLK(n2261), .C(n2262) );
  CKBD0 U2145 ( .CLK(n2262), .C(n2263) );
  CKBD0 U2146 ( .CLK(n2263), .C(n2264) );
  CKBD0 U2147 ( .CLK(n2264), .C(n2265) );
  CKBD0 U2148 ( .CLK(n2265), .C(n2266) );
  CKBD0 U2149 ( .CLK(n2266), .C(n2267) );
  CKBD0 U2150 ( .CLK(n2267), .C(n2268) );
  BUFFD0 U2151 ( .I(n2268), .Z(n2269) );
  CKBD0 U2152 ( .CLK(n2269), .C(n2270) );
  CKBD0 U2153 ( .CLK(n2270), .C(n2271) );
  CKBD0 U2154 ( .CLK(n2271), .C(n2272) );
  BUFFD0 U2155 ( .I(n8846), .Z(n2273) );
  CKBD0 U2156 ( .CLK(FrameSR[16]), .C(n2274) );
  CKBD0 U2157 ( .CLK(n2274), .C(n2275) );
  CKBD0 U2158 ( .CLK(n2275), .C(n2276) );
  BUFFD0 U2159 ( .I(n2276), .Z(n2277) );
  CKBD0 U2160 ( .CLK(n2277), .C(n2278) );
  CKBD0 U2161 ( .CLK(n2278), .C(n2279) );
  CKBD0 U2162 ( .CLK(n2279), .C(n2280) );
  CKBD0 U2163 ( .CLK(n2280), .C(n2281) );
  CKBD0 U2164 ( .CLK(n2281), .C(n2282) );
  CKBD0 U2165 ( .CLK(n2282), .C(n2283) );
  CKBD0 U2166 ( .CLK(n2283), .C(n2284) );
  CKBD0 U2167 ( .CLK(n2284), .C(n2285) );
  CKBD0 U2168 ( .CLK(n2285), .C(n2286) );
  CKBD0 U2169 ( .CLK(n2286), .C(n2287) );
  BUFFD0 U2170 ( .I(n2287), .Z(n2288) );
  CKBD0 U2171 ( .CLK(n2288), .C(n2289) );
  CKBD0 U2172 ( .CLK(n2289), .C(n2290) );
  CKBD0 U2173 ( .CLK(n2290), .C(n2291) );
  CKBD0 U2174 ( .CLK(n2291), .C(n2292) );
  CKBD0 U2175 ( .CLK(n2292), .C(n2293) );
  CKBD0 U2176 ( .CLK(n2293), .C(n2294) );
  CKBD0 U2177 ( .CLK(n2294), .C(n2295) );
  CKBD0 U2178 ( .CLK(n2295), .C(n2296) );
  CKBD0 U2179 ( .CLK(n2296), .C(n2297) );
  CKBD0 U2180 ( .CLK(n2297), .C(n2298) );
  BUFFD0 U2181 ( .I(n2298), .Z(n2299) );
  CKBD0 U2182 ( .CLK(n2299), .C(n2300) );
  CKBD0 U2183 ( .CLK(n2300), .C(n2301) );
  CKBD0 U2184 ( .CLK(n2301), .C(n2302) );
  CKBD0 U2185 ( .CLK(n2302), .C(n2303) );
  CKBD0 U2186 ( .CLK(n2303), .C(n2304) );
  CKBD0 U2187 ( .CLK(n2304), .C(n2305) );
  CKBD0 U2188 ( .CLK(n2305), .C(n2306) );
  CKBD0 U2189 ( .CLK(n2306), .C(n2307) );
  CKBD0 U2190 ( .CLK(n2307), .C(n2308) );
  CKBD0 U2191 ( .CLK(n2308), .C(n2309) );
  BUFFD0 U2192 ( .I(n2309), .Z(n2310) );
  CKBD0 U2193 ( .CLK(n2310), .C(n2311) );
  CKBD0 U2194 ( .CLK(n2311), .C(n2312) );
  CKBD0 U2195 ( .CLK(n2312), .C(n2313) );
  CKBD0 U2196 ( .CLK(n2313), .C(n2314) );
  CKBD0 U2197 ( .CLK(n2314), .C(n2315) );
  CKBD0 U2198 ( .CLK(n2315), .C(n2316) );
  CKBD0 U2199 ( .CLK(n2316), .C(n2317) );
  CKBD0 U2200 ( .CLK(n2317), .C(n2318) );
  CKBD0 U2201 ( .CLK(n2318), .C(n2319) );
  CKBD0 U2202 ( .CLK(n2319), .C(n2320) );
  BUFFD0 U2203 ( .I(n2320), .Z(n2321) );
  CKBD0 U2204 ( .CLK(n2321), .C(n2322) );
  CKBD0 U2205 ( .CLK(n2322), .C(n2323) );
  CKBD0 U2206 ( .CLK(n2323), .C(n2324) );
  CKBD0 U2207 ( .CLK(n2324), .C(n2325) );
  CKBD0 U2208 ( .CLK(n2325), .C(n2326) );
  CKBD0 U2209 ( .CLK(n2326), .C(n2327) );
  CKBD0 U2210 ( .CLK(n2327), .C(n2328) );
  CKBD0 U2211 ( .CLK(n2328), .C(n2329) );
  CKBD0 U2212 ( .CLK(n2329), .C(n2330) );
  BUFFD0 U2213 ( .I(n2330), .Z(n2331) );
  CKBD0 U2214 ( .CLK(n2331), .C(n2332) );
  CKBD0 U2215 ( .CLK(n2332), .C(n2333) );
  CKBD0 U2216 ( .CLK(n2333), .C(n2334) );
  CKBD0 U2217 ( .CLK(n2334), .C(n2335) );
  CKBD0 U2218 ( .CLK(n2335), .C(n2336) );
  CKBD0 U2219 ( .CLK(n2336), .C(n2337) );
  CKBD0 U2220 ( .CLK(n2337), .C(n2338) );
  CKBD0 U2221 ( .CLK(n2338), .C(n2339) );
  CKBD0 U2222 ( .CLK(n2339), .C(n2340) );
  CKBD0 U2223 ( .CLK(n2340), .C(n2341) );
  BUFFD0 U2224 ( .I(n2341), .Z(n2342) );
  CKBD0 U2225 ( .CLK(n2342), .C(n2343) );
  CKBD0 U2226 ( .CLK(n2343), .C(n2344) );
  CKBD0 U2227 ( .CLK(n2344), .C(n2345) );
  CKBD0 U2228 ( .CLK(n2345), .C(n2346) );
  CKBD0 U2229 ( .CLK(n2346), .C(n2347) );
  CKBD0 U2230 ( .CLK(n2347), .C(n2348) );
  CKBD0 U2231 ( .CLK(n2348), .C(n2349) );
  CKBD0 U2232 ( .CLK(n2349), .C(n2350) );
  CKBD0 U2233 ( .CLK(n2350), .C(n2351) );
  CKBD0 U2234 ( .CLK(n2351), .C(n2352) );
  BUFFD0 U2235 ( .I(n2352), .Z(n2353) );
  CKBD0 U2236 ( .CLK(n2353), .C(n2354) );
  CKBD0 U2237 ( .CLK(n2354), .C(n2355) );
  CKBD0 U2238 ( .CLK(n2355), .C(n2356) );
  CKBD0 U2239 ( .CLK(n2356), .C(n2357) );
  CKBD0 U2240 ( .CLK(n2357), .C(n2358) );
  CKBD0 U2241 ( .CLK(n2358), .C(n2359) );
  CKBD0 U2242 ( .CLK(n2359), .C(n2360) );
  CKBD0 U2243 ( .CLK(n2360), .C(n2361) );
  BUFFD0 U2244 ( .I(n5764), .Z(n2362) );
  CKBD0 U2245 ( .CLK(FrameSR[15]), .C(n2363) );
  BUFFD0 U2246 ( .I(N42), .Z(n2364) );
  BUFFD0 U2247 ( .I(n2496), .Z(n2365) );
  CKBD0 U2248 ( .CLK(FrameSR[63]), .C(n2366) );
  CKBD0 U2249 ( .CLK(n2366), .C(n2367) );
  CKBD0 U2250 ( .CLK(n2367), .C(n2368) );
  CKBD0 U2251 ( .CLK(n2368), .C(n2369) );
  CKBD0 U2252 ( .CLK(n2369), .C(n2370) );
  CKBD0 U2253 ( .CLK(n2370), .C(n2371) );
  CKBD0 U2254 ( .CLK(n2371), .C(n2372) );
  CKBD0 U2255 ( .CLK(n2372), .C(n2373) );
  CKBD0 U2256 ( .CLK(n2373), .C(n2374) );
  CKBD0 U2257 ( .CLK(n2374), .C(n2375) );
  BUFFD0 U2258 ( .I(n2375), .Z(n2376) );
  CKBD0 U2259 ( .CLK(n2376), .C(n2377) );
  CKBD0 U2260 ( .CLK(n2377), .C(n2378) );
  CKBD0 U2261 ( .CLK(n2378), .C(n2379) );
  CKBD0 U2262 ( .CLK(n2379), .C(n2380) );
  CKBD0 U2263 ( .CLK(n2380), .C(n2381) );
  CKBD0 U2264 ( .CLK(n2381), .C(n2382) );
  CKBD0 U2265 ( .CLK(n2382), .C(n2383) );
  CKBD0 U2266 ( .CLK(n2383), .C(n2384) );
  CKBD0 U2267 ( .CLK(n2384), .C(n2385) );
  CKBD0 U2268 ( .CLK(n2385), .C(n2386) );
  BUFFD0 U2269 ( .I(n2386), .Z(n2387) );
  CKBD0 U2270 ( .CLK(n2387), .C(n2388) );
  CKBD0 U2271 ( .CLK(n2388), .C(n2389) );
  CKBD0 U2272 ( .CLK(n2389), .C(n2390) );
  CKBD0 U2273 ( .CLK(n2390), .C(n2391) );
  CKBD0 U2274 ( .CLK(n2391), .C(n2392) );
  CKBD0 U2275 ( .CLK(n2392), .C(n2393) );
  CKBD0 U2276 ( .CLK(n2393), .C(n2394) );
  CKBD0 U2277 ( .CLK(n2394), .C(n2395) );
  CKBD0 U2278 ( .CLK(n2395), .C(n2396) );
  CKBD0 U2279 ( .CLK(n2396), .C(n2397) );
  BUFFD0 U2280 ( .I(n2397), .Z(n2398) );
  CKBD0 U2281 ( .CLK(n2398), .C(n2399) );
  CKBD0 U2282 ( .CLK(n2399), .C(n2400) );
  CKBD0 U2283 ( .CLK(n2400), .C(n2401) );
  CKBD0 U2284 ( .CLK(n2401), .C(n2402) );
  CKBD0 U2285 ( .CLK(n2402), .C(n2403) );
  CKBD0 U2286 ( .CLK(n2403), .C(n2404) );
  CKBD0 U2287 ( .CLK(n2404), .C(n2405) );
  CKBD0 U2288 ( .CLK(n2405), .C(n2406) );
  CKBD0 U2289 ( .CLK(n2406), .C(n2407) );
  CKBD0 U2290 ( .CLK(n2407), .C(n2408) );
  BUFFD0 U2291 ( .I(n2408), .Z(n2409) );
  CKBD0 U2292 ( .CLK(n2409), .C(n2410) );
  CKBD0 U2293 ( .CLK(n2410), .C(n2411) );
  CKBD0 U2294 ( .CLK(n2411), .C(n2412) );
  CKBD0 U2295 ( .CLK(n2412), .C(n2413) );
  CKBD0 U2296 ( .CLK(n2413), .C(n2414) );
  CKBD0 U2297 ( .CLK(n2414), .C(n2415) );
  CKBD0 U2298 ( .CLK(n2415), .C(n2416) );
  CKBD0 U2299 ( .CLK(n2416), .C(n2417) );
  CKBD0 U2300 ( .CLK(n2417), .C(n2418) );
  CKBD0 U2301 ( .CLK(n2418), .C(n2419) );
  BUFFD0 U2302 ( .I(n2419), .Z(n2420) );
  CKBD0 U2303 ( .CLK(n2420), .C(n2421) );
  CKBD0 U2304 ( .CLK(n2421), .C(n2422) );
  CKBD0 U2305 ( .CLK(n2422), .C(n2423) );
  CKBD0 U2306 ( .CLK(n2423), .C(n2424) );
  CKBD0 U2307 ( .CLK(n2424), .C(n2425) );
  CKBD0 U2308 ( .CLK(n2425), .C(n2426) );
  CKBD0 U2309 ( .CLK(n2426), .C(n2427) );
  CKBD0 U2310 ( .CLK(n2427), .C(n2428) );
  CKBD0 U2311 ( .CLK(n2428), .C(n2429) );
  CKBD0 U2312 ( .CLK(n2429), .C(n2430) );
  BUFFD0 U2313 ( .I(n2430), .Z(n2431) );
  CKBD0 U2314 ( .CLK(n2431), .C(n2432) );
  CKBD0 U2315 ( .CLK(n2432), .C(n2433) );
  CKBD0 U2316 ( .CLK(n2433), .C(n2434) );
  CKBD0 U2317 ( .CLK(n2434), .C(n2435) );
  CKBD0 U2318 ( .CLK(n2435), .C(n2436) );
  CKBD0 U2319 ( .CLK(n2436), .C(n2437) );
  CKBD0 U2320 ( .CLK(n2437), .C(n2438) );
  CKBD0 U2321 ( .CLK(n2438), .C(n2439) );
  CKBD0 U2322 ( .CLK(n2439), .C(n2440) );
  BUFFD0 U2323 ( .I(n2440), .Z(n2441) );
  CKBD0 U2324 ( .CLK(n2441), .C(n2442) );
  CKBD0 U2325 ( .CLK(n2442), .C(n2443) );
  CKBD0 U2326 ( .CLK(n2443), .C(n2444) );
  CKBD0 U2327 ( .CLK(n2444), .C(n2445) );
  CKBD0 U2328 ( .CLK(n2445), .C(n2446) );
  CKBD0 U2329 ( .CLK(n2446), .C(n2447) );
  CKBD0 U2330 ( .CLK(n2447), .C(n2448) );
  CKBD0 U2331 ( .CLK(n2448), .C(n2449) );
  CKBD0 U2332 ( .CLK(n2449), .C(n2450) );
  CKBD0 U2333 ( .CLK(n2450), .C(n2451) );
  BUFFD0 U2334 ( .I(n2451), .Z(n2452) );
  CKBD0 U2335 ( .CLK(n2452), .C(n2453) );
  CKBD0 U2336 ( .CLK(n2453), .C(n2454) );
  CKBD0 U2337 ( .CLK(n2454), .C(n2455) );
  CKBD0 U2338 ( .CLK(n2455), .C(n2456) );
  CKBD0 U2339 ( .CLK(n2456), .C(n2457) );
  CKBD0 U2340 ( .CLK(n2457), .C(n2458) );
  CKBD0 U2341 ( .CLK(n2458), .C(n2459) );
  CKBD0 U2342 ( .CLK(n2459), .C(n2460) );
  CKBD0 U2343 ( .CLK(n2460), .C(n2461) );
  CKBD0 U2344 ( .CLK(n2461), .C(n2462) );
  BUFFD0 U2345 ( .I(n2462), .Z(n2463) );
  CKBD0 U2346 ( .CLK(n2463), .C(n2464) );
  CKBD0 U2347 ( .CLK(n2464), .C(n2465) );
  CKBD0 U2348 ( .CLK(n2465), .C(n2466) );
  CKBD0 U2349 ( .CLK(n2466), .C(n2467) );
  BUFFD0 U2350 ( .I(n2467), .Z(n2468) );
  CKBD0 U2351 ( .CLK(n2468), .C(n2469) );
  BUFFD0 U2352 ( .I(n2469), .Z(n2470) );
  CKBD0 U2353 ( .CLK(n2470), .C(n2471) );
  BUFFD0 U2354 ( .I(n2471), .Z(n2472) );
  CKBD0 U2355 ( .CLK(n2472), .C(n2473) );
  BUFFD0 U2356 ( .I(n2473), .Z(n2474) );
  CKBD0 U2357 ( .CLK(n2474), .C(n2475) );
  BUFFD0 U2358 ( .I(n2475), .Z(n2476) );
  CKBD0 U2359 ( .CLK(n2476), .C(n2477) );
  BUFFD0 U2360 ( .I(n2477), .Z(n2478) );
  CKBD0 U2361 ( .CLK(n2478), .C(n2479) );
  BUFFD0 U2362 ( .I(n2479), .Z(n2480) );
  CKBD0 U2363 ( .CLK(n2480), .C(n2481) );
  BUFFD0 U2364 ( .I(n2481), .Z(n2482) );
  CKBD0 U2365 ( .CLK(n2482), .C(n2483) );
  BUFFD0 U2366 ( .I(n2483), .Z(n2484) );
  CKBD0 U2367 ( .CLK(n2484), .C(n2485) );
  BUFFD0 U2368 ( .I(n2485), .Z(n2486) );
  CKBD0 U2369 ( .CLK(n2486), .C(n2487) );
  BUFFD0 U2370 ( .I(n2487), .Z(n2488) );
  CKBD0 U2371 ( .CLK(n2488), .C(n2489) );
  BUFFD0 U2372 ( .I(n2489), .Z(n2490) );
  CKBD0 U2373 ( .CLK(n2490), .C(n2491) );
  BUFFD0 U2374 ( .I(n2491), .Z(n2492) );
  CKBD0 U2375 ( .CLK(n2492), .C(n2493) );
  BUFFD0 U2376 ( .I(n2493), .Z(n2494) );
  CKBD0 U2377 ( .CLK(n2494), .C(n2495) );
  BUFFD0 U2378 ( .I(n2497), .Z(n2496) );
  BUFFD0 U2379 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2380 ( .I(n164), .Z(n2498) );
  BUFFD0 U2381 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2382 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2383 ( .I(n163), .Z(n2501) );
  CKBD0 U2384 ( .CLK(n5), .C(n2502) );
  CKBD0 U2385 ( .CLK(n2502), .C(n2503) );
  CKBD0 U2386 ( .CLK(n2503), .C(n2504) );
  BUFFD0 U2387 ( .I(n2504), .Z(n2505) );
  CKBD0 U2388 ( .CLK(n2505), .C(n2506) );
  CKBD0 U2389 ( .CLK(n2506), .C(n2507) );
  CKBD0 U2390 ( .CLK(n2507), .C(n2508) );
  CKBD0 U2391 ( .CLK(n2508), .C(n2509) );
  CKBD0 U2392 ( .CLK(n2509), .C(n2510) );
  CKBD0 U2393 ( .CLK(n2510), .C(n2511) );
  CKBD0 U2394 ( .CLK(n2511), .C(n2512) );
  CKBD0 U2395 ( .CLK(n2512), .C(n2513) );
  CKBD0 U2396 ( .CLK(n2513), .C(n2514) );
  CKBD0 U2397 ( .CLK(n2514), .C(n2515) );
  BUFFD0 U2398 ( .I(n2515), .Z(n2516) );
  CKBD0 U2399 ( .CLK(n2516), .C(n2517) );
  CKBD0 U2400 ( .CLK(n2517), .C(n2518) );
  CKBD0 U2401 ( .CLK(n2518), .C(n2519) );
  CKBD0 U2402 ( .CLK(n2519), .C(n2520) );
  CKBD0 U2403 ( .CLK(n2520), .C(n2521) );
  CKBD0 U2404 ( .CLK(n2521), .C(n2522) );
  CKBD0 U2405 ( .CLK(n2522), .C(n2523) );
  CKBD0 U2406 ( .CLK(n2523), .C(n2524) );
  CKBD0 U2407 ( .CLK(n2524), .C(n2525) );
  CKBD0 U2408 ( .CLK(n2525), .C(n2526) );
  BUFFD0 U2409 ( .I(n2526), .Z(n2527) );
  CKBD0 U2410 ( .CLK(n2527), .C(n2528) );
  CKBD0 U2411 ( .CLK(n2528), .C(n2529) );
  CKBD0 U2412 ( .CLK(n2529), .C(n2530) );
  CKBD0 U2413 ( .CLK(n2530), .C(n2531) );
  CKBD0 U2414 ( .CLK(n2531), .C(n2532) );
  CKBD0 U2415 ( .CLK(n2532), .C(n2533) );
  CKBD0 U2416 ( .CLK(n2533), .C(n2534) );
  CKBD0 U2417 ( .CLK(n2534), .C(n2535) );
  CKBD0 U2418 ( .CLK(n2535), .C(n2536) );
  CKBD0 U2419 ( .CLK(n2536), .C(n2537) );
  BUFFD0 U2420 ( .I(n2537), .Z(n2538) );
  CKBD0 U2421 ( .CLK(n2538), .C(n2539) );
  CKBD0 U2422 ( .CLK(n2539), .C(n2540) );
  CKBD0 U2423 ( .CLK(n2540), .C(n2541) );
  CKBD0 U2424 ( .CLK(n2541), .C(n2542) );
  CKBD0 U2425 ( .CLK(n2542), .C(n2543) );
  CKBD0 U2426 ( .CLK(n2543), .C(n2544) );
  CKBD0 U2427 ( .CLK(n2544), .C(n2545) );
  CKBD0 U2428 ( .CLK(n2545), .C(n2546) );
  CKBD0 U2429 ( .CLK(n2546), .C(n2547) );
  CKBD0 U2430 ( .CLK(n2547), .C(n2548) );
  BUFFD0 U2431 ( .I(n2548), .Z(n2549) );
  CKBD0 U2432 ( .CLK(n2549), .C(n2550) );
  CKBD0 U2433 ( .CLK(n2550), .C(n2551) );
  CKBD0 U2434 ( .CLK(n2551), .C(n2552) );
  CKBD0 U2435 ( .CLK(n2552), .C(n2553) );
  CKBD0 U2436 ( .CLK(n2553), .C(n2554) );
  CKBD0 U2437 ( .CLK(n2554), .C(n2555) );
  CKBD0 U2438 ( .CLK(n2555), .C(n2556) );
  CKBD0 U2439 ( .CLK(n2556), .C(n2557) );
  CKBD0 U2440 ( .CLK(n2557), .C(n2558) );
  BUFFD0 U2441 ( .I(n2558), .Z(n2559) );
  CKBD0 U2442 ( .CLK(n2559), .C(n2560) );
  CKBD0 U2443 ( .CLK(n2560), .C(n2561) );
  CKBD0 U2444 ( .CLK(n2561), .C(n2562) );
  CKBD0 U2445 ( .CLK(n2562), .C(n2563) );
  CKBD0 U2446 ( .CLK(n2563), .C(n2564) );
  CKBD0 U2447 ( .CLK(n2564), .C(n2565) );
  CKBD0 U2448 ( .CLK(n2565), .C(n2566) );
  CKBD0 U2449 ( .CLK(n2566), .C(n2567) );
  CKBD0 U2450 ( .CLK(n2567), .C(n2568) );
  CKBD0 U2451 ( .CLK(n2568), .C(n2569) );
  CKBD0 U2452 ( .CLK(n2569), .C(n2570) );
  BUFFD0 U2453 ( .I(n2570), .Z(n2571) );
  CKBD0 U2454 ( .CLK(n2571), .C(n2572) );
  CKBD0 U2455 ( .CLK(n2572), .C(n2573) );
  CKBD0 U2456 ( .CLK(n2573), .C(n2574) );
  CKBD0 U2457 ( .CLK(n2574), .C(n2575) );
  CKBD0 U2458 ( .CLK(n2575), .C(n2576) );
  CKBD0 U2459 ( .CLK(n2576), .C(n2577) );
  CKBD0 U2460 ( .CLK(n2577), .C(n2578) );
  CKBD0 U2461 ( .CLK(n2578), .C(n2579) );
  CKBD0 U2462 ( .CLK(n2579), .C(n2580) );
  BUFFD0 U2463 ( .I(n2580), .Z(n2581) );
  CKBD0 U2464 ( .CLK(n2581), .C(n2582) );
  CKBD0 U2465 ( .CLK(n2582), .C(n2583) );
  CKBD0 U2466 ( .CLK(n2583), .C(n2584) );
  CKBD0 U2467 ( .CLK(n2584), .C(n2585) );
  CKBD0 U2468 ( .CLK(n2585), .C(n2586) );
  CKBD0 U2469 ( .CLK(n2586), .C(n2587) );
  CKBD0 U2470 ( .CLK(n2587), .C(n2588) );
  CKBD0 U2471 ( .CLK(n2588), .C(n2589) );
  CKBD0 U2472 ( .CLK(n2589), .C(n2590) );
  CKBD0 U2473 ( .CLK(n2590), .C(n2591) );
  BUFFD0 U2474 ( .I(n2591), .Z(n2592) );
  CKBD0 U2475 ( .CLK(n2592), .C(n2593) );
  CKBD0 U2476 ( .CLK(n2593), .C(n2594) );
  CKBD0 U2477 ( .CLK(n2594), .C(n2595) );
  CKBD0 U2478 ( .CLK(n2595), .C(n2596) );
  CKBD0 U2479 ( .CLK(n2596), .C(n2597) );
  CKBD0 U2480 ( .CLK(n2597), .C(n2598) );
  CKBD0 U2481 ( .CLK(n2598), .C(n2599) );
  CKBD0 U2482 ( .CLK(n2599), .C(n2600) );
  CKBD0 U2483 ( .CLK(n2600), .C(n2601) );
  CKBD0 U2484 ( .CLK(n2601), .C(n2602) );
  BUFFD0 U2485 ( .I(n2602), .Z(n2603) );
  CKBD0 U2486 ( .CLK(n2603), .C(n2604) );
  CKBD0 U2487 ( .CLK(n2604), .C(n2605) );
  CKBD0 U2488 ( .CLK(n2605), .C(n2606) );
  CKBD0 U2489 ( .CLK(n2606), .C(n2607) );
  CKBD0 U2490 ( .CLK(n2607), .C(n2608) );
  CKBD0 U2491 ( .CLK(n2608), .C(n2609) );
  CKBD0 U2492 ( .CLK(n2609), .C(n2610) );
  CKBD0 U2493 ( .CLK(n2610), .C(n2611) );
  CKBD0 U2494 ( .CLK(n2611), .C(n2612) );
  CKBD0 U2495 ( .CLK(n2612), .C(n2613) );
  BUFFD0 U2496 ( .I(n2613), .Z(n2614) );
  CKBD0 U2497 ( .CLK(n2614), .C(n2615) );
  CKBD0 U2498 ( .CLK(n2615), .C(n2616) );
  CKBD0 U2499 ( .CLK(n2616), .C(n2617) );
  CKBD0 U2500 ( .CLK(n2617), .C(n2618) );
  CKBD0 U2501 ( .CLK(n2618), .C(n2619) );
  BUFFD0 U2502 ( .I(n2619), .Z(n2620) );
  CKBD0 U2503 ( .CLK(n2620), .C(n2621) );
  BUFFD0 U2504 ( .I(n2621), .Z(n2622) );
  CKBD0 U2505 ( .CLK(n2622), .C(n2623) );
  BUFFD0 U2506 ( .I(n2623), .Z(n2624) );
  CKBD0 U2507 ( .CLK(n2624), .C(n2625) );
  BUFFD0 U2508 ( .I(n2625), .Z(n2626) );
  CKBD0 U2509 ( .CLK(n2626), .C(n2627) );
  BUFFD0 U2510 ( .I(n2627), .Z(n2628) );
  CKBD0 U2511 ( .CLK(n2628), .C(n2629) );
  BUFFD0 U2512 ( .I(n2629), .Z(n2630) );
  CKBD0 U2513 ( .CLK(n2630), .C(n2631) );
  BUFFD0 U2514 ( .I(n2631), .Z(n2632) );
  CKBD0 U2515 ( .CLK(n2632), .C(n2633) );
  BUFFD0 U2516 ( .I(n2633), .Z(n2634) );
  BUFFD0 U2517 ( .I(n2636), .Z(n2635) );
  BUFFD0 U2518 ( .I(n2637), .Z(n2636) );
  BUFFD0 U2519 ( .I(n162), .Z(n2637) );
  CKBD0 U2520 ( .CLK(n1269), .C(n2638) );
  CKBD0 U2521 ( .CLK(n2638), .C(n2639) );
  CKBD0 U2522 ( .CLK(n2639), .C(n2640) );
  CKBD0 U2523 ( .CLK(n2640), .C(n2641) );
  BUFFD0 U2524 ( .I(n2641), .Z(n2642) );
  CKBD0 U2525 ( .CLK(n2642), .C(n2643) );
  CKBD0 U2526 ( .CLK(n2643), .C(n2644) );
  CKBD0 U2527 ( .CLK(n2644), .C(n2645) );
  CKBD0 U2528 ( .CLK(n2645), .C(n2646) );
  CKBD0 U2529 ( .CLK(n2646), .C(n2647) );
  CKBD0 U2530 ( .CLK(n2647), .C(n2648) );
  CKBD0 U2531 ( .CLK(n2648), .C(n2649) );
  CKBD0 U2532 ( .CLK(n2649), .C(n2650) );
  CKBD0 U2533 ( .CLK(n2650), .C(n2651) );
  BUFFD0 U2534 ( .I(n2651), .Z(n2652) );
  CKBD0 U2535 ( .CLK(n2652), .C(n2653) );
  CKBD0 U2536 ( .CLK(n2653), .C(n2654) );
  CKBD0 U2537 ( .CLK(n2654), .C(n2655) );
  CKBD0 U2538 ( .CLK(n2655), .C(n2656) );
  CKBD0 U2539 ( .CLK(n2656), .C(n2657) );
  CKBD0 U2540 ( .CLK(n2657), .C(n2658) );
  CKBD0 U2541 ( .CLK(n2658), .C(n2659) );
  CKBD0 U2542 ( .CLK(n2659), .C(n2660) );
  CKBD0 U2543 ( .CLK(n2660), .C(n2661) );
  BUFFD0 U2544 ( .I(n2661), .Z(n2662) );
  CKBD0 U2545 ( .CLK(n2662), .C(n2663) );
  CKBD0 U2546 ( .CLK(n2663), .C(n2664) );
  CKBD0 U2547 ( .CLK(n2664), .C(n2665) );
  CKBD0 U2548 ( .CLK(n2665), .C(n2666) );
  CKBD0 U2549 ( .CLK(n2666), .C(n2667) );
  CKBD0 U2550 ( .CLK(n2667), .C(n2668) );
  CKBD0 U2551 ( .CLK(n2668), .C(n2669) );
  CKBD0 U2552 ( .CLK(n2669), .C(n2670) );
  CKBD0 U2553 ( .CLK(n2670), .C(n2671) );
  CKBD0 U2554 ( .CLK(n2671), .C(n2672) );
  CKBD0 U2555 ( .CLK(n2672), .C(n2673) );
  BUFFD0 U2556 ( .I(n2673), .Z(n2674) );
  CKBD0 U2557 ( .CLK(n2674), .C(n2675) );
  CKBD0 U2558 ( .CLK(n2675), .C(n2676) );
  CKBD0 U2559 ( .CLK(n2676), .C(n2677) );
  CKBD0 U2560 ( .CLK(n2677), .C(n2678) );
  CKBD0 U2561 ( .CLK(n2678), .C(n2679) );
  CKBD0 U2562 ( .CLK(n2679), .C(n2680) );
  CKBD0 U2563 ( .CLK(n2680), .C(n2681) );
  CKBD0 U2564 ( .CLK(n2681), .C(n2682) );
  CKBD0 U2565 ( .CLK(n2682), .C(n2683) );
  CKBD0 U2566 ( .CLK(n2683), .C(n2684) );
  BUFFD0 U2567 ( .I(n2684), .Z(n2685) );
  CKBD0 U2568 ( .CLK(n2685), .C(n2686) );
  CKBD0 U2569 ( .CLK(n2686), .C(n2687) );
  CKBD0 U2570 ( .CLK(n2687), .C(n2688) );
  CKBD0 U2571 ( .CLK(n2688), .C(n2689) );
  CKBD0 U2572 ( .CLK(n2689), .C(n2690) );
  CKBD0 U2573 ( .CLK(n2690), .C(n2691) );
  CKBD0 U2574 ( .CLK(n2691), .C(n2692) );
  CKBD0 U2575 ( .CLK(n2692), .C(n2693) );
  CKBD0 U2576 ( .CLK(n2693), .C(n2694) );
  BUFFD0 U2577 ( .I(n2694), .Z(n2695) );
  CKBD0 U2578 ( .CLK(n2695), .C(n2696) );
  CKBD0 U2579 ( .CLK(n2696), .C(n2697) );
  CKBD0 U2580 ( .CLK(n2697), .C(n2698) );
  CKBD0 U2581 ( .CLK(n2698), .C(n2699) );
  CKBD0 U2582 ( .CLK(n2699), .C(n2700) );
  CKBD0 U2583 ( .CLK(n2700), .C(n2701) );
  CKBD0 U2584 ( .CLK(n2701), .C(n2702) );
  CKBD0 U2585 ( .CLK(n2702), .C(n2703) );
  CKBD0 U2586 ( .CLK(n2703), .C(n2704) );
  CKBD0 U2587 ( .CLK(n2704), .C(n2705) );
  CKBD0 U2588 ( .CLK(n2705), .C(n2706) );
  BUFFD0 U2589 ( .I(n2706), .Z(n2707) );
  CKBD0 U2590 ( .CLK(n2707), .C(n2708) );
  CKBD0 U2591 ( .CLK(n2708), .C(n2709) );
  CKBD0 U2592 ( .CLK(n2709), .C(n2710) );
  CKBD0 U2593 ( .CLK(n2710), .C(n2711) );
  CKBD0 U2594 ( .CLK(n2711), .C(n2712) );
  CKBD0 U2595 ( .CLK(n2712), .C(n2713) );
  CKBD0 U2596 ( .CLK(n2713), .C(n2714) );
  CKBD0 U2597 ( .CLK(n2714), .C(n2715) );
  CKBD0 U2598 ( .CLK(n2715), .C(n2716) );
  BUFFD0 U2599 ( .I(n2716), .Z(n2717) );
  CKBD0 U2600 ( .CLK(n2717), .C(n2718) );
  CKBD0 U2601 ( .CLK(n2718), .C(n2719) );
  CKBD0 U2602 ( .CLK(n2719), .C(n2720) );
  CKBD0 U2603 ( .CLK(n2720), .C(n2721) );
  CKBD0 U2604 ( .CLK(n2721), .C(n2722) );
  CKBD0 U2605 ( .CLK(n2722), .C(n2723) );
  CKBD0 U2606 ( .CLK(n2723), .C(n2724) );
  CKBD0 U2607 ( .CLK(n2724), .C(n2725) );
  CKBD0 U2608 ( .CLK(n2725), .C(n2726) );
  BUFFD0 U2609 ( .I(n2726), .Z(n2727) );
  CKBD0 U2610 ( .CLK(n2727), .C(n2728) );
  CKBD0 U2611 ( .CLK(n2728), .C(n2729) );
  CKBD0 U2612 ( .CLK(n2729), .C(n2730) );
  CKBD0 U2613 ( .CLK(n2730), .C(n2731) );
  CKBD0 U2614 ( .CLK(n2731), .C(n2732) );
  CKBD0 U2615 ( .CLK(n2732), .C(n2733) );
  CKBD0 U2616 ( .CLK(n2733), .C(n2734) );
  CKBD0 U2617 ( .CLK(n2734), .C(n2735) );
  CKBD0 U2618 ( .CLK(n2735), .C(n2736) );
  CKBD0 U2619 ( .CLK(n2736), .C(n2737) );
  CKBD0 U2620 ( .CLK(n2737), .C(n2738) );
  BUFFD0 U2621 ( .I(n2738), .Z(n2739) );
  CKBD0 U2622 ( .CLK(n2739), .C(n2740) );
  CKBD0 U2623 ( .CLK(n2740), .C(n2741) );
  CKBD0 U2624 ( .CLK(n2741), .C(n2742) );
  CKBD0 U2625 ( .CLK(n2742), .C(n2743) );
  CKBD0 U2626 ( .CLK(n2743), .C(n2744) );
  CKBD0 U2627 ( .CLK(n2744), .C(n2745) );
  CKBD0 U2628 ( .CLK(n2745), .C(n2746) );
  CKBD0 U2629 ( .CLK(n2746), .C(n2747) );
  CKBD0 U2630 ( .CLK(n2747), .C(n2748) );
  CKBD0 U2631 ( .CLK(n2748), .C(n2749) );
  BUFFD0 U2632 ( .I(n2749), .Z(n2750) );
  CKBD0 U2633 ( .CLK(n2750), .C(n2751) );
  CKBD0 U2634 ( .CLK(n2751), .C(n2752) );
  CKBD0 U2635 ( .CLK(n2752), .C(n2753) );
  CKBD0 U2636 ( .CLK(n2753), .C(n2754) );
  CKBD0 U2637 ( .CLK(n2754), .C(n2755) );
  BUFFD0 U2638 ( .I(n2755), .Z(n2756) );
  CKBD0 U2639 ( .CLK(n2756), .C(n2757) );
  BUFFD0 U2640 ( .I(n2757), .Z(n2758) );
  CKBD0 U2641 ( .CLK(n2758), .C(n2759) );
  BUFFD0 U2642 ( .I(n2759), .Z(n2760) );
  CKBD0 U2643 ( .CLK(n2760), .C(n2761) );
  BUFFD0 U2644 ( .I(n2761), .Z(n2762) );
  CKBD0 U2645 ( .CLK(n2762), .C(n2763) );
  BUFFD0 U2646 ( .I(n2763), .Z(n2764) );
  CKBD0 U2647 ( .CLK(n2764), .C(n2765) );
  BUFFD0 U2648 ( .I(n2765), .Z(n2766) );
  CKBD0 U2649 ( .CLK(n2766), .C(n2767) );
  BUFFD0 U2650 ( .I(n2767), .Z(n2768) );
  CKBD0 U2651 ( .CLK(n2768), .C(n2769) );
  BUFFD0 U2652 ( .I(n2769), .Z(n2770) );
  BUFFD0 U2653 ( .I(n2772), .Z(n2771) );
  BUFFD0 U2654 ( .I(n2773), .Z(n2772) );
  BUFFD0 U2655 ( .I(n161), .Z(n2773) );
  CKBD0 U2656 ( .CLK(n1267), .C(n2774) );
  CKBD0 U2657 ( .CLK(n2774), .C(n2775) );
  CKBD0 U2658 ( .CLK(n2775), .C(n2776) );
  BUFFD0 U2659 ( .I(n2776), .Z(n2777) );
  CKBD0 U2660 ( .CLK(n2777), .C(n2778) );
  CKBD0 U2661 ( .CLK(n2778), .C(n2779) );
  CKBD0 U2662 ( .CLK(n2779), .C(n2780) );
  CKBD0 U2663 ( .CLK(n2780), .C(n2781) );
  CKBD0 U2664 ( .CLK(n2781), .C(n2782) );
  CKBD0 U2665 ( .CLK(n2782), .C(n2783) );
  CKBD0 U2666 ( .CLK(n2783), .C(n2784) );
  CKBD0 U2667 ( .CLK(n2784), .C(n2785) );
  CKBD0 U2668 ( .CLK(n2785), .C(n2786) );
  CKBD0 U2669 ( .CLK(n2786), .C(n2787) );
  BUFFD0 U2670 ( .I(n2787), .Z(n2788) );
  CKBD0 U2671 ( .CLK(n2788), .C(n2789) );
  CKBD0 U2672 ( .CLK(n2789), .C(n2790) );
  CKBD0 U2673 ( .CLK(n2790), .C(n2791) );
  CKBD0 U2674 ( .CLK(n2791), .C(n2792) );
  CKBD0 U2675 ( .CLK(n2792), .C(n2793) );
  CKBD0 U2676 ( .CLK(n2793), .C(n2794) );
  CKBD0 U2677 ( .CLK(n2794), .C(n2795) );
  CKBD0 U2678 ( .CLK(n2795), .C(n2796) );
  CKBD0 U2679 ( .CLK(n2796), .C(n2797) );
  CKBD0 U2680 ( .CLK(n2797), .C(n2798) );
  BUFFD0 U2681 ( .I(n2798), .Z(n2799) );
  CKBD0 U2682 ( .CLK(n2799), .C(n2800) );
  CKBD0 U2683 ( .CLK(n2800), .C(n2801) );
  CKBD0 U2684 ( .CLK(n2801), .C(n2802) );
  CKBD0 U2685 ( .CLK(n2802), .C(n2803) );
  CKBD0 U2686 ( .CLK(n2803), .C(n2804) );
  CKBD0 U2687 ( .CLK(n2804), .C(n2805) );
  CKBD0 U2688 ( .CLK(n2805), .C(n2806) );
  CKBD0 U2689 ( .CLK(n2806), .C(n2807) );
  CKBD0 U2690 ( .CLK(n2807), .C(n2808) );
  CKBD0 U2691 ( .CLK(n2808), .C(n2809) );
  BUFFD0 U2692 ( .I(n2809), .Z(n2810) );
  CKBD0 U2693 ( .CLK(n2810), .C(n2811) );
  CKBD0 U2694 ( .CLK(n2811), .C(n2812) );
  CKBD0 U2695 ( .CLK(n2812), .C(n2813) );
  CKBD0 U2696 ( .CLK(n2813), .C(n2814) );
  CKBD0 U2697 ( .CLK(n2814), .C(n2815) );
  CKBD0 U2698 ( .CLK(n2815), .C(n2816) );
  CKBD0 U2699 ( .CLK(n2816), .C(n2817) );
  CKBD0 U2700 ( .CLK(n2817), .C(n2818) );
  CKBD0 U2701 ( .CLK(n2818), .C(n2819) );
  BUFFD0 U2702 ( .I(n2819), .Z(n2820) );
  CKBD0 U2703 ( .CLK(n2820), .C(n2821) );
  CKBD0 U2704 ( .CLK(n2821), .C(n2822) );
  CKBD0 U2705 ( .CLK(n2822), .C(n2823) );
  CKBD0 U2706 ( .CLK(n2823), .C(n2824) );
  CKBD0 U2707 ( .CLK(n2824), .C(n2825) );
  CKBD0 U2708 ( .CLK(n2825), .C(n2826) );
  CKBD0 U2709 ( .CLK(n2826), .C(n2827) );
  CKBD0 U2710 ( .CLK(n2827), .C(n2828) );
  CKBD0 U2711 ( .CLK(n2828), .C(n2829) );
  CKBD0 U2712 ( .CLK(n2829), .C(n2830) );
  CKBD0 U2713 ( .CLK(n2830), .C(n2831) );
  BUFFD0 U2714 ( .I(n2831), .Z(n2832) );
  CKBD0 U2715 ( .CLK(n2832), .C(n2833) );
  CKBD0 U2716 ( .CLK(n2833), .C(n2834) );
  CKBD0 U2717 ( .CLK(n2834), .C(n2835) );
  CKBD0 U2718 ( .CLK(n2835), .C(n2836) );
  CKBD0 U2719 ( .CLK(n2836), .C(n2837) );
  CKBD0 U2720 ( .CLK(n2837), .C(n2838) );
  CKBD0 U2721 ( .CLK(n2838), .C(n2839) );
  CKBD0 U2722 ( .CLK(n2839), .C(n2840) );
  CKBD0 U2723 ( .CLK(n2840), .C(n2841) );
  BUFFD0 U2724 ( .I(n2841), .Z(n2842) );
  CKBD0 U2725 ( .CLK(n2842), .C(n2843) );
  CKBD0 U2726 ( .CLK(n2843), .C(n2844) );
  CKBD0 U2727 ( .CLK(n2844), .C(n2845) );
  CKBD0 U2728 ( .CLK(n2845), .C(n2846) );
  CKBD0 U2729 ( .CLK(n2846), .C(n2847) );
  CKBD0 U2730 ( .CLK(n2847), .C(n2848) );
  CKBD0 U2731 ( .CLK(n2848), .C(n2849) );
  CKBD0 U2732 ( .CLK(n2849), .C(n2850) );
  CKBD0 U2733 ( .CLK(n2850), .C(n2851) );
  CKBD0 U2734 ( .CLK(n2851), .C(n2852) );
  BUFFD0 U2735 ( .I(n2852), .Z(n2853) );
  CKBD0 U2736 ( .CLK(n2853), .C(n2854) );
  CKBD0 U2737 ( .CLK(n2854), .C(n2855) );
  CKBD0 U2738 ( .CLK(n2855), .C(n2856) );
  CKBD0 U2739 ( .CLK(n2856), .C(n2857) );
  CKBD0 U2740 ( .CLK(n2857), .C(n2858) );
  CKBD0 U2741 ( .CLK(n2858), .C(n2859) );
  CKBD0 U2742 ( .CLK(n2859), .C(n2860) );
  CKBD0 U2743 ( .CLK(n2860), .C(n2861) );
  CKBD0 U2744 ( .CLK(n2861), .C(n2862) );
  CKBD0 U2745 ( .CLK(n2862), .C(n2863) );
  CKBD0 U2746 ( .CLK(n2863), .C(n2864) );
  BUFFD0 U2747 ( .I(n2864), .Z(n2865) );
  CKBD0 U2748 ( .CLK(n2865), .C(n2866) );
  CKBD0 U2749 ( .CLK(n2866), .C(n2867) );
  CKBD0 U2750 ( .CLK(n2867), .C(n2868) );
  CKBD0 U2751 ( .CLK(n2868), .C(n2869) );
  CKBD0 U2752 ( .CLK(n2869), .C(n2870) );
  CKBD0 U2753 ( .CLK(n2870), .C(n2871) );
  CKBD0 U2754 ( .CLK(n2871), .C(n2872) );
  CKBD0 U2755 ( .CLK(n2872), .C(n2873) );
  CKBD0 U2756 ( .CLK(n2873), .C(n2874) );
  BUFFD0 U2757 ( .I(n2874), .Z(n2875) );
  CKBD0 U2758 ( .CLK(n2875), .C(n2876) );
  CKBD0 U2759 ( .CLK(n2876), .C(n2877) );
  CKBD0 U2760 ( .CLK(n2877), .C(n2878) );
  CKBD0 U2761 ( .CLK(n2878), .C(n2879) );
  CKBD0 U2762 ( .CLK(n2879), .C(n2880) );
  CKBD0 U2763 ( .CLK(n2880), .C(n2881) );
  CKBD0 U2764 ( .CLK(n2881), .C(n2882) );
  CKBD0 U2765 ( .CLK(n2882), .C(n2883) );
  CKBD0 U2766 ( .CLK(n2883), .C(n2884) );
  BUFFD0 U2767 ( .I(n2884), .Z(n2885) );
  CKBD0 U2768 ( .CLK(n2885), .C(n2886) );
  CKBD0 U2769 ( .CLK(n2886), .C(n2887) );
  CKBD0 U2770 ( .CLK(n2887), .C(n2888) );
  CKBD0 U2771 ( .CLK(n2888), .C(n2889) );
  CKBD0 U2772 ( .CLK(n2889), .C(n2890) );
  CKBD0 U2773 ( .CLK(n2890), .C(n2891) );
  BUFFD0 U2774 ( .I(n2891), .Z(n2892) );
  CKBD0 U2775 ( .CLK(n2892), .C(n2893) );
  BUFFD0 U2776 ( .I(n2893), .Z(n2894) );
  CKBD0 U2777 ( .CLK(n2894), .C(n2895) );
  BUFFD0 U2778 ( .I(n2895), .Z(n2896) );
  CKBD0 U2779 ( .CLK(n2896), .C(n2897) );
  BUFFD0 U2780 ( .I(n2897), .Z(n2898) );
  CKBD0 U2781 ( .CLK(n2898), .C(n2899) );
  BUFFD0 U2782 ( .I(n2899), .Z(n2900) );
  CKBD0 U2783 ( .CLK(n2900), .C(n2901) );
  BUFFD0 U2784 ( .I(n2901), .Z(n2902) );
  CKBD0 U2785 ( .CLK(n2902), .C(n2903) );
  BUFFD0 U2786 ( .I(n2903), .Z(n2904) );
  CKBD0 U2787 ( .CLK(n2904), .C(n2905) );
  BUFFD0 U2788 ( .I(n2905), .Z(n2906) );
  BUFFD0 U2789 ( .I(n2908), .Z(n2907) );
  BUFFD0 U2790 ( .I(n2909), .Z(n2908) );
  BUFFD0 U2791 ( .I(n160), .Z(n2909) );
  CKBD0 U2792 ( .CLK(n1265), .C(n2910) );
  CKBD0 U2793 ( .CLK(n2910), .C(n2911) );
  CKBD0 U2794 ( .CLK(n2911), .C(n2912) );
  BUFFD0 U2795 ( .I(n2912), .Z(n2913) );
  CKBD0 U2796 ( .CLK(n2913), .C(n2914) );
  CKBD0 U2797 ( .CLK(n2914), .C(n2915) );
  CKBD0 U2798 ( .CLK(n2915), .C(n2916) );
  CKBD0 U2799 ( .CLK(n2916), .C(n2917) );
  CKBD0 U2800 ( .CLK(n2917), .C(n2918) );
  CKBD0 U2801 ( .CLK(n2918), .C(n2919) );
  CKBD0 U2802 ( .CLK(n2919), .C(n2920) );
  CKBD0 U2803 ( .CLK(n2920), .C(n2921) );
  CKBD0 U2804 ( .CLK(n2921), .C(n2922) );
  CKBD0 U2805 ( .CLK(n2922), .C(n2923) );
  BUFFD0 U2806 ( .I(n2923), .Z(n2924) );
  CKBD0 U2807 ( .CLK(n2924), .C(n2925) );
  CKBD0 U2808 ( .CLK(n2925), .C(n2926) );
  CKBD0 U2809 ( .CLK(n2926), .C(n2927) );
  CKBD0 U2810 ( .CLK(n2927), .C(n2928) );
  CKBD0 U2811 ( .CLK(n2928), .C(n2929) );
  CKBD0 U2812 ( .CLK(n2929), .C(n2930) );
  CKBD0 U2813 ( .CLK(n2930), .C(n2931) );
  CKBD0 U2814 ( .CLK(n2931), .C(n2932) );
  CKBD0 U2815 ( .CLK(n2932), .C(n2933) );
  CKBD0 U2816 ( .CLK(n2933), .C(n2934) );
  BUFFD0 U2817 ( .I(n2934), .Z(n2935) );
  CKBD0 U2818 ( .CLK(n2935), .C(n2936) );
  CKBD0 U2819 ( .CLK(n2936), .C(n2937) );
  CKBD0 U2820 ( .CLK(n2937), .C(n2938) );
  CKBD0 U2821 ( .CLK(n2938), .C(n2939) );
  CKBD0 U2822 ( .CLK(n2939), .C(n2940) );
  CKBD0 U2823 ( .CLK(n2940), .C(n2941) );
  CKBD0 U2824 ( .CLK(n2941), .C(n2942) );
  CKBD0 U2825 ( .CLK(n2942), .C(n2943) );
  CKBD0 U2826 ( .CLK(n2943), .C(n2944) );
  CKBD0 U2827 ( .CLK(n2944), .C(n2945) );
  BUFFD0 U2828 ( .I(n2945), .Z(n2946) );
  CKBD0 U2829 ( .CLK(n2946), .C(n2947) );
  CKBD0 U2830 ( .CLK(n2947), .C(n2948) );
  CKBD0 U2831 ( .CLK(n2948), .C(n2949) );
  CKBD0 U2832 ( .CLK(n2949), .C(n2950) );
  CKBD0 U2833 ( .CLK(n2950), .C(n2951) );
  CKBD0 U2834 ( .CLK(n2951), .C(n2952) );
  CKBD0 U2835 ( .CLK(n2952), .C(n2953) );
  CKBD0 U2836 ( .CLK(n2953), .C(n2954) );
  CKBD0 U2837 ( .CLK(n2954), .C(n2955) );
  BUFFD0 U2838 ( .I(n2955), .Z(n2956) );
  CKBD0 U2839 ( .CLK(n2956), .C(n2957) );
  CKBD0 U2840 ( .CLK(n2957), .C(n2958) );
  CKBD0 U2841 ( .CLK(n2958), .C(n2959) );
  CKBD0 U2842 ( .CLK(n2959), .C(n2960) );
  CKBD0 U2843 ( .CLK(n2960), .C(n2961) );
  CKBD0 U2844 ( .CLK(n2961), .C(n2962) );
  CKBD0 U2845 ( .CLK(n2962), .C(n2963) );
  CKBD0 U2846 ( .CLK(n2963), .C(n2964) );
  CKBD0 U2847 ( .CLK(n2964), .C(n2965) );
  CKBD0 U2848 ( .CLK(n2965), .C(n2966) );
  CKBD0 U2849 ( .CLK(n2966), .C(n2967) );
  BUFFD0 U2850 ( .I(n2967), .Z(n2968) );
  CKBD0 U2851 ( .CLK(n2968), .C(n2969) );
  CKBD0 U2852 ( .CLK(n2969), .C(n2970) );
  CKBD0 U2853 ( .CLK(n2970), .C(n2971) );
  CKBD0 U2854 ( .CLK(n2971), .C(n2972) );
  CKBD0 U2855 ( .CLK(n2972), .C(n2973) );
  CKBD0 U2856 ( .CLK(n2973), .C(n2974) );
  CKBD0 U2857 ( .CLK(n2974), .C(n2975) );
  CKBD0 U2858 ( .CLK(n2975), .C(n2976) );
  CKBD0 U2859 ( .CLK(n2976), .C(n2977) );
  BUFFD0 U2860 ( .I(n2977), .Z(n2978) );
  CKBD0 U2861 ( .CLK(n2978), .C(n2979) );
  CKBD0 U2862 ( .CLK(n2979), .C(n2980) );
  CKBD0 U2863 ( .CLK(n2980), .C(n2981) );
  CKBD0 U2864 ( .CLK(n2981), .C(n2982) );
  CKBD0 U2865 ( .CLK(n2982), .C(n2983) );
  CKBD0 U2866 ( .CLK(n2983), .C(n2984) );
  CKBD0 U2867 ( .CLK(n2984), .C(n2985) );
  CKBD0 U2868 ( .CLK(n2985), .C(n2986) );
  CKBD0 U2869 ( .CLK(n2986), .C(n2987) );
  CKBD0 U2870 ( .CLK(n2987), .C(n2988) );
  BUFFD0 U2871 ( .I(n2988), .Z(n2989) );
  CKBD0 U2872 ( .CLK(n2989), .C(n2990) );
  CKBD0 U2873 ( .CLK(n2990), .C(n2991) );
  CKBD0 U2874 ( .CLK(n2991), .C(n2992) );
  CKBD0 U2875 ( .CLK(n2992), .C(n2993) );
  CKBD0 U2876 ( .CLK(n2993), .C(n2994) );
  CKBD0 U2877 ( .CLK(n2994), .C(n2995) );
  CKBD0 U2878 ( .CLK(n2995), .C(n2996) );
  CKBD0 U2879 ( .CLK(n2996), .C(n2997) );
  CKBD0 U2880 ( .CLK(n2997), .C(n2998) );
  CKBD0 U2881 ( .CLK(n2998), .C(n2999) );
  BUFFD0 U2882 ( .I(n2999), .Z(n3000) );
  CKBD0 U2883 ( .CLK(n3000), .C(n3001) );
  CKBD0 U2884 ( .CLK(n3001), .C(n3002) );
  CKBD0 U2885 ( .CLK(n3002), .C(n3003) );
  CKBD0 U2886 ( .CLK(n3003), .C(n3004) );
  CKBD0 U2887 ( .CLK(n3004), .C(n3005) );
  CKBD0 U2888 ( .CLK(n3005), .C(n3006) );
  CKBD0 U2889 ( .CLK(n3006), .C(n3007) );
  CKBD0 U2890 ( .CLK(n3007), .C(n3008) );
  CKBD0 U2891 ( .CLK(n3008), .C(n3009) );
  CKBD0 U2892 ( .CLK(n3009), .C(n3010) );
  BUFFD0 U2893 ( .I(n3010), .Z(n3011) );
  CKBD0 U2894 ( .CLK(n3011), .C(n3012) );
  CKBD0 U2895 ( .CLK(n3012), .C(n3013) );
  CKBD0 U2896 ( .CLK(n3013), .C(n3014) );
  CKBD0 U2897 ( .CLK(n3014), .C(n3015) );
  CKBD0 U2898 ( .CLK(n3015), .C(n3016) );
  CKBD0 U2899 ( .CLK(n3016), .C(n3017) );
  CKBD0 U2900 ( .CLK(n3017), .C(n3018) );
  CKBD0 U2901 ( .CLK(n3018), .C(n3019) );
  CKBD0 U2902 ( .CLK(n3019), .C(n3020) );
  BUFFD0 U2903 ( .I(n3020), .Z(n3021) );
  CKBD0 U2904 ( .CLK(n3021), .C(n3022) );
  CKBD0 U2905 ( .CLK(n3022), .C(n3023) );
  CKBD0 U2906 ( .CLK(n3023), .C(n3024) );
  CKBD0 U2907 ( .CLK(n3024), .C(n3025) );
  CKBD0 U2908 ( .CLK(n3025), .C(n3026) );
  CKBD0 U2909 ( .CLK(n3026), .C(n3027) );
  BUFFD0 U2910 ( .I(n3027), .Z(n3028) );
  CKBD0 U2911 ( .CLK(n3028), .C(n3029) );
  BUFFD0 U2912 ( .I(n3029), .Z(n3030) );
  CKBD0 U2913 ( .CLK(n3030), .C(n3031) );
  BUFFD0 U2914 ( .I(n3031), .Z(n3032) );
  CKBD0 U2915 ( .CLK(n3032), .C(n3033) );
  BUFFD0 U2916 ( .I(n3033), .Z(n3034) );
  CKBD0 U2917 ( .CLK(n3034), .C(n3035) );
  BUFFD0 U2918 ( .I(n3035), .Z(n3036) );
  CKBD0 U2919 ( .CLK(n3036), .C(n3037) );
  BUFFD0 U2920 ( .I(n3037), .Z(n3038) );
  CKBD0 U2921 ( .CLK(n3038), .C(n3039) );
  BUFFD0 U2922 ( .I(n3039), .Z(n3040) );
  CKBD0 U2923 ( .CLK(n3040), .C(n3041) );
  BUFFD0 U2924 ( .I(n3041), .Z(n3042) );
  BUFFD0 U2925 ( .I(n3044), .Z(n3043) );
  BUFFD0 U2926 ( .I(n3045), .Z(n3044) );
  BUFFD0 U2927 ( .I(n159), .Z(n3045) );
  CKBD0 U2928 ( .CLK(n1263), .C(n3046) );
  CKBD0 U2929 ( .CLK(n3046), .C(n3047) );
  CKBD0 U2930 ( .CLK(n3047), .C(n3048) );
  BUFFD0 U2931 ( .I(n3048), .Z(n3049) );
  CKBD0 U2932 ( .CLK(n3049), .C(n3050) );
  CKBD0 U2933 ( .CLK(n3050), .C(n3051) );
  CKBD0 U2934 ( .CLK(n3051), .C(n3052) );
  CKBD0 U2935 ( .CLK(n3052), .C(n3053) );
  CKBD0 U2936 ( .CLK(n3053), .C(n3054) );
  CKBD0 U2937 ( .CLK(n3054), .C(n3055) );
  CKBD0 U2938 ( .CLK(n3055), .C(n3056) );
  CKBD0 U2939 ( .CLK(n3056), .C(n3057) );
  CKBD0 U2940 ( .CLK(n3057), .C(n3058) );
  BUFFD0 U2941 ( .I(n3058), .Z(n3059) );
  CKBD0 U2942 ( .CLK(n3059), .C(n3060) );
  CKBD0 U2943 ( .CLK(n3060), .C(n3061) );
  CKBD0 U2944 ( .CLK(n3061), .C(n3062) );
  CKBD0 U2945 ( .CLK(n3062), .C(n3063) );
  CKBD0 U2946 ( .CLK(n3063), .C(n3064) );
  CKBD0 U2947 ( .CLK(n3064), .C(n3065) );
  CKBD0 U2948 ( .CLK(n3065), .C(n3066) );
  CKBD0 U2949 ( .CLK(n3066), .C(n3067) );
  CKBD0 U2950 ( .CLK(n3067), .C(n3068) );
  CKBD0 U2951 ( .CLK(n3068), .C(n3069) );
  CKBD0 U2952 ( .CLK(n3069), .C(n3070) );
  BUFFD0 U2953 ( .I(n3070), .Z(n3071) );
  CKBD0 U2954 ( .CLK(n3071), .C(n3072) );
  CKBD0 U2955 ( .CLK(n3072), .C(n3073) );
  CKBD0 U2956 ( .CLK(n3073), .C(n3074) );
  CKBD0 U2957 ( .CLK(n3074), .C(n3075) );
  CKBD0 U2958 ( .CLK(n3075), .C(n3076) );
  CKBD0 U2959 ( .CLK(n3076), .C(n3077) );
  CKBD0 U2960 ( .CLK(n3077), .C(n3078) );
  CKBD0 U2961 ( .CLK(n3078), .C(n3079) );
  CKBD0 U2962 ( .CLK(n3079), .C(n3080) );
  CKBD0 U2963 ( .CLK(n3080), .C(n3081) );
  BUFFD0 U2964 ( .I(n3081), .Z(n3082) );
  CKBD0 U2965 ( .CLK(n3082), .C(n3083) );
  CKBD0 U2966 ( .CLK(n3083), .C(n3084) );
  CKBD0 U2967 ( .CLK(n3084), .C(n3085) );
  CKBD0 U2968 ( .CLK(n3085), .C(n3086) );
  CKBD0 U2969 ( .CLK(n3086), .C(n3087) );
  CKBD0 U2970 ( .CLK(n3087), .C(n3088) );
  CKBD0 U2971 ( .CLK(n3088), .C(n3089) );
  CKBD0 U2972 ( .CLK(n3089), .C(n3090) );
  CKBD0 U2973 ( .CLK(n3090), .C(n3091) );
  CKBD0 U2974 ( .CLK(n3091), .C(n3092) );
  BUFFD0 U2975 ( .I(n3092), .Z(n3093) );
  CKBD0 U2976 ( .CLK(n3093), .C(n3094) );
  CKBD0 U2977 ( .CLK(n3094), .C(n3095) );
  CKBD0 U2978 ( .CLK(n3095), .C(n3096) );
  CKBD0 U2979 ( .CLK(n3096), .C(n3097) );
  CKBD0 U2980 ( .CLK(n3097), .C(n3098) );
  CKBD0 U2981 ( .CLK(n3098), .C(n3099) );
  CKBD0 U2982 ( .CLK(n3099), .C(n3100) );
  CKBD0 U2983 ( .CLK(n3100), .C(n3101) );
  CKBD0 U2984 ( .CLK(n3101), .C(n3102) );
  CKBD0 U2985 ( .CLK(n3102), .C(n3103) );
  BUFFD0 U2986 ( .I(n3103), .Z(n3104) );
  CKBD0 U2987 ( .CLK(n3104), .C(n3105) );
  CKBD0 U2988 ( .CLK(n3105), .C(n3106) );
  CKBD0 U2989 ( .CLK(n3106), .C(n3107) );
  CKBD0 U2990 ( .CLK(n3107), .C(n3108) );
  CKBD0 U2991 ( .CLK(n3108), .C(n3109) );
  CKBD0 U2992 ( .CLK(n3109), .C(n3110) );
  CKBD0 U2993 ( .CLK(n3110), .C(n3111) );
  CKBD0 U2994 ( .CLK(n3111), .C(n3112) );
  CKBD0 U2995 ( .CLK(n3112), .C(n3113) );
  BUFFD0 U2996 ( .I(n3113), .Z(n3114) );
  CKBD0 U2997 ( .CLK(n3114), .C(n3115) );
  CKBD0 U2998 ( .CLK(n3115), .C(n3116) );
  CKBD0 U2999 ( .CLK(n3116), .C(n3117) );
  CKBD0 U3000 ( .CLK(n3117), .C(n3118) );
  CKBD0 U3001 ( .CLK(n3118), .C(n3119) );
  CKBD0 U3002 ( .CLK(n3119), .C(n3120) );
  CKBD0 U3003 ( .CLK(n3120), .C(n3121) );
  CKBD0 U3004 ( .CLK(n3121), .C(n3122) );
  CKBD0 U3005 ( .CLK(n3122), .C(n3123) );
  CKBD0 U3006 ( .CLK(n3123), .C(n3124) );
  CKBD0 U3007 ( .CLK(n3124), .C(n3125) );
  BUFFD0 U3008 ( .I(n3125), .Z(n3126) );
  CKBD0 U3009 ( .CLK(n3126), .C(n3127) );
  CKBD0 U3010 ( .CLK(n3127), .C(n3128) );
  CKBD0 U3011 ( .CLK(n3128), .C(n3129) );
  CKBD0 U3012 ( .CLK(n3129), .C(n3130) );
  CKBD0 U3013 ( .CLK(n3130), .C(n3131) );
  CKBD0 U3014 ( .CLK(n3131), .C(n3132) );
  CKBD0 U3015 ( .CLK(n3132), .C(n3133) );
  CKBD0 U3016 ( .CLK(n3133), .C(n3134) );
  CKBD0 U3017 ( .CLK(n3134), .C(n3135) );
  BUFFD0 U3018 ( .I(n3135), .Z(n3136) );
  CKBD0 U3019 ( .CLK(n3136), .C(n3137) );
  CKBD0 U3020 ( .CLK(n3137), .C(n3138) );
  CKBD0 U3021 ( .CLK(n3138), .C(n3139) );
  CKBD0 U3022 ( .CLK(n3139), .C(n3140) );
  CKBD0 U3023 ( .CLK(n3140), .C(n3141) );
  CKBD0 U3024 ( .CLK(n3141), .C(n3142) );
  CKBD0 U3025 ( .CLK(n3142), .C(n3143) );
  CKBD0 U3026 ( .CLK(n3143), .C(n3144) );
  CKBD0 U3027 ( .CLK(n3144), .C(n3145) );
  CKBD0 U3028 ( .CLK(n3145), .C(n3146) );
  BUFFD0 U3029 ( .I(n3146), .Z(n3147) );
  CKBD0 U3030 ( .CLK(n3147), .C(n3148) );
  CKBD0 U3031 ( .CLK(n3148), .C(n3149) );
  CKBD0 U3032 ( .CLK(n3149), .C(n3150) );
  CKBD0 U3033 ( .CLK(n3150), .C(n3151) );
  CKBD0 U3034 ( .CLK(n3151), .C(n3152) );
  CKBD0 U3035 ( .CLK(n3152), .C(n3153) );
  CKBD0 U3036 ( .CLK(n3153), .C(n3154) );
  CKBD0 U3037 ( .CLK(n3154), .C(n3155) );
  CKBD0 U3038 ( .CLK(n3155), .C(n3156) );
  CKBD0 U3039 ( .CLK(n3156), .C(n3157) );
  BUFFD0 U3040 ( .I(n3157), .Z(n3158) );
  CKBD0 U3041 ( .CLK(n3158), .C(n3159) );
  CKBD0 U3042 ( .CLK(n3159), .C(n3160) );
  CKBD0 U3043 ( .CLK(n3160), .C(n3161) );
  CKBD0 U3044 ( .CLK(n3161), .C(n3162) );
  CKBD0 U3045 ( .CLK(n3162), .C(n3163) );
  BUFFD0 U3046 ( .I(n3163), .Z(n3164) );
  CKBD0 U3047 ( .CLK(n3164), .C(n3165) );
  BUFFD0 U3048 ( .I(n3165), .Z(n3166) );
  CKBD0 U3049 ( .CLK(n3166), .C(n3167) );
  BUFFD0 U3050 ( .I(n3167), .Z(n3168) );
  CKBD0 U3051 ( .CLK(n3168), .C(n3169) );
  BUFFD0 U3052 ( .I(n3169), .Z(n3170) );
  CKBD0 U3053 ( .CLK(n3170), .C(n3171) );
  BUFFD0 U3054 ( .I(n3171), .Z(n3172) );
  CKBD0 U3055 ( .CLK(n3172), .C(n3173) );
  BUFFD0 U3056 ( .I(n3173), .Z(n3174) );
  CKBD0 U3057 ( .CLK(n3174), .C(n3175) );
  BUFFD0 U3058 ( .I(n3175), .Z(n3176) );
  CKBD0 U3059 ( .CLK(n3176), .C(n3177) );
  BUFFD0 U3060 ( .I(n3177), .Z(n3178) );
  BUFFD0 U3061 ( .I(n3180), .Z(n3179) );
  BUFFD0 U3062 ( .I(n3181), .Z(n3180) );
  BUFFD0 U3063 ( .I(n158), .Z(n3181) );
  CKBD0 U3064 ( .CLK(n1261), .C(n3182) );
  CKBD0 U3065 ( .CLK(n3182), .C(n3183) );
  CKBD0 U3066 ( .CLK(n3183), .C(n3184) );
  BUFFD0 U3067 ( .I(n3184), .Z(n3185) );
  CKBD0 U3068 ( .CLK(n3185), .C(n3186) );
  CKBD0 U3069 ( .CLK(n3186), .C(n3187) );
  CKBD0 U3070 ( .CLK(n3187), .C(n3188) );
  CKBD0 U3071 ( .CLK(n3188), .C(n3189) );
  CKBD0 U3072 ( .CLK(n3189), .C(n3190) );
  CKBD0 U3073 ( .CLK(n3190), .C(n3191) );
  CKBD0 U3074 ( .CLK(n3191), .C(n3192) );
  CKBD0 U3075 ( .CLK(n3192), .C(n3193) );
  CKBD0 U3076 ( .CLK(n3193), .C(n3194) );
  CKBD0 U3077 ( .CLK(n3194), .C(n3195) );
  CKBD0 U3078 ( .CLK(n3195), .C(n3196) );
  BUFFD0 U3079 ( .I(n3196), .Z(n3197) );
  CKBD0 U3080 ( .CLK(n3197), .C(n3198) );
  CKBD0 U3081 ( .CLK(n3198), .C(n3199) );
  CKBD0 U3082 ( .CLK(n3199), .C(n3200) );
  CKBD0 U3083 ( .CLK(n3200), .C(n3201) );
  CKBD0 U3084 ( .CLK(n3201), .C(n3202) );
  CKBD0 U3085 ( .CLK(n3202), .C(n3203) );
  CKBD0 U3086 ( .CLK(n3203), .C(n3204) );
  CKBD0 U3087 ( .CLK(n3204), .C(n3205) );
  CKBD0 U3088 ( .CLK(n3205), .C(n3206) );
  BUFFD0 U3089 ( .I(n3206), .Z(n3207) );
  CKBD0 U3090 ( .CLK(n3207), .C(n3208) );
  CKBD0 U3091 ( .CLK(n3208), .C(n3209) );
  CKBD0 U3092 ( .CLK(n3209), .C(n3210) );
  CKBD0 U3093 ( .CLK(n3210), .C(n3211) );
  CKBD0 U3094 ( .CLK(n3211), .C(n3212) );
  CKBD0 U3095 ( .CLK(n3212), .C(n3213) );
  CKBD0 U3096 ( .CLK(n3213), .C(n3214) );
  CKBD0 U3097 ( .CLK(n3214), .C(n3215) );
  CKBD0 U3098 ( .CLK(n3215), .C(n3216) );
  BUFFD0 U3099 ( .I(n3216), .Z(n3217) );
  CKBD0 U3100 ( .CLK(n3217), .C(n3218) );
  CKBD0 U3101 ( .CLK(n3218), .C(n3219) );
  CKBD0 U3102 ( .CLK(n3219), .C(n3220) );
  CKBD0 U3103 ( .CLK(n3220), .C(n3221) );
  CKBD0 U3104 ( .CLK(n3221), .C(n3222) );
  CKBD0 U3105 ( .CLK(n3222), .C(n3223) );
  CKBD0 U3106 ( .CLK(n3223), .C(n3224) );
  CKBD0 U3107 ( .CLK(n3224), .C(n3225) );
  CKBD0 U3108 ( .CLK(n3225), .C(n3226) );
  CKBD0 U3109 ( .CLK(n3226), .C(n3227) );
  CKBD0 U3110 ( .CLK(n3227), .C(n3228) );
  BUFFD0 U3111 ( .I(n3228), .Z(n3229) );
  CKBD0 U3112 ( .CLK(n3229), .C(n3230) );
  CKBD0 U3113 ( .CLK(n3230), .C(n3231) );
  CKBD0 U3114 ( .CLK(n3231), .C(n3232) );
  CKBD0 U3115 ( .CLK(n3232), .C(n3233) );
  CKBD0 U3116 ( .CLK(n3233), .C(n3234) );
  CKBD0 U3117 ( .CLK(n3234), .C(n3235) );
  CKBD0 U3118 ( .CLK(n3235), .C(n3236) );
  CKBD0 U3119 ( .CLK(n3236), .C(n3237) );
  CKBD0 U3120 ( .CLK(n3237), .C(n3238) );
  BUFFD0 U3121 ( .I(n3238), .Z(n3239) );
  CKBD0 U3122 ( .CLK(n3239), .C(n3240) );
  CKBD0 U3123 ( .CLK(n3240), .C(n3241) );
  CKBD0 U3124 ( .CLK(n3241), .C(n3242) );
  CKBD0 U3125 ( .CLK(n3242), .C(n3243) );
  CKBD0 U3126 ( .CLK(n3243), .C(n3244) );
  CKBD0 U3127 ( .CLK(n3244), .C(n3245) );
  CKBD0 U3128 ( .CLK(n3245), .C(n3246) );
  CKBD0 U3129 ( .CLK(n3246), .C(n3247) );
  CKBD0 U3130 ( .CLK(n3247), .C(n3248) );
  CKBD0 U3131 ( .CLK(n3248), .C(n3249) );
  BUFFD0 U3132 ( .I(n3249), .Z(n3250) );
  CKBD0 U3133 ( .CLK(n3250), .C(n3251) );
  CKBD0 U3134 ( .CLK(n3251), .C(n3252) );
  CKBD0 U3135 ( .CLK(n3252), .C(n3253) );
  CKBD0 U3136 ( .CLK(n3253), .C(n3254) );
  CKBD0 U3137 ( .CLK(n3254), .C(n3255) );
  CKBD0 U3138 ( .CLK(n3255), .C(n3256) );
  CKBD0 U3139 ( .CLK(n3256), .C(n3257) );
  CKBD0 U3140 ( .CLK(n3257), .C(n3258) );
  CKBD0 U3141 ( .CLK(n3258), .C(n3259) );
  CKBD0 U3142 ( .CLK(n3259), .C(n3260) );
  CKBD0 U3143 ( .CLK(n3260), .C(n3261) );
  BUFFD0 U3144 ( .I(n3261), .Z(n3262) );
  CKBD0 U3145 ( .CLK(n3262), .C(n3263) );
  CKBD0 U3146 ( .CLK(n3263), .C(n3264) );
  CKBD0 U3147 ( .CLK(n3264), .C(n3265) );
  CKBD0 U3148 ( .CLK(n3265), .C(n3266) );
  CKBD0 U3149 ( .CLK(n3266), .C(n3267) );
  CKBD0 U3150 ( .CLK(n3267), .C(n3268) );
  CKBD0 U3151 ( .CLK(n3268), .C(n3269) );
  CKBD0 U3152 ( .CLK(n3269), .C(n3270) );
  CKBD0 U3153 ( .CLK(n3270), .C(n3271) );
  BUFFD0 U3154 ( .I(n3271), .Z(n3272) );
  CKBD0 U3155 ( .CLK(n3272), .C(n3273) );
  CKBD0 U3156 ( .CLK(n3273), .C(n3274) );
  CKBD0 U3157 ( .CLK(n3274), .C(n3275) );
  CKBD0 U3158 ( .CLK(n3275), .C(n3276) );
  CKBD0 U3159 ( .CLK(n3276), .C(n3277) );
  CKBD0 U3160 ( .CLK(n3277), .C(n3278) );
  CKBD0 U3161 ( .CLK(n3278), .C(n3279) );
  CKBD0 U3162 ( .CLK(n3279), .C(n3280) );
  CKBD0 U3163 ( .CLK(n3280), .C(n3281) );
  BUFFD0 U3164 ( .I(n3281), .Z(n3282) );
  CKBD0 U3165 ( .CLK(n3282), .C(n3283) );
  CKBD0 U3166 ( .CLK(n3283), .C(n3284) );
  CKBD0 U3167 ( .CLK(n3284), .C(n3285) );
  CKBD0 U3168 ( .CLK(n3285), .C(n3286) );
  CKBD0 U3169 ( .CLK(n3286), .C(n3287) );
  CKBD0 U3170 ( .CLK(n3287), .C(n3288) );
  CKBD0 U3171 ( .CLK(n3288), .C(n3289) );
  CKBD0 U3172 ( .CLK(n3289), .C(n3290) );
  CKBD0 U3173 ( .CLK(n3290), .C(n3291) );
  CKBD0 U3174 ( .CLK(n3291), .C(n3292) );
  CKBD0 U3175 ( .CLK(n3292), .C(n3293) );
  BUFFD0 U3176 ( .I(n3293), .Z(n3294) );
  CKBD0 U3177 ( .CLK(n3294), .C(n3295) );
  CKBD0 U3178 ( .CLK(n3295), .C(n3296) );
  CKBD0 U3179 ( .CLK(n3296), .C(n3297) );
  CKBD0 U3180 ( .CLK(n3297), .C(n3298) );
  CKBD0 U3181 ( .CLK(n3298), .C(n3299) );
  BUFFD0 U3182 ( .I(n3299), .Z(n3300) );
  CKBD0 U3183 ( .CLK(n3300), .C(n3301) );
  BUFFD0 U3184 ( .I(n3301), .Z(n3302) );
  CKBD0 U3185 ( .CLK(n3302), .C(n3303) );
  BUFFD0 U3186 ( .I(n3303), .Z(n3304) );
  CKBD0 U3187 ( .CLK(n3304), .C(n3305) );
  BUFFD0 U3188 ( .I(n3305), .Z(n3306) );
  CKBD0 U3189 ( .CLK(n3306), .C(n3307) );
  BUFFD0 U3190 ( .I(n3307), .Z(n3308) );
  CKBD0 U3191 ( .CLK(n3308), .C(n3309) );
  BUFFD0 U3192 ( .I(n3309), .Z(n3310) );
  CKBD0 U3193 ( .CLK(n3310), .C(n3311) );
  BUFFD0 U3194 ( .I(n3311), .Z(n3312) );
  CKBD0 U3195 ( .CLK(n3312), .C(n3313) );
  BUFFD0 U3196 ( .I(n3313), .Z(n3314) );
  BUFFD0 U3197 ( .I(n3316), .Z(n3315) );
  BUFFD0 U3198 ( .I(n3317), .Z(n3316) );
  BUFFD0 U3199 ( .I(n157), .Z(n3317) );
  CKBD0 U3200 ( .CLK(n1259), .C(n3318) );
  CKBD0 U3201 ( .CLK(n3318), .C(n3319) );
  CKBD0 U3202 ( .CLK(n3319), .C(n3320) );
  BUFFD0 U3203 ( .I(n3320), .Z(n3321) );
  CKBD0 U3204 ( .CLK(n3321), .C(n3322) );
  CKBD0 U3205 ( .CLK(n3322), .C(n3323) );
  CKBD0 U3206 ( .CLK(n3323), .C(n3324) );
  CKBD0 U3207 ( .CLK(n3324), .C(n3325) );
  CKBD0 U3208 ( .CLK(n3325), .C(n3326) );
  CKBD0 U3209 ( .CLK(n3326), .C(n3327) );
  CKBD0 U3210 ( .CLK(n3327), .C(n3328) );
  CKBD0 U3211 ( .CLK(n3328), .C(n3329) );
  CKBD0 U3212 ( .CLK(n3329), .C(n3330) );
  CKBD0 U3213 ( .CLK(n3330), .C(n3331) );
  BUFFD0 U3214 ( .I(n3331), .Z(n3332) );
  CKBD0 U3215 ( .CLK(n3332), .C(n3333) );
  CKBD0 U3216 ( .CLK(n3333), .C(n3334) );
  CKBD0 U3217 ( .CLK(n3334), .C(n3335) );
  CKBD0 U3218 ( .CLK(n3335), .C(n3336) );
  CKBD0 U3219 ( .CLK(n3336), .C(n3337) );
  CKBD0 U3220 ( .CLK(n3337), .C(n3338) );
  CKBD0 U3221 ( .CLK(n3338), .C(n3339) );
  CKBD0 U3222 ( .CLK(n3339), .C(n3340) );
  CKBD0 U3223 ( .CLK(n3340), .C(n3341) );
  CKBD0 U3224 ( .CLK(n3341), .C(n3342) );
  BUFFD0 U3225 ( .I(n3342), .Z(n3343) );
  CKBD0 U3226 ( .CLK(n3343), .C(n3344) );
  CKBD0 U3227 ( .CLK(n3344), .C(n3345) );
  CKBD0 U3228 ( .CLK(n3345), .C(n3346) );
  CKBD0 U3229 ( .CLK(n3346), .C(n3347) );
  CKBD0 U3230 ( .CLK(n3347), .C(n3348) );
  CKBD0 U3231 ( .CLK(n3348), .C(n3349) );
  CKBD0 U3232 ( .CLK(n3349), .C(n3350) );
  CKBD0 U3233 ( .CLK(n3350), .C(n3351) );
  CKBD0 U3234 ( .CLK(n3351), .C(n3352) );
  BUFFD0 U3235 ( .I(n3352), .Z(n3353) );
  CKBD0 U3236 ( .CLK(n3353), .C(n3354) );
  CKBD0 U3237 ( .CLK(n3354), .C(n3355) );
  CKBD0 U3238 ( .CLK(n3355), .C(n3356) );
  CKBD0 U3239 ( .CLK(n3356), .C(n3357) );
  CKBD0 U3240 ( .CLK(n3357), .C(n3358) );
  CKBD0 U3241 ( .CLK(n3358), .C(n3359) );
  CKBD0 U3242 ( .CLK(n3359), .C(n3360) );
  CKBD0 U3243 ( .CLK(n3360), .C(n3361) );
  CKBD0 U3244 ( .CLK(n3361), .C(n3362) );
  CKBD0 U3245 ( .CLK(n3362), .C(n3363) );
  CKBD0 U3246 ( .CLK(n3363), .C(n3364) );
  BUFFD0 U3247 ( .I(n3364), .Z(n3365) );
  CKBD0 U3248 ( .CLK(n3365), .C(n3366) );
  CKBD0 U3249 ( .CLK(n3366), .C(n3367) );
  CKBD0 U3250 ( .CLK(n3367), .C(n3368) );
  CKBD0 U3251 ( .CLK(n3368), .C(n3369) );
  CKBD0 U3252 ( .CLK(n3369), .C(n3370) );
  CKBD0 U3253 ( .CLK(n3370), .C(n3371) );
  CKBD0 U3254 ( .CLK(n3371), .C(n3372) );
  CKBD0 U3255 ( .CLK(n3372), .C(n3373) );
  CKBD0 U3256 ( .CLK(n3373), .C(n3374) );
  BUFFD0 U3257 ( .I(n3374), .Z(n3375) );
  CKBD0 U3258 ( .CLK(n3375), .C(n3376) );
  CKBD0 U3259 ( .CLK(n3376), .C(n3377) );
  CKBD0 U3260 ( .CLK(n3377), .C(n3378) );
  CKBD0 U3261 ( .CLK(n3378), .C(n3379) );
  CKBD0 U3262 ( .CLK(n3379), .C(n3380) );
  CKBD0 U3263 ( .CLK(n3380), .C(n3381) );
  CKBD0 U3264 ( .CLK(n3381), .C(n3382) );
  CKBD0 U3265 ( .CLK(n3382), .C(n3383) );
  CKBD0 U3266 ( .CLK(n3383), .C(n3384) );
  CKBD0 U3267 ( .CLK(n3384), .C(n3385) );
  CKBD0 U3268 ( .CLK(n3385), .C(n3386) );
  BUFFD0 U3269 ( .I(n3386), .Z(n3387) );
  CKBD0 U3270 ( .CLK(n3387), .C(n3388) );
  CKBD0 U3271 ( .CLK(n3388), .C(n3389) );
  CKBD0 U3272 ( .CLK(n3389), .C(n3390) );
  CKBD0 U3273 ( .CLK(n3390), .C(n3391) );
  CKBD0 U3274 ( .CLK(n3391), .C(n3392) );
  CKBD0 U3275 ( .CLK(n3392), .C(n3393) );
  CKBD0 U3276 ( .CLK(n3393), .C(n3394) );
  CKBD0 U3277 ( .CLK(n3394), .C(n3395) );
  CKBD0 U3278 ( .CLK(n3395), .C(n3396) );
  BUFFD0 U3279 ( .I(n3396), .Z(n3397) );
  CKBD0 U3280 ( .CLK(n3397), .C(n3398) );
  CKBD0 U3281 ( .CLK(n3398), .C(n3399) );
  CKBD0 U3282 ( .CLK(n3399), .C(n3400) );
  CKBD0 U3283 ( .CLK(n3400), .C(n3401) );
  CKBD0 U3284 ( .CLK(n3401), .C(n3402) );
  CKBD0 U3285 ( .CLK(n3402), .C(n3403) );
  CKBD0 U3286 ( .CLK(n3403), .C(n3404) );
  CKBD0 U3287 ( .CLK(n3404), .C(n3405) );
  CKBD0 U3288 ( .CLK(n3405), .C(n3406) );
  CKBD0 U3289 ( .CLK(n3406), .C(n3407) );
  BUFFD0 U3290 ( .I(n3407), .Z(n3408) );
  CKBD0 U3291 ( .CLK(n3408), .C(n3409) );
  CKBD0 U3292 ( .CLK(n3409), .C(n3410) );
  CKBD0 U3293 ( .CLK(n3410), .C(n3411) );
  CKBD0 U3294 ( .CLK(n3411), .C(n3412) );
  CKBD0 U3295 ( .CLK(n3412), .C(n3413) );
  CKBD0 U3296 ( .CLK(n3413), .C(n3414) );
  CKBD0 U3297 ( .CLK(n3414), .C(n3415) );
  CKBD0 U3298 ( .CLK(n3415), .C(n3416) );
  CKBD0 U3299 ( .CLK(n3416), .C(n3417) );
  CKBD0 U3300 ( .CLK(n3417), .C(n3418) );
  BUFFD0 U3301 ( .I(n3418), .Z(n3419) );
  CKBD0 U3302 ( .CLK(n3419), .C(n3420) );
  CKBD0 U3303 ( .CLK(n3420), .C(n3421) );
  CKBD0 U3304 ( .CLK(n3421), .C(n3422) );
  CKBD0 U3305 ( .CLK(n3422), .C(n3423) );
  CKBD0 U3306 ( .CLK(n3423), .C(n3424) );
  CKBD0 U3307 ( .CLK(n3424), .C(n3425) );
  CKBD0 U3308 ( .CLK(n3425), .C(n3426) );
  CKBD0 U3309 ( .CLK(n3426), .C(n3427) );
  CKBD0 U3310 ( .CLK(n3427), .C(n3428) );
  CKBD0 U3311 ( .CLK(n3428), .C(n3429) );
  BUFFD0 U3312 ( .I(n3429), .Z(n3430) );
  CKBD0 U3313 ( .CLK(n3430), .C(n3431) );
  CKBD0 U3314 ( .CLK(n3431), .C(n3432) );
  CKBD0 U3315 ( .CLK(n3432), .C(n3433) );
  CKBD0 U3316 ( .CLK(n3433), .C(n3434) );
  CKBD0 U3317 ( .CLK(n3434), .C(n3435) );
  BUFFD0 U3318 ( .I(n3435), .Z(n3436) );
  CKBD0 U3319 ( .CLK(n3436), .C(n3437) );
  BUFFD0 U3320 ( .I(n3437), .Z(n3438) );
  CKBD0 U3321 ( .CLK(n3438), .C(n3439) );
  BUFFD0 U3322 ( .I(n3439), .Z(n3440) );
  CKBD0 U3323 ( .CLK(n3440), .C(n3441) );
  BUFFD0 U3324 ( .I(n3441), .Z(n3442) );
  CKBD0 U3325 ( .CLK(n3442), .C(n3443) );
  BUFFD0 U3326 ( .I(n3443), .Z(n3444) );
  CKBD0 U3327 ( .CLK(n3444), .C(n3445) );
  BUFFD0 U3328 ( .I(n3445), .Z(n3446) );
  CKBD0 U3329 ( .CLK(n3446), .C(n3447) );
  BUFFD0 U3330 ( .I(n3447), .Z(n3448) );
  CKBD0 U3331 ( .CLK(n3448), .C(n3449) );
  BUFFD0 U3332 ( .I(n3449), .Z(n3450) );
  BUFFD0 U3333 ( .I(n3452), .Z(n3451) );
  BUFFD0 U3334 ( .I(n3453), .Z(n3452) );
  BUFFD0 U3335 ( .I(n156), .Z(n3453) );
  CKBD0 U3336 ( .CLK(n1726), .C(n3454) );
  CKBD0 U3337 ( .CLK(n3454), .C(n3455) );
  CKBD0 U3338 ( .CLK(n3455), .C(n3456) );
  CKBD0 U3339 ( .CLK(n3456), .C(n3457) );
  BUFFD0 U3340 ( .I(n3457), .Z(n3458) );
  CKBD0 U3341 ( .CLK(n3458), .C(n3459) );
  CKBD0 U3342 ( .CLK(n3459), .C(n3460) );
  CKBD0 U3343 ( .CLK(n3460), .C(n3461) );
  CKBD0 U3344 ( .CLK(n3461), .C(n3462) );
  CKBD0 U3345 ( .CLK(n3462), .C(n3463) );
  CKBD0 U3346 ( .CLK(n3463), .C(n3464) );
  CKBD0 U3347 ( .CLK(n3464), .C(n3465) );
  CKBD0 U3348 ( .CLK(n3465), .C(n3466) );
  CKBD0 U3349 ( .CLK(n3466), .C(n3467) );
  BUFFD0 U3350 ( .I(n3467), .Z(n3468) );
  CKBD0 U3351 ( .CLK(n3468), .C(n3469) );
  CKBD0 U3352 ( .CLK(n3469), .C(n3470) );
  CKBD0 U3353 ( .CLK(n3470), .C(n3471) );
  CKBD0 U3354 ( .CLK(n3471), .C(n3472) );
  CKBD0 U3355 ( .CLK(n3472), .C(n3473) );
  CKBD0 U3356 ( .CLK(n3473), .C(n3474) );
  CKBD0 U3357 ( .CLK(n3474), .C(n3475) );
  CKBD0 U3358 ( .CLK(n3475), .C(n3476) );
  CKBD0 U3359 ( .CLK(n3476), .C(n3477) );
  CKBD0 U3360 ( .CLK(n3477), .C(n3478) );
  BUFFD0 U3361 ( .I(n3478), .Z(n3479) );
  CKBD0 U3362 ( .CLK(n3479), .C(n3480) );
  CKBD0 U3363 ( .CLK(n3480), .C(n3481) );
  CKBD0 U3364 ( .CLK(n3481), .C(n3482) );
  CKBD0 U3365 ( .CLK(n3482), .C(n3483) );
  CKBD0 U3366 ( .CLK(n3483), .C(n3484) );
  CKBD0 U3367 ( .CLK(n3484), .C(n3485) );
  CKBD0 U3368 ( .CLK(n3485), .C(n3486) );
  CKBD0 U3369 ( .CLK(n3486), .C(n3487) );
  CKBD0 U3370 ( .CLK(n3487), .C(n3488) );
  CKBD0 U3371 ( .CLK(n3488), .C(n3489) );
  BUFFD0 U3372 ( .I(n3489), .Z(n3490) );
  CKBD0 U3373 ( .CLK(n3490), .C(n3491) );
  CKBD0 U3374 ( .CLK(n3491), .C(n3492) );
  CKBD0 U3375 ( .CLK(n3492), .C(n3493) );
  CKBD0 U3376 ( .CLK(n3493), .C(n3494) );
  CKBD0 U3377 ( .CLK(n3494), .C(n3495) );
  CKBD0 U3378 ( .CLK(n3495), .C(n3496) );
  CKBD0 U3379 ( .CLK(n3496), .C(n3497) );
  CKBD0 U3380 ( .CLK(n3497), .C(n3498) );
  CKBD0 U3381 ( .CLK(n3498), .C(n3499) );
  CKBD0 U3382 ( .CLK(n3499), .C(n3500) );
  BUFFD0 U3383 ( .I(n3500), .Z(n3501) );
  CKBD0 U3384 ( .CLK(n3501), .C(n3502) );
  CKBD0 U3385 ( .CLK(n3502), .C(n3503) );
  CKBD0 U3386 ( .CLK(n3503), .C(n3504) );
  CKBD0 U3387 ( .CLK(n3504), .C(n3505) );
  CKBD0 U3388 ( .CLK(n3505), .C(n3506) );
  CKBD0 U3389 ( .CLK(n3506), .C(n3507) );
  CKBD0 U3390 ( .CLK(n3507), .C(n3508) );
  CKBD0 U3391 ( .CLK(n3508), .C(n3509) );
  CKBD0 U3392 ( .CLK(n3509), .C(n3510) );
  BUFFD0 U3393 ( .I(n3510), .Z(n3511) );
  CKBD0 U3394 ( .CLK(n3511), .C(n3512) );
  CKBD0 U3395 ( .CLK(n3512), .C(n3513) );
  CKBD0 U3396 ( .CLK(n3513), .C(n3514) );
  CKBD0 U3397 ( .CLK(n3514), .C(n3515) );
  CKBD0 U3398 ( .CLK(n3515), .C(n3516) );
  CKBD0 U3399 ( .CLK(n3516), .C(n3517) );
  CKBD0 U3400 ( .CLK(n3517), .C(n3518) );
  CKBD0 U3401 ( .CLK(n3518), .C(n3519) );
  CKBD0 U3402 ( .CLK(n3519), .C(n3520) );
  CKBD0 U3403 ( .CLK(n3520), .C(n3521) );
  CKBD0 U3404 ( .CLK(n3521), .C(n3522) );
  BUFFD0 U3405 ( .I(n3522), .Z(n3523) );
  CKBD0 U3406 ( .CLK(n3523), .C(n3524) );
  CKBD0 U3407 ( .CLK(n3524), .C(n3525) );
  CKBD0 U3408 ( .CLK(n3525), .C(n3526) );
  CKBD0 U3409 ( .CLK(n3526), .C(n3527) );
  CKBD0 U3410 ( .CLK(n3527), .C(n3528) );
  CKBD0 U3411 ( .CLK(n3528), .C(n3529) );
  CKBD0 U3412 ( .CLK(n3529), .C(n3530) );
  CKBD0 U3413 ( .CLK(n3530), .C(n3531) );
  CKBD0 U3414 ( .CLK(n3531), .C(n3532) );
  BUFFD0 U3415 ( .I(n3532), .Z(n3533) );
  CKBD0 U3416 ( .CLK(n3533), .C(n3534) );
  CKBD0 U3417 ( .CLK(n3534), .C(n3535) );
  CKBD0 U3418 ( .CLK(n3535), .C(n3536) );
  CKBD0 U3419 ( .CLK(n3536), .C(n3537) );
  CKBD0 U3420 ( .CLK(n3537), .C(n3538) );
  CKBD0 U3421 ( .CLK(n3538), .C(n3539) );
  CKBD0 U3422 ( .CLK(n3539), .C(n3540) );
  CKBD0 U3423 ( .CLK(n3540), .C(n3541) );
  CKBD0 U3424 ( .CLK(n3541), .C(n3542) );
  CKBD0 U3425 ( .CLK(n3542), .C(n3543) );
  BUFFD0 U3426 ( .I(n3543), .Z(n3544) );
  CKBD0 U3427 ( .CLK(n3544), .C(n3545) );
  CKBD0 U3428 ( .CLK(n3545), .C(n3546) );
  CKBD0 U3429 ( .CLK(n3546), .C(n3547) );
  CKBD0 U3430 ( .CLK(n3547), .C(n3548) );
  CKBD0 U3431 ( .CLK(n3548), .C(n3549) );
  CKBD0 U3432 ( .CLK(n3549), .C(n3550) );
  CKBD0 U3433 ( .CLK(n3550), .C(n3551) );
  CKBD0 U3434 ( .CLK(n3551), .C(n3552) );
  CKBD0 U3435 ( .CLK(n3552), .C(n3553) );
  CKBD0 U3436 ( .CLK(n3553), .C(n3554) );
  BUFFD0 U3437 ( .I(n3554), .Z(n3555) );
  CKBD0 U3438 ( .CLK(n3555), .C(n3556) );
  CKBD0 U3439 ( .CLK(n3556), .C(n3557) );
  CKBD0 U3440 ( .CLK(n3557), .C(n3558) );
  CKBD0 U3441 ( .CLK(n3558), .C(n3559) );
  CKBD0 U3442 ( .CLK(n3559), .C(n3560) );
  CKBD0 U3443 ( .CLK(n3560), .C(n3561) );
  CKBD0 U3444 ( .CLK(n3561), .C(n3562) );
  CKBD0 U3445 ( .CLK(n3562), .C(n3563) );
  CKBD0 U3446 ( .CLK(n3563), .C(n3564) );
  CKBD0 U3447 ( .CLK(n3564), .C(n3565) );
  BUFFD0 U3448 ( .I(n3565), .Z(n3566) );
  CKBD0 U3449 ( .CLK(n3566), .C(n3567) );
  CKBD0 U3450 ( .CLK(n3567), .C(n3568) );
  CKBD0 U3451 ( .CLK(n3568), .C(n3569) );
  CKBD0 U3452 ( .CLK(n3569), .C(n3570) );
  CKBD0 U3453 ( .CLK(n3570), .C(n3571) );
  BUFFD0 U3454 ( .I(n3571), .Z(n3572) );
  CKBD0 U3455 ( .CLK(n3572), .C(n3573) );
  BUFFD0 U3456 ( .I(n3573), .Z(n3574) );
  CKBD0 U3457 ( .CLK(n3574), .C(n3575) );
  BUFFD0 U3458 ( .I(n3575), .Z(n3576) );
  CKBD0 U3459 ( .CLK(n3576), .C(n3577) );
  BUFFD0 U3460 ( .I(n3577), .Z(n3578) );
  CKBD0 U3461 ( .CLK(n3578), .C(n3579) );
  BUFFD0 U3462 ( .I(n3579), .Z(n3580) );
  CKBD0 U3463 ( .CLK(n3580), .C(n3581) );
  BUFFD0 U3464 ( .I(n3581), .Z(n3582) );
  CKBD0 U3465 ( .CLK(n3582), .C(n3583) );
  BUFFD0 U3466 ( .I(n3583), .Z(n3584) );
  CKBD0 U3467 ( .CLK(n3584), .C(n3585) );
  BUFFD0 U3468 ( .I(n3585), .Z(n3586) );
  BUFFD0 U3469 ( .I(n3588), .Z(n3587) );
  BUFFD0 U3470 ( .I(n3589), .Z(n3588) );
  BUFFD0 U3471 ( .I(n155), .Z(n3589) );
  CKBD0 U3472 ( .CLK(n1167), .C(n3590) );
  CKBD0 U3473 ( .CLK(n3590), .C(n3591) );
  CKBD0 U3474 ( .CLK(n3591), .C(n3592) );
  CKBD0 U3475 ( .CLK(n3592), .C(n3593) );
  BUFFD0 U3476 ( .I(n3593), .Z(n3594) );
  CKBD0 U3477 ( .CLK(n3594), .C(n3595) );
  CKBD0 U3478 ( .CLK(n3595), .C(n3596) );
  CKBD0 U3479 ( .CLK(n3596), .C(n3597) );
  CKBD0 U3480 ( .CLK(n3597), .C(n3598) );
  CKBD0 U3481 ( .CLK(n3598), .C(n3599) );
  CKBD0 U3482 ( .CLK(n3599), .C(n3600) );
  CKBD0 U3483 ( .CLK(n3600), .C(n3601) );
  CKBD0 U3484 ( .CLK(n3601), .C(n3602) );
  CKBD0 U3485 ( .CLK(n3602), .C(n3603) );
  BUFFD0 U3486 ( .I(n3603), .Z(n3604) );
  CKBD0 U3487 ( .CLK(n3604), .C(n3605) );
  CKBD0 U3488 ( .CLK(n3605), .C(n3606) );
  CKBD0 U3489 ( .CLK(n3606), .C(n3607) );
  CKBD0 U3490 ( .CLK(n3607), .C(n3608) );
  CKBD0 U3491 ( .CLK(n3608), .C(n3609) );
  CKBD0 U3492 ( .CLK(n3609), .C(n3610) );
  CKBD0 U3493 ( .CLK(n3610), .C(n3611) );
  CKBD0 U3494 ( .CLK(n3611), .C(n3612) );
  CKBD0 U3495 ( .CLK(n3612), .C(n3613) );
  BUFFD0 U3496 ( .I(n3613), .Z(n3614) );
  CKBD0 U3497 ( .CLK(n3614), .C(n3615) );
  CKBD0 U3498 ( .CLK(n3615), .C(n3616) );
  CKBD0 U3499 ( .CLK(n3616), .C(n3617) );
  CKBD0 U3500 ( .CLK(n3617), .C(n3618) );
  CKBD0 U3501 ( .CLK(n3618), .C(n3619) );
  CKBD0 U3502 ( .CLK(n3619), .C(n3620) );
  CKBD0 U3503 ( .CLK(n3620), .C(n3621) );
  CKBD0 U3504 ( .CLK(n3621), .C(n3622) );
  CKBD0 U3505 ( .CLK(n3622), .C(n3623) );
  CKBD0 U3506 ( .CLK(n3623), .C(n3624) );
  CKBD0 U3507 ( .CLK(n3624), .C(n3625) );
  BUFFD0 U3508 ( .I(n3625), .Z(n3626) );
  CKBD0 U3509 ( .CLK(n3626), .C(n3627) );
  CKBD0 U3510 ( .CLK(n3627), .C(n3628) );
  CKBD0 U3511 ( .CLK(n3628), .C(n3629) );
  CKBD0 U3512 ( .CLK(n3629), .C(n3630) );
  CKBD0 U3513 ( .CLK(n3630), .C(n3631) );
  CKBD0 U3514 ( .CLK(n3631), .C(n3632) );
  CKBD0 U3515 ( .CLK(n3632), .C(n3633) );
  CKBD0 U3516 ( .CLK(n3633), .C(n3634) );
  CKBD0 U3517 ( .CLK(n3634), .C(n3635) );
  BUFFD0 U3518 ( .I(n3635), .Z(n3636) );
  CKBD0 U3519 ( .CLK(n3636), .C(n3637) );
  CKBD0 U3520 ( .CLK(n3637), .C(n3638) );
  CKBD0 U3521 ( .CLK(n3638), .C(n3639) );
  CKBD0 U3522 ( .CLK(n3639), .C(n3640) );
  CKBD0 U3523 ( .CLK(n3640), .C(n3641) );
  CKBD0 U3524 ( .CLK(n3641), .C(n3642) );
  CKBD0 U3525 ( .CLK(n3642), .C(n3643) );
  CKBD0 U3526 ( .CLK(n3643), .C(n3644) );
  CKBD0 U3527 ( .CLK(n3644), .C(n3645) );
  CKBD0 U3528 ( .CLK(n3645), .C(n3646) );
  BUFFD0 U3529 ( .I(n3646), .Z(n3647) );
  CKBD0 U3530 ( .CLK(n3647), .C(n3648) );
  CKBD0 U3531 ( .CLK(n3648), .C(n3649) );
  CKBD0 U3532 ( .CLK(n3649), .C(n3650) );
  CKBD0 U3533 ( .CLK(n3650), .C(n3651) );
  CKBD0 U3534 ( .CLK(n3651), .C(n3652) );
  CKBD0 U3535 ( .CLK(n3652), .C(n3653) );
  CKBD0 U3536 ( .CLK(n3653), .C(n3654) );
  CKBD0 U3537 ( .CLK(n3654), .C(n3655) );
  CKBD0 U3538 ( .CLK(n3655), .C(n3656) );
  CKBD0 U3539 ( .CLK(n3656), .C(n3657) );
  CKBD0 U3540 ( .CLK(n3657), .C(n3658) );
  BUFFD0 U3541 ( .I(n3658), .Z(n3659) );
  CKBD0 U3542 ( .CLK(n3659), .C(n3660) );
  CKBD0 U3543 ( .CLK(n3660), .C(n3661) );
  CKBD0 U3544 ( .CLK(n3661), .C(n3662) );
  CKBD0 U3545 ( .CLK(n3662), .C(n3663) );
  CKBD0 U3546 ( .CLK(n3663), .C(n3664) );
  CKBD0 U3547 ( .CLK(n3664), .C(n3665) );
  CKBD0 U3548 ( .CLK(n3665), .C(n3666) );
  CKBD0 U3549 ( .CLK(n3666), .C(n3667) );
  CKBD0 U3550 ( .CLK(n3667), .C(n3668) );
  BUFFD0 U3551 ( .I(n3668), .Z(n3669) );
  CKBD0 U3552 ( .CLK(n3669), .C(n3670) );
  CKBD0 U3553 ( .CLK(n3670), .C(n3671) );
  CKBD0 U3554 ( .CLK(n3671), .C(n3672) );
  CKBD0 U3555 ( .CLK(n3672), .C(n3673) );
  CKBD0 U3556 ( .CLK(n3673), .C(n3674) );
  CKBD0 U3557 ( .CLK(n3674), .C(n3675) );
  CKBD0 U3558 ( .CLK(n3675), .C(n3676) );
  CKBD0 U3559 ( .CLK(n3676), .C(n3677) );
  CKBD0 U3560 ( .CLK(n3677), .C(n3678) );
  CKBD0 U3561 ( .CLK(n3678), .C(n3679) );
  CKBD0 U3562 ( .CLK(n3679), .C(n3680) );
  BUFFD0 U3563 ( .I(n3680), .Z(n3681) );
  CKBD0 U3564 ( .CLK(n3681), .C(n3682) );
  CKBD0 U3565 ( .CLK(n3682), .C(n3683) );
  CKBD0 U3566 ( .CLK(n3683), .C(n3684) );
  CKBD0 U3567 ( .CLK(n3684), .C(n3685) );
  CKBD0 U3568 ( .CLK(n3685), .C(n3686) );
  CKBD0 U3569 ( .CLK(n3686), .C(n3687) );
  CKBD0 U3570 ( .CLK(n3687), .C(n3688) );
  CKBD0 U3571 ( .CLK(n3688), .C(n3689) );
  CKBD0 U3572 ( .CLK(n3689), .C(n3690) );
  BUFFD0 U3573 ( .I(n3690), .Z(n3691) );
  CKBD0 U3574 ( .CLK(n3691), .C(n3692) );
  CKBD0 U3575 ( .CLK(n3692), .C(n3693) );
  CKBD0 U3576 ( .CLK(n3693), .C(n3694) );
  CKBD0 U3577 ( .CLK(n3694), .C(n3695) );
  CKBD0 U3578 ( .CLK(n3695), .C(n3696) );
  CKBD0 U3579 ( .CLK(n3696), .C(n3697) );
  CKBD0 U3580 ( .CLK(n3697), .C(n3698) );
  CKBD0 U3581 ( .CLK(n3698), .C(n3699) );
  CKBD0 U3582 ( .CLK(n3699), .C(n3700) );
  BUFFD0 U3583 ( .I(n3700), .Z(n3701) );
  CKBD0 U3584 ( .CLK(n3701), .C(n3702) );
  CKBD0 U3585 ( .CLK(n3702), .C(n3703) );
  CKBD0 U3586 ( .CLK(n3703), .C(n3704) );
  CKBD0 U3587 ( .CLK(n3704), .C(n3705) );
  CKBD0 U3588 ( .CLK(n3705), .C(n3706) );
  CKBD0 U3589 ( .CLK(n3706), .C(n3707) );
  BUFFD0 U3590 ( .I(n3707), .Z(n3708) );
  CKBD0 U3591 ( .CLK(n3708), .C(n3709) );
  BUFFD0 U3592 ( .I(n3709), .Z(n3710) );
  CKBD0 U3593 ( .CLK(n3710), .C(n3711) );
  BUFFD0 U3594 ( .I(n3711), .Z(n3712) );
  CKBD0 U3595 ( .CLK(n3712), .C(n3713) );
  BUFFD0 U3596 ( .I(n3713), .Z(n3714) );
  CKBD0 U3597 ( .CLK(n3714), .C(n3715) );
  BUFFD0 U3598 ( .I(n3715), .Z(n3716) );
  CKBD0 U3599 ( .CLK(n3716), .C(n3717) );
  BUFFD0 U3600 ( .I(n3717), .Z(n3718) );
  CKBD0 U3601 ( .CLK(n3718), .C(n3719) );
  BUFFD0 U3602 ( .I(n3719), .Z(n3720) );
  CKBD0 U3603 ( .CLK(n3720), .C(n3721) );
  BUFFD0 U3604 ( .I(n3721), .Z(n3722) );
  BUFFD0 U3605 ( .I(n3724), .Z(n3723) );
  BUFFD0 U3606 ( .I(n3725), .Z(n3724) );
  BUFFD0 U3607 ( .I(n154), .Z(n3725) );
  CKBD0 U3608 ( .CLK(n1165), .C(n3726) );
  CKBD0 U3609 ( .CLK(n3726), .C(n3727) );
  CKBD0 U3610 ( .CLK(n3727), .C(n3728) );
  BUFFD0 U3611 ( .I(n3728), .Z(n3729) );
  CKBD0 U3612 ( .CLK(n3729), .C(n3730) );
  CKBD0 U3613 ( .CLK(n3730), .C(n3731) );
  CKBD0 U3614 ( .CLK(n3731), .C(n3732) );
  CKBD0 U3615 ( .CLK(n3732), .C(n3733) );
  CKBD0 U3616 ( .CLK(n3733), .C(n3734) );
  CKBD0 U3617 ( .CLK(n3734), .C(n3735) );
  CKBD0 U3618 ( .CLK(n3735), .C(n3736) );
  CKBD0 U3619 ( .CLK(n3736), .C(n3737) );
  CKBD0 U3620 ( .CLK(n3737), .C(n3738) );
  CKBD0 U3621 ( .CLK(n3738), .C(n3739) );
  BUFFD0 U3622 ( .I(n3739), .Z(n3740) );
  CKBD0 U3623 ( .CLK(n3740), .C(n3741) );
  CKBD0 U3624 ( .CLK(n3741), .C(n3742) );
  CKBD0 U3625 ( .CLK(n3742), .C(n3743) );
  CKBD0 U3626 ( .CLK(n3743), .C(n3744) );
  CKBD0 U3627 ( .CLK(n3744), .C(n3745) );
  CKBD0 U3628 ( .CLK(n3745), .C(n3746) );
  CKBD0 U3629 ( .CLK(n3746), .C(n3747) );
  CKBD0 U3630 ( .CLK(n3747), .C(n3748) );
  CKBD0 U3631 ( .CLK(n3748), .C(n3749) );
  CKBD0 U3632 ( .CLK(n3749), .C(n3750) );
  BUFFD0 U3633 ( .I(n3750), .Z(n3751) );
  CKBD0 U3634 ( .CLK(n3751), .C(n3752) );
  CKBD0 U3635 ( .CLK(n3752), .C(n3753) );
  CKBD0 U3636 ( .CLK(n3753), .C(n3754) );
  CKBD0 U3637 ( .CLK(n3754), .C(n3755) );
  CKBD0 U3638 ( .CLK(n3755), .C(n3756) );
  CKBD0 U3639 ( .CLK(n3756), .C(n3757) );
  CKBD0 U3640 ( .CLK(n3757), .C(n3758) );
  CKBD0 U3641 ( .CLK(n3758), .C(n3759) );
  CKBD0 U3642 ( .CLK(n3759), .C(n3760) );
  CKBD0 U3643 ( .CLK(n3760), .C(n3761) );
  BUFFD0 U3644 ( .I(n3761), .Z(n3762) );
  CKBD0 U3645 ( .CLK(n3762), .C(n3763) );
  CKBD0 U3646 ( .CLK(n3763), .C(n3764) );
  CKBD0 U3647 ( .CLK(n3764), .C(n3765) );
  CKBD0 U3648 ( .CLK(n3765), .C(n3766) );
  CKBD0 U3649 ( .CLK(n3766), .C(n3767) );
  CKBD0 U3650 ( .CLK(n3767), .C(n3768) );
  CKBD0 U3651 ( .CLK(n3768), .C(n3769) );
  CKBD0 U3652 ( .CLK(n3769), .C(n3770) );
  CKBD0 U3653 ( .CLK(n3770), .C(n3771) );
  BUFFD0 U3654 ( .I(n3771), .Z(n3772) );
  CKBD0 U3655 ( .CLK(n3772), .C(n3773) );
  CKBD0 U3656 ( .CLK(n3773), .C(n3774) );
  CKBD0 U3657 ( .CLK(n3774), .C(n3775) );
  CKBD0 U3658 ( .CLK(n3775), .C(n3776) );
  CKBD0 U3659 ( .CLK(n3776), .C(n3777) );
  CKBD0 U3660 ( .CLK(n3777), .C(n3778) );
  CKBD0 U3661 ( .CLK(n3778), .C(n3779) );
  CKBD0 U3662 ( .CLK(n3779), .C(n3780) );
  CKBD0 U3663 ( .CLK(n3780), .C(n3781) );
  CKBD0 U3664 ( .CLK(n3781), .C(n3782) );
  CKBD0 U3665 ( .CLK(n3782), .C(n3783) );
  BUFFD0 U3666 ( .I(n3783), .Z(n3784) );
  CKBD0 U3667 ( .CLK(n3784), .C(n3785) );
  CKBD0 U3668 ( .CLK(n3785), .C(n3786) );
  CKBD0 U3669 ( .CLK(n3786), .C(n3787) );
  CKBD0 U3670 ( .CLK(n3787), .C(n3788) );
  CKBD0 U3671 ( .CLK(n3788), .C(n3789) );
  CKBD0 U3672 ( .CLK(n3789), .C(n3790) );
  CKBD0 U3673 ( .CLK(n3790), .C(n3791) );
  CKBD0 U3674 ( .CLK(n3791), .C(n3792) );
  CKBD0 U3675 ( .CLK(n3792), .C(n3793) );
  BUFFD0 U3676 ( .I(n3793), .Z(n3794) );
  CKBD0 U3677 ( .CLK(n3794), .C(n3795) );
  CKBD0 U3678 ( .CLK(n3795), .C(n3796) );
  CKBD0 U3679 ( .CLK(n3796), .C(n3797) );
  CKBD0 U3680 ( .CLK(n3797), .C(n3798) );
  CKBD0 U3681 ( .CLK(n3798), .C(n3799) );
  CKBD0 U3682 ( .CLK(n3799), .C(n3800) );
  CKBD0 U3683 ( .CLK(n3800), .C(n3801) );
  CKBD0 U3684 ( .CLK(n3801), .C(n3802) );
  CKBD0 U3685 ( .CLK(n3802), .C(n3803) );
  CKBD0 U3686 ( .CLK(n3803), .C(n3804) );
  BUFFD0 U3687 ( .I(n3804), .Z(n3805) );
  CKBD0 U3688 ( .CLK(n3805), .C(n3806) );
  CKBD0 U3689 ( .CLK(n3806), .C(n3807) );
  CKBD0 U3690 ( .CLK(n3807), .C(n3808) );
  CKBD0 U3691 ( .CLK(n3808), .C(n3809) );
  CKBD0 U3692 ( .CLK(n3809), .C(n3810) );
  CKBD0 U3693 ( .CLK(n3810), .C(n3811) );
  CKBD0 U3694 ( .CLK(n3811), .C(n3812) );
  CKBD0 U3695 ( .CLK(n3812), .C(n3813) );
  CKBD0 U3696 ( .CLK(n3813), .C(n3814) );
  CKBD0 U3697 ( .CLK(n3814), .C(n3815) );
  BUFFD0 U3698 ( .I(n3815), .Z(n3816) );
  CKBD0 U3699 ( .CLK(n3816), .C(n3817) );
  CKBD0 U3700 ( .CLK(n3817), .C(n3818) );
  CKBD0 U3701 ( .CLK(n3818), .C(n3819) );
  CKBD0 U3702 ( .CLK(n3819), .C(n3820) );
  CKBD0 U3703 ( .CLK(n3820), .C(n3821) );
  CKBD0 U3704 ( .CLK(n3821), .C(n3822) );
  CKBD0 U3705 ( .CLK(n3822), .C(n3823) );
  CKBD0 U3706 ( .CLK(n3823), .C(n3824) );
  CKBD0 U3707 ( .CLK(n3824), .C(n3825) );
  CKBD0 U3708 ( .CLK(n3825), .C(n3826) );
  BUFFD0 U3709 ( .I(n3826), .Z(n3827) );
  CKBD0 U3710 ( .CLK(n3827), .C(n3828) );
  CKBD0 U3711 ( .CLK(n3828), .C(n3829) );
  CKBD0 U3712 ( .CLK(n3829), .C(n3830) );
  CKBD0 U3713 ( .CLK(n3830), .C(n3831) );
  CKBD0 U3714 ( .CLK(n3831), .C(n3832) );
  CKBD0 U3715 ( .CLK(n3832), .C(n3833) );
  CKBD0 U3716 ( .CLK(n3833), .C(n3834) );
  CKBD0 U3717 ( .CLK(n3834), .C(n3835) );
  CKBD0 U3718 ( .CLK(n3835), .C(n3836) );
  BUFFD0 U3719 ( .I(n3836), .Z(n3837) );
  CKBD0 U3720 ( .CLK(n3837), .C(n3838) );
  CKBD0 U3721 ( .CLK(n3838), .C(n3839) );
  CKBD0 U3722 ( .CLK(n3839), .C(n3840) );
  CKBD0 U3723 ( .CLK(n3840), .C(n3841) );
  CKBD0 U3724 ( .CLK(n3841), .C(n3842) );
  CKBD0 U3725 ( .CLK(n3842), .C(n3843) );
  BUFFD0 U3726 ( .I(n3843), .Z(n3844) );
  CKBD0 U3727 ( .CLK(n3844), .C(n3845) );
  BUFFD0 U3728 ( .I(n3845), .Z(n3846) );
  CKBD0 U3729 ( .CLK(n3846), .C(n3847) );
  BUFFD0 U3730 ( .I(n3847), .Z(n3848) );
  CKBD0 U3731 ( .CLK(n3848), .C(n3849) );
  BUFFD0 U3732 ( .I(n3849), .Z(n3850) );
  CKBD0 U3733 ( .CLK(n3850), .C(n3851) );
  BUFFD0 U3734 ( .I(n3851), .Z(n3852) );
  CKBD0 U3735 ( .CLK(n3852), .C(n3853) );
  BUFFD0 U3736 ( .I(n3853), .Z(n3854) );
  CKBD0 U3737 ( .CLK(n3854), .C(n3855) );
  BUFFD0 U3738 ( .I(n3855), .Z(n3856) );
  CKBD0 U3739 ( .CLK(n3856), .C(n3857) );
  BUFFD0 U3740 ( .I(n3857), .Z(n3858) );
  BUFFD0 U3741 ( .I(n3860), .Z(n3859) );
  BUFFD0 U3742 ( .I(n3861), .Z(n3860) );
  BUFFD0 U3743 ( .I(n153), .Z(n3861) );
  CKBD0 U3744 ( .CLK(n1163), .C(n3862) );
  CKBD0 U3745 ( .CLK(n3862), .C(n3863) );
  CKBD0 U3746 ( .CLK(n3863), .C(n3864) );
  BUFFD0 U3747 ( .I(n3864), .Z(n3865) );
  CKBD0 U3748 ( .CLK(n3865), .C(n3866) );
  CKBD0 U3749 ( .CLK(n3866), .C(n3867) );
  CKBD0 U3750 ( .CLK(n3867), .C(n3868) );
  CKBD0 U3751 ( .CLK(n3868), .C(n3869) );
  CKBD0 U3752 ( .CLK(n3869), .C(n3870) );
  CKBD0 U3753 ( .CLK(n3870), .C(n3871) );
  CKBD0 U3754 ( .CLK(n3871), .C(n3872) );
  CKBD0 U3755 ( .CLK(n3872), .C(n3873) );
  CKBD0 U3756 ( .CLK(n3873), .C(n3874) );
  CKBD0 U3757 ( .CLK(n3874), .C(n3875) );
  BUFFD0 U3758 ( .I(n3875), .Z(n3876) );
  CKBD0 U3759 ( .CLK(n3876), .C(n3877) );
  CKBD0 U3760 ( .CLK(n3877), .C(n3878) );
  CKBD0 U3761 ( .CLK(n3878), .C(n3879) );
  CKBD0 U3762 ( .CLK(n3879), .C(n3880) );
  CKBD0 U3763 ( .CLK(n3880), .C(n3881) );
  CKBD0 U3764 ( .CLK(n3881), .C(n3882) );
  CKBD0 U3765 ( .CLK(n3882), .C(n3883) );
  CKBD0 U3766 ( .CLK(n3883), .C(n3884) );
  CKBD0 U3767 ( .CLK(n3884), .C(n3885) );
  CKBD0 U3768 ( .CLK(n3885), .C(n3886) );
  BUFFD0 U3769 ( .I(n3886), .Z(n3887) );
  CKBD0 U3770 ( .CLK(n3887), .C(n3888) );
  CKBD0 U3771 ( .CLK(n3888), .C(n3889) );
  CKBD0 U3772 ( .CLK(n3889), .C(n3890) );
  CKBD0 U3773 ( .CLK(n3890), .C(n3891) );
  CKBD0 U3774 ( .CLK(n3891), .C(n3892) );
  CKBD0 U3775 ( .CLK(n3892), .C(n3893) );
  CKBD0 U3776 ( .CLK(n3893), .C(n3894) );
  CKBD0 U3777 ( .CLK(n3894), .C(n3895) );
  CKBD0 U3778 ( .CLK(n3895), .C(n3896) );
  CKBD0 U3779 ( .CLK(n3896), .C(n3897) );
  BUFFD0 U3780 ( .I(n3897), .Z(n3898) );
  CKBD0 U3781 ( .CLK(n3898), .C(n3899) );
  CKBD0 U3782 ( .CLK(n3899), .C(n3900) );
  CKBD0 U3783 ( .CLK(n3900), .C(n3901) );
  CKBD0 U3784 ( .CLK(n3901), .C(n3902) );
  CKBD0 U3785 ( .CLK(n3902), .C(n3903) );
  CKBD0 U3786 ( .CLK(n3903), .C(n3904) );
  CKBD0 U3787 ( .CLK(n3904), .C(n3905) );
  CKBD0 U3788 ( .CLK(n3905), .C(n3906) );
  CKBD0 U3789 ( .CLK(n3906), .C(n3907) );
  BUFFD0 U3790 ( .I(n3907), .Z(n3908) );
  CKBD0 U3791 ( .CLK(n3908), .C(n3909) );
  CKBD0 U3792 ( .CLK(n3909), .C(n3910) );
  CKBD0 U3793 ( .CLK(n3910), .C(n3911) );
  CKBD0 U3794 ( .CLK(n3911), .C(n3912) );
  CKBD0 U3795 ( .CLK(n3912), .C(n3913) );
  CKBD0 U3796 ( .CLK(n3913), .C(n3914) );
  CKBD0 U3797 ( .CLK(n3914), .C(n3915) );
  CKBD0 U3798 ( .CLK(n3915), .C(n3916) );
  CKBD0 U3799 ( .CLK(n3916), .C(n3917) );
  CKBD0 U3800 ( .CLK(n3917), .C(n3918) );
  CKBD0 U3801 ( .CLK(n3918), .C(n3919) );
  BUFFD0 U3802 ( .I(n3919), .Z(n3920) );
  CKBD0 U3803 ( .CLK(n3920), .C(n3921) );
  CKBD0 U3804 ( .CLK(n3921), .C(n3922) );
  CKBD0 U3805 ( .CLK(n3922), .C(n3923) );
  CKBD0 U3806 ( .CLK(n3923), .C(n3924) );
  CKBD0 U3807 ( .CLK(n3924), .C(n3925) );
  CKBD0 U3808 ( .CLK(n3925), .C(n3926) );
  CKBD0 U3809 ( .CLK(n3926), .C(n3927) );
  CKBD0 U3810 ( .CLK(n3927), .C(n3928) );
  CKBD0 U3811 ( .CLK(n3928), .C(n3929) );
  BUFFD0 U3812 ( .I(n3929), .Z(n3930) );
  CKBD0 U3813 ( .CLK(n3930), .C(n3931) );
  CKBD0 U3814 ( .CLK(n3931), .C(n3932) );
  CKBD0 U3815 ( .CLK(n3932), .C(n3933) );
  CKBD0 U3816 ( .CLK(n3933), .C(n3934) );
  CKBD0 U3817 ( .CLK(n3934), .C(n3935) );
  CKBD0 U3818 ( .CLK(n3935), .C(n3936) );
  CKBD0 U3819 ( .CLK(n3936), .C(n3937) );
  CKBD0 U3820 ( .CLK(n3937), .C(n3938) );
  CKBD0 U3821 ( .CLK(n3938), .C(n3939) );
  CKBD0 U3822 ( .CLK(n3939), .C(n3940) );
  BUFFD0 U3823 ( .I(n3940), .Z(n3941) );
  CKBD0 U3824 ( .CLK(n3941), .C(n3942) );
  CKBD0 U3825 ( .CLK(n3942), .C(n3943) );
  CKBD0 U3826 ( .CLK(n3943), .C(n3944) );
  CKBD0 U3827 ( .CLK(n3944), .C(n3945) );
  CKBD0 U3828 ( .CLK(n3945), .C(n3946) );
  CKBD0 U3829 ( .CLK(n3946), .C(n3947) );
  CKBD0 U3830 ( .CLK(n3947), .C(n3948) );
  CKBD0 U3831 ( .CLK(n3948), .C(n3949) );
  CKBD0 U3832 ( .CLK(n3949), .C(n3950) );
  CKBD0 U3833 ( .CLK(n3950), .C(n3951) );
  BUFFD0 U3834 ( .I(n3951), .Z(n3952) );
  CKBD0 U3835 ( .CLK(n3952), .C(n3953) );
  CKBD0 U3836 ( .CLK(n3953), .C(n3954) );
  CKBD0 U3837 ( .CLK(n3954), .C(n3955) );
  CKBD0 U3838 ( .CLK(n3955), .C(n3956) );
  CKBD0 U3839 ( .CLK(n3956), .C(n3957) );
  CKBD0 U3840 ( .CLK(n3957), .C(n3958) );
  CKBD0 U3841 ( .CLK(n3958), .C(n3959) );
  CKBD0 U3842 ( .CLK(n3959), .C(n3960) );
  CKBD0 U3843 ( .CLK(n3960), .C(n3961) );
  CKBD0 U3844 ( .CLK(n3961), .C(n3962) );
  BUFFD0 U3845 ( .I(n3962), .Z(n3963) );
  CKBD0 U3846 ( .CLK(n3963), .C(n3964) );
  CKBD0 U3847 ( .CLK(n3964), .C(n3965) );
  CKBD0 U3848 ( .CLK(n3965), .C(n3966) );
  CKBD0 U3849 ( .CLK(n3966), .C(n3967) );
  CKBD0 U3850 ( .CLK(n3967), .C(n3968) );
  CKBD0 U3851 ( .CLK(n3968), .C(n3969) );
  CKBD0 U3852 ( .CLK(n3969), .C(n3970) );
  CKBD0 U3853 ( .CLK(n3970), .C(n3971) );
  CKBD0 U3854 ( .CLK(n3971), .C(n3972) );
  CKBD0 U3855 ( .CLK(n3972), .C(n3973) );
  BUFFD0 U3856 ( .I(n3973), .Z(n3974) );
  CKBD0 U3857 ( .CLK(n3974), .C(n3975) );
  CKBD0 U3858 ( .CLK(n3975), .C(n3976) );
  CKBD0 U3859 ( .CLK(n3976), .C(n3977) );
  CKBD0 U3860 ( .CLK(n3977), .C(n3978) );
  CKBD0 U3861 ( .CLK(n3978), .C(n3979) );
  BUFFD0 U3862 ( .I(n3979), .Z(n3980) );
  CKBD0 U3863 ( .CLK(n3980), .C(n3981) );
  BUFFD0 U3864 ( .I(n3981), .Z(n3982) );
  CKBD0 U3865 ( .CLK(n3982), .C(n3983) );
  BUFFD0 U3866 ( .I(n3983), .Z(n3984) );
  CKBD0 U3867 ( .CLK(n3984), .C(n3985) );
  BUFFD0 U3868 ( .I(n3985), .Z(n3986) );
  CKBD0 U3869 ( .CLK(n3986), .C(n3987) );
  BUFFD0 U3870 ( .I(n3987), .Z(n3988) );
  CKBD0 U3871 ( .CLK(n3988), .C(n3989) );
  BUFFD0 U3872 ( .I(n3989), .Z(n3990) );
  CKBD0 U3873 ( .CLK(n3990), .C(n3991) );
  BUFFD0 U3874 ( .I(n3991), .Z(n3992) );
  CKBD0 U3875 ( .CLK(n3992), .C(n3993) );
  BUFFD0 U3876 ( .I(n3993), .Z(n3994) );
  BUFFD0 U3877 ( .I(n3996), .Z(n3995) );
  BUFFD0 U3878 ( .I(n3997), .Z(n3996) );
  BUFFD0 U3879 ( .I(n152), .Z(n3997) );
  CKBD0 U3880 ( .CLK(n1161), .C(n3998) );
  CKBD0 U3881 ( .CLK(n3998), .C(n3999) );
  CKBD0 U3882 ( .CLK(n3999), .C(n4000) );
  BUFFD0 U3883 ( .I(n4000), .Z(n4001) );
  CKBD0 U3884 ( .CLK(n4001), .C(n4002) );
  CKBD0 U3885 ( .CLK(n4002), .C(n4003) );
  CKBD0 U3886 ( .CLK(n4003), .C(n4004) );
  CKBD0 U3887 ( .CLK(n4004), .C(n4005) );
  CKBD0 U3888 ( .CLK(n4005), .C(n4006) );
  CKBD0 U3889 ( .CLK(n4006), .C(n4007) );
  CKBD0 U3890 ( .CLK(n4007), .C(n4008) );
  CKBD0 U3891 ( .CLK(n4008), .C(n4009) );
  CKBD0 U3892 ( .CLK(n4009), .C(n4010) );
  CKBD0 U3893 ( .CLK(n4010), .C(n4011) );
  CKBD0 U3894 ( .CLK(n4011), .C(n4012) );
  BUFFD0 U3895 ( .I(n4012), .Z(n4013) );
  CKBD0 U3896 ( .CLK(n4013), .C(n4014) );
  CKBD0 U3897 ( .CLK(n4014), .C(n4015) );
  CKBD0 U3898 ( .CLK(n4015), .C(n4016) );
  CKBD0 U3899 ( .CLK(n4016), .C(n4017) );
  CKBD0 U3900 ( .CLK(n4017), .C(n4018) );
  CKBD0 U3901 ( .CLK(n4018), .C(n4019) );
  CKBD0 U3902 ( .CLK(n4019), .C(n4020) );
  CKBD0 U3903 ( .CLK(n4020), .C(n4021) );
  CKBD0 U3904 ( .CLK(n4021), .C(n4022) );
  BUFFD0 U3905 ( .I(n4022), .Z(n4023) );
  CKBD0 U3906 ( .CLK(n4023), .C(n4024) );
  CKBD0 U3907 ( .CLK(n4024), .C(n4025) );
  CKBD0 U3908 ( .CLK(n4025), .C(n4026) );
  CKBD0 U3909 ( .CLK(n4026), .C(n4027) );
  CKBD0 U3910 ( .CLK(n4027), .C(n4028) );
  CKBD0 U3911 ( .CLK(n4028), .C(n4029) );
  CKBD0 U3912 ( .CLK(n4029), .C(n4030) );
  CKBD0 U3913 ( .CLK(n4030), .C(n4031) );
  CKBD0 U3914 ( .CLK(n4031), .C(n4032) );
  BUFFD0 U3915 ( .I(n4032), .Z(n4033) );
  CKBD0 U3916 ( .CLK(n4033), .C(n4034) );
  CKBD0 U3917 ( .CLK(n4034), .C(n4035) );
  CKBD0 U3918 ( .CLK(n4035), .C(n4036) );
  CKBD0 U3919 ( .CLK(n4036), .C(n4037) );
  CKBD0 U3920 ( .CLK(n4037), .C(n4038) );
  CKBD0 U3921 ( .CLK(n4038), .C(n4039) );
  CKBD0 U3922 ( .CLK(n4039), .C(n4040) );
  CKBD0 U3923 ( .CLK(n4040), .C(n4041) );
  CKBD0 U3924 ( .CLK(n4041), .C(n4042) );
  CKBD0 U3925 ( .CLK(n4042), .C(n4043) );
  CKBD0 U3926 ( .CLK(n4043), .C(n4044) );
  BUFFD0 U3927 ( .I(n4044), .Z(n4045) );
  CKBD0 U3928 ( .CLK(n4045), .C(n4046) );
  CKBD0 U3929 ( .CLK(n4046), .C(n4047) );
  CKBD0 U3930 ( .CLK(n4047), .C(n4048) );
  CKBD0 U3931 ( .CLK(n4048), .C(n4049) );
  CKBD0 U3932 ( .CLK(n4049), .C(n4050) );
  CKBD0 U3933 ( .CLK(n4050), .C(n4051) );
  CKBD0 U3934 ( .CLK(n4051), .C(n4052) );
  CKBD0 U3935 ( .CLK(n4052), .C(n4053) );
  CKBD0 U3936 ( .CLK(n4053), .C(n4054) );
  CKBD0 U3937 ( .CLK(n4054), .C(n4055) );
  BUFFD0 U3938 ( .I(n4055), .Z(n4056) );
  CKBD0 U3939 ( .CLK(n4056), .C(n4057) );
  CKBD0 U3940 ( .CLK(n4057), .C(n4058) );
  CKBD0 U3941 ( .CLK(n4058), .C(n4059) );
  CKBD0 U3942 ( .CLK(n4059), .C(n4060) );
  CKBD0 U3943 ( .CLK(n4060), .C(n4061) );
  CKBD0 U3944 ( .CLK(n4061), .C(n4062) );
  CKBD0 U3945 ( .CLK(n4062), .C(n4063) );
  CKBD0 U3946 ( .CLK(n4063), .C(n4064) );
  CKBD0 U3947 ( .CLK(n4064), .C(n4065) );
  BUFFD0 U3948 ( .I(n4065), .Z(n4066) );
  CKBD0 U3949 ( .CLK(n4066), .C(n4067) );
  CKBD0 U3950 ( .CLK(n4067), .C(n4068) );
  CKBD0 U3951 ( .CLK(n4068), .C(n4069) );
  CKBD0 U3952 ( .CLK(n4069), .C(n4070) );
  CKBD0 U3953 ( .CLK(n4070), .C(n4071) );
  CKBD0 U3954 ( .CLK(n4071), .C(n4072) );
  CKBD0 U3955 ( .CLK(n4072), .C(n4073) );
  CKBD0 U3956 ( .CLK(n4073), .C(n4074) );
  CKBD0 U3957 ( .CLK(n4074), .C(n4075) );
  CKBD0 U3958 ( .CLK(n4075), .C(n4076) );
  CKBD0 U3959 ( .CLK(n4076), .C(n4077) );
  BUFFD0 U3960 ( .I(n4077), .Z(n4078) );
  CKBD0 U3961 ( .CLK(n4078), .C(n4079) );
  CKBD0 U3962 ( .CLK(n4079), .C(n4080) );
  CKBD0 U3963 ( .CLK(n4080), .C(n4081) );
  CKBD0 U3964 ( .CLK(n4081), .C(n4082) );
  CKBD0 U3965 ( .CLK(n4082), .C(n4083) );
  CKBD0 U3966 ( .CLK(n4083), .C(n4084) );
  CKBD0 U3967 ( .CLK(n4084), .C(n4085) );
  CKBD0 U3968 ( .CLK(n4085), .C(n4086) );
  CKBD0 U3969 ( .CLK(n4086), .C(n4087) );
  BUFFD0 U3970 ( .I(n4087), .Z(n4088) );
  CKBD0 U3971 ( .CLK(n4088), .C(n4089) );
  CKBD0 U3972 ( .CLK(n4089), .C(n4090) );
  CKBD0 U3973 ( .CLK(n4090), .C(n4091) );
  CKBD0 U3974 ( .CLK(n4091), .C(n4092) );
  CKBD0 U3975 ( .CLK(n4092), .C(n4093) );
  CKBD0 U3976 ( .CLK(n4093), .C(n4094) );
  CKBD0 U3977 ( .CLK(n4094), .C(n4095) );
  CKBD0 U3978 ( .CLK(n4095), .C(n4096) );
  CKBD0 U3979 ( .CLK(n4096), .C(n4097) );
  BUFFD0 U3980 ( .I(n4097), .Z(n4098) );
  CKBD0 U3981 ( .CLK(n4098), .C(n4099) );
  CKBD0 U3982 ( .CLK(n4099), .C(n4100) );
  CKBD0 U3983 ( .CLK(n4100), .C(n4101) );
  CKBD0 U3984 ( .CLK(n4101), .C(n4102) );
  CKBD0 U3985 ( .CLK(n4102), .C(n4103) );
  CKBD0 U3986 ( .CLK(n4103), .C(n4104) );
  CKBD0 U3987 ( .CLK(n4104), .C(n4105) );
  CKBD0 U3988 ( .CLK(n4105), .C(n4106) );
  CKBD0 U3989 ( .CLK(n4106), .C(n4107) );
  CKBD0 U3990 ( .CLK(n4107), .C(n4108) );
  CKBD0 U3991 ( .CLK(n4108), .C(n4109) );
  BUFFD0 U3992 ( .I(n4109), .Z(n4110) );
  CKBD0 U3993 ( .CLK(n4110), .C(n4111) );
  CKBD0 U3994 ( .CLK(n4111), .C(n4112) );
  CKBD0 U3995 ( .CLK(n4112), .C(n4113) );
  CKBD0 U3996 ( .CLK(n4113), .C(n4114) );
  CKBD0 U3997 ( .CLK(n4114), .C(n4115) );
  BUFFD0 U3998 ( .I(n4115), .Z(n4116) );
  CKBD0 U3999 ( .CLK(n4116), .C(n4117) );
  BUFFD0 U4000 ( .I(n4117), .Z(n4118) );
  CKBD0 U4001 ( .CLK(n4118), .C(n4119) );
  BUFFD0 U4002 ( .I(n4119), .Z(n4120) );
  CKBD0 U4003 ( .CLK(n4120), .C(n4121) );
  BUFFD0 U4004 ( .I(n4121), .Z(n4122) );
  CKBD0 U4005 ( .CLK(n4122), .C(n4123) );
  BUFFD0 U4006 ( .I(n4123), .Z(n4124) );
  CKBD0 U4007 ( .CLK(n4124), .C(n4125) );
  BUFFD0 U4008 ( .I(n4125), .Z(n4126) );
  CKBD0 U4009 ( .CLK(n4126), .C(n4127) );
  BUFFD0 U4010 ( .I(n4127), .Z(n4128) );
  CKBD0 U4011 ( .CLK(n4128), .C(n4129) );
  BUFFD0 U4012 ( .I(n4129), .Z(n4130) );
  BUFFD0 U4013 ( .I(n4132), .Z(n4131) );
  BUFFD0 U4014 ( .I(n4133), .Z(n4132) );
  BUFFD0 U4015 ( .I(n151), .Z(n4133) );
  CKBD0 U4016 ( .CLK(n1159), .C(n4134) );
  CKBD0 U4017 ( .CLK(n4134), .C(n4135) );
  CKBD0 U4018 ( .CLK(n4135), .C(n4136) );
  BUFFD0 U4019 ( .I(n4136), .Z(n4137) );
  CKBD0 U4020 ( .CLK(n4137), .C(n4138) );
  CKBD0 U4021 ( .CLK(n4138), .C(n4139) );
  CKBD0 U4022 ( .CLK(n4139), .C(n4140) );
  CKBD0 U4023 ( .CLK(n4140), .C(n4141) );
  CKBD0 U4024 ( .CLK(n4141), .C(n4142) );
  CKBD0 U4025 ( .CLK(n4142), .C(n4143) );
  CKBD0 U4026 ( .CLK(n4143), .C(n4144) );
  CKBD0 U4027 ( .CLK(n4144), .C(n4145) );
  CKBD0 U4028 ( .CLK(n4145), .C(n4146) );
  CKBD0 U4029 ( .CLK(n4146), .C(n4147) );
  BUFFD0 U4030 ( .I(n4147), .Z(n4148) );
  CKBD0 U4031 ( .CLK(n4148), .C(n4149) );
  CKBD0 U4032 ( .CLK(n4149), .C(n4150) );
  CKBD0 U4033 ( .CLK(n4150), .C(n4151) );
  CKBD0 U4034 ( .CLK(n4151), .C(n4152) );
  CKBD0 U4035 ( .CLK(n4152), .C(n4153) );
  CKBD0 U4036 ( .CLK(n4153), .C(n4154) );
  CKBD0 U4037 ( .CLK(n4154), .C(n4155) );
  CKBD0 U4038 ( .CLK(n4155), .C(n4156) );
  CKBD0 U4039 ( .CLK(n4156), .C(n4157) );
  CKBD0 U4040 ( .CLK(n4157), .C(n4158) );
  BUFFD0 U4041 ( .I(n4158), .Z(n4159) );
  CKBD0 U4042 ( .CLK(n4159), .C(n4160) );
  CKBD0 U4043 ( .CLK(n4160), .C(n4161) );
  CKBD0 U4044 ( .CLK(n4161), .C(n4162) );
  CKBD0 U4045 ( .CLK(n4162), .C(n4163) );
  CKBD0 U4046 ( .CLK(n4163), .C(n4164) );
  CKBD0 U4047 ( .CLK(n4164), .C(n4165) );
  CKBD0 U4048 ( .CLK(n4165), .C(n4166) );
  CKBD0 U4049 ( .CLK(n4166), .C(n4167) );
  CKBD0 U4050 ( .CLK(n4167), .C(n4168) );
  BUFFD0 U4051 ( .I(n4168), .Z(n4169) );
  CKBD0 U4052 ( .CLK(n4169), .C(n4170) );
  CKBD0 U4053 ( .CLK(n4170), .C(n4171) );
  CKBD0 U4054 ( .CLK(n4171), .C(n4172) );
  CKBD0 U4055 ( .CLK(n4172), .C(n4173) );
  CKBD0 U4056 ( .CLK(n4173), .C(n4174) );
  CKBD0 U4057 ( .CLK(n4174), .C(n4175) );
  CKBD0 U4058 ( .CLK(n4175), .C(n4176) );
  CKBD0 U4059 ( .CLK(n4176), .C(n4177) );
  CKBD0 U4060 ( .CLK(n4177), .C(n4178) );
  CKBD0 U4061 ( .CLK(n4178), .C(n4179) );
  CKBD0 U4062 ( .CLK(n4179), .C(n4180) );
  BUFFD0 U4063 ( .I(n4180), .Z(n4181) );
  CKBD0 U4064 ( .CLK(n4181), .C(n4182) );
  CKBD0 U4065 ( .CLK(n4182), .C(n4183) );
  CKBD0 U4066 ( .CLK(n4183), .C(n4184) );
  CKBD0 U4067 ( .CLK(n4184), .C(n4185) );
  CKBD0 U4068 ( .CLK(n4185), .C(n4186) );
  CKBD0 U4069 ( .CLK(n4186), .C(n4187) );
  CKBD0 U4070 ( .CLK(n4187), .C(n4188) );
  CKBD0 U4071 ( .CLK(n4188), .C(n4189) );
  CKBD0 U4072 ( .CLK(n4189), .C(n4190) );
  BUFFD0 U4073 ( .I(n4190), .Z(n4191) );
  CKBD0 U4074 ( .CLK(n4191), .C(n4192) );
  CKBD0 U4075 ( .CLK(n4192), .C(n4193) );
  CKBD0 U4076 ( .CLK(n4193), .C(n4194) );
  CKBD0 U4077 ( .CLK(n4194), .C(n4195) );
  CKBD0 U4078 ( .CLK(n4195), .C(n4196) );
  CKBD0 U4079 ( .CLK(n4196), .C(n4197) );
  CKBD0 U4080 ( .CLK(n4197), .C(n4198) );
  CKBD0 U4081 ( .CLK(n4198), .C(n4199) );
  CKBD0 U4082 ( .CLK(n4199), .C(n4200) );
  CKBD0 U4083 ( .CLK(n4200), .C(n4201) );
  BUFFD0 U4084 ( .I(n4201), .Z(n4202) );
  CKBD0 U4085 ( .CLK(n4202), .C(n4203) );
  CKBD0 U4086 ( .CLK(n4203), .C(n4204) );
  CKBD0 U4087 ( .CLK(n4204), .C(n4205) );
  CKBD0 U4088 ( .CLK(n4205), .C(n4206) );
  CKBD0 U4089 ( .CLK(n4206), .C(n4207) );
  CKBD0 U4090 ( .CLK(n4207), .C(n4208) );
  CKBD0 U4091 ( .CLK(n4208), .C(n4209) );
  CKBD0 U4092 ( .CLK(n4209), .C(n4210) );
  CKBD0 U4093 ( .CLK(n4210), .C(n4211) );
  CKBD0 U4094 ( .CLK(n4211), .C(n4212) );
  BUFFD0 U4095 ( .I(n4212), .Z(n4213) );
  CKBD0 U4096 ( .CLK(n4213), .C(n4214) );
  CKBD0 U4097 ( .CLK(n4214), .C(n4215) );
  CKBD0 U4098 ( .CLK(n4215), .C(n4216) );
  CKBD0 U4099 ( .CLK(n4216), .C(n4217) );
  CKBD0 U4100 ( .CLK(n4217), .C(n4218) );
  CKBD0 U4101 ( .CLK(n4218), .C(n4219) );
  CKBD0 U4102 ( .CLK(n4219), .C(n4220) );
  CKBD0 U4103 ( .CLK(n4220), .C(n4221) );
  CKBD0 U4104 ( .CLK(n4221), .C(n4222) );
  CKBD0 U4105 ( .CLK(n4222), .C(n4223) );
  BUFFD0 U4106 ( .I(n4223), .Z(n4224) );
  CKBD0 U4107 ( .CLK(n4224), .C(n4225) );
  CKBD0 U4108 ( .CLK(n4225), .C(n4226) );
  CKBD0 U4109 ( .CLK(n4226), .C(n4227) );
  CKBD0 U4110 ( .CLK(n4227), .C(n4228) );
  CKBD0 U4111 ( .CLK(n4228), .C(n4229) );
  CKBD0 U4112 ( .CLK(n4229), .C(n4230) );
  CKBD0 U4113 ( .CLK(n4230), .C(n4231) );
  CKBD0 U4114 ( .CLK(n4231), .C(n4232) );
  CKBD0 U4115 ( .CLK(n4232), .C(n4233) );
  CKBD0 U4116 ( .CLK(n4233), .C(n4234) );
  BUFFD0 U4117 ( .I(n4234), .Z(n4235) );
  CKBD0 U4118 ( .CLK(n4235), .C(n4236) );
  CKBD0 U4119 ( .CLK(n4236), .C(n4237) );
  CKBD0 U4120 ( .CLK(n4237), .C(n4238) );
  CKBD0 U4121 ( .CLK(n4238), .C(n4239) );
  CKBD0 U4122 ( .CLK(n4239), .C(n4240) );
  CKBD0 U4123 ( .CLK(n4240), .C(n4241) );
  CKBD0 U4124 ( .CLK(n4241), .C(n4242) );
  CKBD0 U4125 ( .CLK(n4242), .C(n4243) );
  CKBD0 U4126 ( .CLK(n4243), .C(n4244) );
  CKBD0 U4127 ( .CLK(n4244), .C(n4245) );
  BUFFD0 U4128 ( .I(n4245), .Z(n4246) );
  CKBD0 U4129 ( .CLK(n4246), .C(n4247) );
  CKBD0 U4130 ( .CLK(n4247), .C(n4248) );
  CKBD0 U4131 ( .CLK(n4248), .C(n4249) );
  CKBD0 U4132 ( .CLK(n4249), .C(n4250) );
  CKBD0 U4133 ( .CLK(n4250), .C(n4251) );
  BUFFD0 U4134 ( .I(n4251), .Z(n4252) );
  CKBD0 U4135 ( .CLK(n4252), .C(n4253) );
  BUFFD0 U4136 ( .I(n4253), .Z(n4254) );
  CKBD0 U4137 ( .CLK(n4254), .C(n4255) );
  BUFFD0 U4138 ( .I(n4255), .Z(n4256) );
  CKBD0 U4139 ( .CLK(n4256), .C(n4257) );
  BUFFD0 U4140 ( .I(n4257), .Z(n4258) );
  CKBD0 U4141 ( .CLK(n4258), .C(n4259) );
  BUFFD0 U4142 ( .I(n4259), .Z(n4260) );
  CKBD0 U4143 ( .CLK(n4260), .C(n4261) );
  BUFFD0 U4144 ( .I(n4261), .Z(n4262) );
  CKBD0 U4145 ( .CLK(n4262), .C(n4263) );
  BUFFD0 U4146 ( .I(n4263), .Z(n4264) );
  CKBD0 U4147 ( .CLK(n4264), .C(n4265) );
  BUFFD0 U4148 ( .I(n4265), .Z(n4266) );
  BUFFD0 U4149 ( .I(n4268), .Z(n4267) );
  BUFFD0 U4150 ( .I(n4269), .Z(n4268) );
  BUFFD0 U4151 ( .I(n150), .Z(n4269) );
  CKBD0 U4152 ( .CLK(n1157), .C(n4270) );
  CKBD0 U4153 ( .CLK(n4270), .C(n4271) );
  CKBD0 U4154 ( .CLK(n4271), .C(n4272) );
  BUFFD0 U4155 ( .I(n4272), .Z(n4273) );
  CKBD0 U4156 ( .CLK(n4273), .C(n4274) );
  CKBD0 U4157 ( .CLK(n4274), .C(n4275) );
  CKBD0 U4158 ( .CLK(n4275), .C(n4276) );
  CKBD0 U4159 ( .CLK(n4276), .C(n4277) );
  CKBD0 U4160 ( .CLK(n4277), .C(n4278) );
  CKBD0 U4161 ( .CLK(n4278), .C(n4279) );
  CKBD0 U4162 ( .CLK(n4279), .C(n4280) );
  CKBD0 U4163 ( .CLK(n4280), .C(n4281) );
  CKBD0 U4164 ( .CLK(n4281), .C(n4282) );
  CKBD0 U4165 ( .CLK(n4282), .C(n4283) );
  BUFFD0 U4166 ( .I(n4283), .Z(n4284) );
  CKBD0 U4167 ( .CLK(n4284), .C(n4285) );
  CKBD0 U4168 ( .CLK(n4285), .C(n4286) );
  CKBD0 U4169 ( .CLK(n4286), .C(n4287) );
  CKBD0 U4170 ( .CLK(n4287), .C(n4288) );
  CKBD0 U4171 ( .CLK(n4288), .C(n4289) );
  CKBD0 U4172 ( .CLK(n4289), .C(n4290) );
  CKBD0 U4173 ( .CLK(n4290), .C(n4291) );
  CKBD0 U4174 ( .CLK(n4291), .C(n4292) );
  CKBD0 U4175 ( .CLK(n4292), .C(n4293) );
  CKBD0 U4176 ( .CLK(n4293), .C(n4294) );
  BUFFD0 U4177 ( .I(n4294), .Z(n4295) );
  CKBD0 U4178 ( .CLK(n4295), .C(n4296) );
  CKBD0 U4179 ( .CLK(n4296), .C(n4297) );
  CKBD0 U4180 ( .CLK(n4297), .C(n4298) );
  CKBD0 U4181 ( .CLK(n4298), .C(n4299) );
  CKBD0 U4182 ( .CLK(n4299), .C(n4300) );
  CKBD0 U4183 ( .CLK(n4300), .C(n4301) );
  CKBD0 U4184 ( .CLK(n4301), .C(n4302) );
  CKBD0 U4185 ( .CLK(n4302), .C(n4303) );
  CKBD0 U4186 ( .CLK(n4303), .C(n4304) );
  CKBD0 U4187 ( .CLK(n4304), .C(n4305) );
  BUFFD0 U4188 ( .I(n4305), .Z(n4306) );
  CKBD0 U4189 ( .CLK(n4306), .C(n4307) );
  CKBD0 U4190 ( .CLK(n4307), .C(n4308) );
  CKBD0 U4191 ( .CLK(n4308), .C(n4309) );
  CKBD0 U4192 ( .CLK(n4309), .C(n4310) );
  CKBD0 U4193 ( .CLK(n4310), .C(n4311) );
  CKBD0 U4194 ( .CLK(n4311), .C(n4312) );
  CKBD0 U4195 ( .CLK(n4312), .C(n4313) );
  CKBD0 U4196 ( .CLK(n4313), .C(n4314) );
  CKBD0 U4197 ( .CLK(n4314), .C(n4315) );
  CKBD0 U4198 ( .CLK(n4315), .C(n4316) );
  BUFFD0 U4199 ( .I(n4316), .Z(n4317) );
  CKBD0 U4200 ( .CLK(n4317), .C(n4318) );
  CKBD0 U4201 ( .CLK(n4318), .C(n4319) );
  CKBD0 U4202 ( .CLK(n4319), .C(n4320) );
  CKBD0 U4203 ( .CLK(n4320), .C(n4321) );
  CKBD0 U4204 ( .CLK(n4321), .C(n4322) );
  CKBD0 U4205 ( .CLK(n4322), .C(n4323) );
  CKBD0 U4206 ( .CLK(n4323), .C(n4324) );
  CKBD0 U4207 ( .CLK(n4324), .C(n4325) );
  CKBD0 U4208 ( .CLK(n4325), .C(n4326) );
  BUFFD0 U4209 ( .I(n4326), .Z(n4327) );
  CKBD0 U4210 ( .CLK(n4327), .C(n4328) );
  CKBD0 U4211 ( .CLK(n4328), .C(n4329) );
  CKBD0 U4212 ( .CLK(n4329), .C(n4330) );
  CKBD0 U4213 ( .CLK(n4330), .C(n4331) );
  CKBD0 U4214 ( .CLK(n4331), .C(n4332) );
  CKBD0 U4215 ( .CLK(n4332), .C(n4333) );
  CKBD0 U4216 ( .CLK(n4333), .C(n4334) );
  CKBD0 U4217 ( .CLK(n4334), .C(n4335) );
  CKBD0 U4218 ( .CLK(n4335), .C(n4336) );
  CKBD0 U4219 ( .CLK(n4336), .C(n4337) );
  CKBD0 U4220 ( .CLK(n4337), .C(n4338) );
  BUFFD0 U4221 ( .I(n4338), .Z(n4339) );
  CKBD0 U4222 ( .CLK(n4339), .C(n4340) );
  CKBD0 U4223 ( .CLK(n4340), .C(n4341) );
  CKBD0 U4224 ( .CLK(n4341), .C(n4342) );
  CKBD0 U4225 ( .CLK(n4342), .C(n4343) );
  CKBD0 U4226 ( .CLK(n4343), .C(n4344) );
  CKBD0 U4227 ( .CLK(n4344), .C(n4345) );
  CKBD0 U4228 ( .CLK(n4345), .C(n4346) );
  CKBD0 U4229 ( .CLK(n4346), .C(n4347) );
  CKBD0 U4230 ( .CLK(n4347), .C(n4348) );
  BUFFD0 U4231 ( .I(n4348), .Z(n4349) );
  CKBD0 U4232 ( .CLK(n4349), .C(n4350) );
  CKBD0 U4233 ( .CLK(n4350), .C(n4351) );
  CKBD0 U4234 ( .CLK(n4351), .C(n4352) );
  CKBD0 U4235 ( .CLK(n4352), .C(n4353) );
  CKBD0 U4236 ( .CLK(n4353), .C(n4354) );
  CKBD0 U4237 ( .CLK(n4354), .C(n4355) );
  CKBD0 U4238 ( .CLK(n4355), .C(n4356) );
  CKBD0 U4239 ( .CLK(n4356), .C(n4357) );
  CKBD0 U4240 ( .CLK(n4357), .C(n4358) );
  CKBD0 U4241 ( .CLK(n4358), .C(n4359) );
  BUFFD0 U4242 ( .I(n4359), .Z(n4360) );
  CKBD0 U4243 ( .CLK(n4360), .C(n4361) );
  CKBD0 U4244 ( .CLK(n4361), .C(n4362) );
  CKBD0 U4245 ( .CLK(n4362), .C(n4363) );
  CKBD0 U4246 ( .CLK(n4363), .C(n4364) );
  CKBD0 U4247 ( .CLK(n4364), .C(n4365) );
  CKBD0 U4248 ( .CLK(n4365), .C(n4366) );
  CKBD0 U4249 ( .CLK(n4366), .C(n4367) );
  CKBD0 U4250 ( .CLK(n4367), .C(n4368) );
  CKBD0 U4251 ( .CLK(n4368), .C(n4369) );
  CKBD0 U4252 ( .CLK(n4369), .C(n4370) );
  BUFFD0 U4253 ( .I(n4370), .Z(n4371) );
  CKBD0 U4254 ( .CLK(n4371), .C(n4372) );
  CKBD0 U4255 ( .CLK(n4372), .C(n4373) );
  CKBD0 U4256 ( .CLK(n4373), .C(n4374) );
  CKBD0 U4257 ( .CLK(n4374), .C(n4375) );
  CKBD0 U4258 ( .CLK(n4375), .C(n4376) );
  CKBD0 U4259 ( .CLK(n4376), .C(n4377) );
  CKBD0 U4260 ( .CLK(n4377), .C(n4378) );
  CKBD0 U4261 ( .CLK(n4378), .C(n4379) );
  CKBD0 U4262 ( .CLK(n4379), .C(n4380) );
  CKBD0 U4263 ( .CLK(n4380), .C(n4381) );
  BUFFD0 U4264 ( .I(n4381), .Z(n4382) );
  CKBD0 U4265 ( .CLK(n4382), .C(n4383) );
  CKBD0 U4266 ( .CLK(n4383), .C(n4384) );
  CKBD0 U4267 ( .CLK(n4384), .C(n4385) );
  CKBD0 U4268 ( .CLK(n4385), .C(n4386) );
  CKBD0 U4269 ( .CLK(n4386), .C(n4387) );
  BUFFD0 U4270 ( .I(n4387), .Z(n4388) );
  CKBD0 U4271 ( .CLK(n4388), .C(n4389) );
  BUFFD0 U4272 ( .I(n4389), .Z(n4390) );
  CKBD0 U4273 ( .CLK(n4390), .C(n4391) );
  BUFFD0 U4274 ( .I(n4391), .Z(n4392) );
  CKBD0 U4275 ( .CLK(n4392), .C(n4393) );
  BUFFD0 U4276 ( .I(n4393), .Z(n4394) );
  CKBD0 U4277 ( .CLK(n4394), .C(n4395) );
  BUFFD0 U4278 ( .I(n4395), .Z(n4396) );
  CKBD0 U4279 ( .CLK(n4396), .C(n4397) );
  BUFFD0 U4280 ( .I(n4397), .Z(n4398) );
  CKBD0 U4281 ( .CLK(n4398), .C(n4399) );
  BUFFD0 U4282 ( .I(n4399), .Z(n4400) );
  CKBD0 U4283 ( .CLK(n4400), .C(n4401) );
  BUFFD0 U4284 ( .I(n4401), .Z(n4402) );
  BUFFD0 U4285 ( .I(n4404), .Z(n4403) );
  BUFFD0 U4286 ( .I(n4405), .Z(n4404) );
  BUFFD0 U4287 ( .I(n149), .Z(n4405) );
  CKBD0 U4288 ( .CLK(n1155), .C(n4406) );
  CKBD0 U4289 ( .CLK(n4406), .C(n4407) );
  CKBD0 U4290 ( .CLK(n4407), .C(n4408) );
  CKBD0 U4291 ( .CLK(n4408), .C(n4409) );
  BUFFD0 U4292 ( .I(n4409), .Z(n4410) );
  CKBD0 U4293 ( .CLK(n4410), .C(n4411) );
  CKBD0 U4294 ( .CLK(n4411), .C(n4412) );
  CKBD0 U4295 ( .CLK(n4412), .C(n4413) );
  CKBD0 U4296 ( .CLK(n4413), .C(n4414) );
  CKBD0 U4297 ( .CLK(n4414), .C(n4415) );
  CKBD0 U4298 ( .CLK(n4415), .C(n4416) );
  CKBD0 U4299 ( .CLK(n4416), .C(n4417) );
  CKBD0 U4300 ( .CLK(n4417), .C(n4418) );
  CKBD0 U4301 ( .CLK(n4418), .C(n4419) );
  BUFFD0 U4302 ( .I(n4419), .Z(n4420) );
  CKBD0 U4303 ( .CLK(n4420), .C(n4421) );
  CKBD0 U4304 ( .CLK(n4421), .C(n4422) );
  CKBD0 U4305 ( .CLK(n4422), .C(n4423) );
  CKBD0 U4306 ( .CLK(n4423), .C(n4424) );
  CKBD0 U4307 ( .CLK(n4424), .C(n4425) );
  CKBD0 U4308 ( .CLK(n4425), .C(n4426) );
  CKBD0 U4309 ( .CLK(n4426), .C(n4427) );
  CKBD0 U4310 ( .CLK(n4427), .C(n4428) );
  CKBD0 U4311 ( .CLK(n4428), .C(n4429) );
  BUFFD0 U4312 ( .I(n4429), .Z(n4430) );
  CKBD0 U4313 ( .CLK(n4430), .C(n4431) );
  CKBD0 U4314 ( .CLK(n4431), .C(n4432) );
  CKBD0 U4315 ( .CLK(n4432), .C(n4433) );
  CKBD0 U4316 ( .CLK(n4433), .C(n4434) );
  CKBD0 U4317 ( .CLK(n4434), .C(n4435) );
  CKBD0 U4318 ( .CLK(n4435), .C(n4436) );
  CKBD0 U4319 ( .CLK(n4436), .C(n4437) );
  CKBD0 U4320 ( .CLK(n4437), .C(n4438) );
  CKBD0 U4321 ( .CLK(n4438), .C(n4439) );
  CKBD0 U4322 ( .CLK(n4439), .C(n4440) );
  CKBD0 U4323 ( .CLK(n4440), .C(n4441) );
  BUFFD0 U4324 ( .I(n4441), .Z(n4442) );
  CKBD0 U4325 ( .CLK(n4442), .C(n4443) );
  CKBD0 U4326 ( .CLK(n4443), .C(n4444) );
  CKBD0 U4327 ( .CLK(n4444), .C(n4445) );
  CKBD0 U4328 ( .CLK(n4445), .C(n4446) );
  CKBD0 U4329 ( .CLK(n4446), .C(n4447) );
  CKBD0 U4330 ( .CLK(n4447), .C(n4448) );
  CKBD0 U4331 ( .CLK(n4448), .C(n4449) );
  CKBD0 U4332 ( .CLK(n4449), .C(n4450) );
  CKBD0 U4333 ( .CLK(n4450), .C(n4451) );
  CKBD0 U4334 ( .CLK(n4451), .C(n4452) );
  BUFFD0 U4335 ( .I(n4452), .Z(n4453) );
  CKBD0 U4336 ( .CLK(n4453), .C(n4454) );
  CKBD0 U4337 ( .CLK(n4454), .C(n4455) );
  CKBD0 U4338 ( .CLK(n4455), .C(n4456) );
  CKBD0 U4339 ( .CLK(n4456), .C(n4457) );
  CKBD0 U4340 ( .CLK(n4457), .C(n4458) );
  CKBD0 U4341 ( .CLK(n4458), .C(n4459) );
  CKBD0 U4342 ( .CLK(n4459), .C(n4460) );
  CKBD0 U4343 ( .CLK(n4460), .C(n4461) );
  CKBD0 U4344 ( .CLK(n4461), .C(n4462) );
  BUFFD0 U4345 ( .I(n4462), .Z(n4463) );
  CKBD0 U4346 ( .CLK(n4463), .C(n4464) );
  CKBD0 U4347 ( .CLK(n4464), .C(n4465) );
  CKBD0 U4348 ( .CLK(n4465), .C(n4466) );
  CKBD0 U4349 ( .CLK(n4466), .C(n4467) );
  CKBD0 U4350 ( .CLK(n4467), .C(n4468) );
  CKBD0 U4351 ( .CLK(n4468), .C(n4469) );
  CKBD0 U4352 ( .CLK(n4469), .C(n4470) );
  CKBD0 U4353 ( .CLK(n4470), .C(n4471) );
  CKBD0 U4354 ( .CLK(n4471), .C(n4472) );
  CKBD0 U4355 ( .CLK(n4472), .C(n4473) );
  CKBD0 U4356 ( .CLK(n4473), .C(n4474) );
  BUFFD0 U4357 ( .I(n4474), .Z(n4475) );
  CKBD0 U4358 ( .CLK(n4475), .C(n4476) );
  CKBD0 U4359 ( .CLK(n4476), .C(n4477) );
  CKBD0 U4360 ( .CLK(n4477), .C(n4478) );
  CKBD0 U4361 ( .CLK(n4478), .C(n4479) );
  CKBD0 U4362 ( .CLK(n4479), .C(n4480) );
  CKBD0 U4363 ( .CLK(n4480), .C(n4481) );
  CKBD0 U4364 ( .CLK(n4481), .C(n4482) );
  CKBD0 U4365 ( .CLK(n4482), .C(n4483) );
  CKBD0 U4366 ( .CLK(n4483), .C(n4484) );
  BUFFD0 U4367 ( .I(n4484), .Z(n4485) );
  CKBD0 U4368 ( .CLK(n4485), .C(n4486) );
  CKBD0 U4369 ( .CLK(n4486), .C(n4487) );
  CKBD0 U4370 ( .CLK(n4487), .C(n4488) );
  CKBD0 U4371 ( .CLK(n4488), .C(n4489) );
  CKBD0 U4372 ( .CLK(n4489), .C(n4490) );
  CKBD0 U4373 ( .CLK(n4490), .C(n4491) );
  CKBD0 U4374 ( .CLK(n4491), .C(n4492) );
  CKBD0 U4375 ( .CLK(n4492), .C(n4493) );
  CKBD0 U4376 ( .CLK(n4493), .C(n4494) );
  CKBD0 U4377 ( .CLK(n4494), .C(n4495) );
  BUFFD0 U4378 ( .I(n4495), .Z(n4496) );
  CKBD0 U4379 ( .CLK(n4496), .C(n4497) );
  CKBD0 U4380 ( .CLK(n4497), .C(n4498) );
  CKBD0 U4381 ( .CLK(n4498), .C(n4499) );
  CKBD0 U4382 ( .CLK(n4499), .C(n4500) );
  CKBD0 U4383 ( .CLK(n4500), .C(n4501) );
  CKBD0 U4384 ( .CLK(n4501), .C(n4502) );
  CKBD0 U4385 ( .CLK(n4502), .C(n4503) );
  CKBD0 U4386 ( .CLK(n4503), .C(n4504) );
  CKBD0 U4387 ( .CLK(n4504), .C(n4505) );
  CKBD0 U4388 ( .CLK(n4505), .C(n4506) );
  BUFFD0 U4389 ( .I(n4506), .Z(n4507) );
  CKBD0 U4390 ( .CLK(n4507), .C(n4508) );
  CKBD0 U4391 ( .CLK(n4508), .C(n4509) );
  CKBD0 U4392 ( .CLK(n4509), .C(n4510) );
  CKBD0 U4393 ( .CLK(n4510), .C(n4511) );
  CKBD0 U4394 ( .CLK(n4511), .C(n4512) );
  CKBD0 U4395 ( .CLK(n4512), .C(n4513) );
  CKBD0 U4396 ( .CLK(n4513), .C(n4514) );
  CKBD0 U4397 ( .CLK(n4514), .C(n4515) );
  CKBD0 U4398 ( .CLK(n4515), .C(n4516) );
  BUFFD0 U4399 ( .I(n4516), .Z(n4517) );
  CKBD0 U4400 ( .CLK(n4517), .C(n4518) );
  CKBD0 U4401 ( .CLK(n4518), .C(n4519) );
  CKBD0 U4402 ( .CLK(n4519), .C(n4520) );
  CKBD0 U4403 ( .CLK(n4520), .C(n4521) );
  CKBD0 U4404 ( .CLK(n4521), .C(n4522) );
  CKBD0 U4405 ( .CLK(n4522), .C(n4523) );
  BUFFD0 U4406 ( .I(n4523), .Z(n4524) );
  CKBD0 U4407 ( .CLK(n4524), .C(n4525) );
  BUFFD0 U4408 ( .I(n4525), .Z(n4526) );
  CKBD0 U4409 ( .CLK(n4526), .C(n4527) );
  BUFFD0 U4410 ( .I(n4527), .Z(n4528) );
  CKBD0 U4411 ( .CLK(n4528), .C(n4529) );
  BUFFD0 U4412 ( .I(n4529), .Z(n4530) );
  CKBD0 U4413 ( .CLK(n4530), .C(n4531) );
  BUFFD0 U4414 ( .I(n4531), .Z(n4532) );
  CKBD0 U4415 ( .CLK(n4532), .C(n4533) );
  BUFFD0 U4416 ( .I(n4533), .Z(n4534) );
  CKBD0 U4417 ( .CLK(n4534), .C(n4535) );
  BUFFD0 U4418 ( .I(n4535), .Z(n4536) );
  CKBD0 U4419 ( .CLK(n4536), .C(n4537) );
  BUFFD0 U4420 ( .I(n4537), .Z(n4538) );
  BUFFD0 U4421 ( .I(n4540), .Z(n4539) );
  BUFFD0 U4422 ( .I(n4541), .Z(n4540) );
  BUFFD0 U4423 ( .I(n148), .Z(n4541) );
  CKBD0 U4424 ( .CLK(n672), .C(n4542) );
  CKBD0 U4425 ( .CLK(n4542), .C(n4543) );
  CKBD0 U4426 ( .CLK(n4543), .C(n4544) );
  BUFFD0 U4427 ( .I(n4544), .Z(n4545) );
  CKBD0 U4428 ( .CLK(n4545), .C(n4546) );
  CKBD0 U4429 ( .CLK(n4546), .C(n4547) );
  CKBD0 U4430 ( .CLK(n4547), .C(n4548) );
  CKBD0 U4431 ( .CLK(n4548), .C(n4549) );
  CKBD0 U4432 ( .CLK(n4549), .C(n4550) );
  CKBD0 U4433 ( .CLK(n4550), .C(n4551) );
  CKBD0 U4434 ( .CLK(n4551), .C(n4552) );
  CKBD0 U4435 ( .CLK(n4552), .C(n4553) );
  CKBD0 U4436 ( .CLK(n4553), .C(n4554) );
  CKBD0 U4437 ( .CLK(n4554), .C(n4555) );
  BUFFD0 U4438 ( .I(n4555), .Z(n4556) );
  CKBD0 U4439 ( .CLK(n4556), .C(n4557) );
  CKBD0 U4440 ( .CLK(n4557), .C(n4558) );
  CKBD0 U4441 ( .CLK(n4558), .C(n4559) );
  CKBD0 U4442 ( .CLK(n4559), .C(n4560) );
  CKBD0 U4443 ( .CLK(n4560), .C(n4561) );
  CKBD0 U4444 ( .CLK(n4561), .C(n4562) );
  CKBD0 U4445 ( .CLK(n4562), .C(n4563) );
  CKBD0 U4446 ( .CLK(n4563), .C(n4564) );
  CKBD0 U4447 ( .CLK(n4564), .C(n4565) );
  CKBD0 U4448 ( .CLK(n4565), .C(n4566) );
  BUFFD0 U4449 ( .I(n4566), .Z(n4567) );
  CKBD0 U4450 ( .CLK(n4567), .C(n4568) );
  CKBD0 U4451 ( .CLK(n4568), .C(n4569) );
  CKBD0 U4452 ( .CLK(n4569), .C(n4570) );
  CKBD0 U4453 ( .CLK(n4570), .C(n4571) );
  CKBD0 U4454 ( .CLK(n4571), .C(n4572) );
  CKBD0 U4455 ( .CLK(n4572), .C(n4573) );
  CKBD0 U4456 ( .CLK(n4573), .C(n4574) );
  CKBD0 U4457 ( .CLK(n4574), .C(n4575) );
  CKBD0 U4458 ( .CLK(n4575), .C(n4576) );
  CKBD0 U4459 ( .CLK(n4576), .C(n4577) );
  BUFFD0 U4460 ( .I(n4577), .Z(n4578) );
  CKBD0 U4461 ( .CLK(n4578), .C(n4579) );
  CKBD0 U4462 ( .CLK(n4579), .C(n4580) );
  CKBD0 U4463 ( .CLK(n4580), .C(n4581) );
  CKBD0 U4464 ( .CLK(n4581), .C(n4582) );
  CKBD0 U4465 ( .CLK(n4582), .C(n4583) );
  CKBD0 U4466 ( .CLK(n4583), .C(n4584) );
  CKBD0 U4467 ( .CLK(n4584), .C(n4585) );
  CKBD0 U4468 ( .CLK(n4585), .C(n4586) );
  CKBD0 U4469 ( .CLK(n4586), .C(n4587) );
  BUFFD0 U4470 ( .I(n4587), .Z(n4588) );
  CKBD0 U4471 ( .CLK(n4588), .C(n4589) );
  CKBD0 U4472 ( .CLK(n4589), .C(n4590) );
  CKBD0 U4473 ( .CLK(n4590), .C(n4591) );
  CKBD0 U4474 ( .CLK(n4591), .C(n4592) );
  CKBD0 U4475 ( .CLK(n4592), .C(n4593) );
  CKBD0 U4476 ( .CLK(n4593), .C(n4594) );
  CKBD0 U4477 ( .CLK(n4594), .C(n4595) );
  CKBD0 U4478 ( .CLK(n4595), .C(n4596) );
  CKBD0 U4479 ( .CLK(n4596), .C(n4597) );
  CKBD0 U4480 ( .CLK(n4597), .C(n4598) );
  CKBD0 U4481 ( .CLK(n4598), .C(n4599) );
  BUFFD0 U4482 ( .I(n4599), .Z(n4600) );
  CKBD0 U4483 ( .CLK(n4600), .C(n4601) );
  CKBD0 U4484 ( .CLK(n4601), .C(n4602) );
  CKBD0 U4485 ( .CLK(n4602), .C(n4603) );
  CKBD0 U4486 ( .CLK(n4603), .C(n4604) );
  CKBD0 U4487 ( .CLK(n4604), .C(n4605) );
  CKBD0 U4488 ( .CLK(n4605), .C(n4606) );
  CKBD0 U4489 ( .CLK(n4606), .C(n4607) );
  CKBD0 U4490 ( .CLK(n4607), .C(n4608) );
  CKBD0 U4491 ( .CLK(n4608), .C(n4609) );
  BUFFD0 U4492 ( .I(n4609), .Z(n4610) );
  CKBD0 U4493 ( .CLK(n4610), .C(n4611) );
  CKBD0 U4494 ( .CLK(n4611), .C(n4612) );
  CKBD0 U4495 ( .CLK(n4612), .C(n4613) );
  CKBD0 U4496 ( .CLK(n4613), .C(n4614) );
  CKBD0 U4497 ( .CLK(n4614), .C(n4615) );
  CKBD0 U4498 ( .CLK(n4615), .C(n4616) );
  CKBD0 U4499 ( .CLK(n4616), .C(n4617) );
  CKBD0 U4500 ( .CLK(n4617), .C(n4618) );
  CKBD0 U4501 ( .CLK(n4618), .C(n4619) );
  CKBD0 U4502 ( .CLK(n4619), .C(n4620) );
  BUFFD0 U4503 ( .I(n4620), .Z(n4621) );
  CKBD0 U4504 ( .CLK(n4621), .C(n4622) );
  CKBD0 U4505 ( .CLK(n4622), .C(n4623) );
  CKBD0 U4506 ( .CLK(n4623), .C(n4624) );
  CKBD0 U4507 ( .CLK(n4624), .C(n4625) );
  CKBD0 U4508 ( .CLK(n4625), .C(n4626) );
  CKBD0 U4509 ( .CLK(n4626), .C(n4627) );
  CKBD0 U4510 ( .CLK(n4627), .C(n4628) );
  CKBD0 U4511 ( .CLK(n4628), .C(n4629) );
  CKBD0 U4512 ( .CLK(n4629), .C(n4630) );
  CKBD0 U4513 ( .CLK(n4630), .C(n4631) );
  BUFFD0 U4514 ( .I(n4631), .Z(n4632) );
  CKBD0 U4515 ( .CLK(n4632), .C(n4633) );
  CKBD0 U4516 ( .CLK(n4633), .C(n4634) );
  CKBD0 U4517 ( .CLK(n4634), .C(n4635) );
  CKBD0 U4518 ( .CLK(n4635), .C(n4636) );
  CKBD0 U4519 ( .CLK(n4636), .C(n4637) );
  CKBD0 U4520 ( .CLK(n4637), .C(n4638) );
  CKBD0 U4521 ( .CLK(n4638), .C(n4639) );
  CKBD0 U4522 ( .CLK(n4639), .C(n4640) );
  CKBD0 U4523 ( .CLK(n4640), .C(n4641) );
  CKBD0 U4524 ( .CLK(n4641), .C(n4642) );
  BUFFD0 U4525 ( .I(n4642), .Z(n4643) );
  CKBD0 U4526 ( .CLK(n4643), .C(n4644) );
  CKBD0 U4527 ( .CLK(n4644), .C(n4645) );
  CKBD0 U4528 ( .CLK(n4645), .C(n4646) );
  CKBD0 U4529 ( .CLK(n4646), .C(n4647) );
  CKBD0 U4530 ( .CLK(n4647), .C(n4648) );
  CKBD0 U4531 ( .CLK(n4648), .C(n4649) );
  CKBD0 U4532 ( .CLK(n4649), .C(n4650) );
  CKBD0 U4533 ( .CLK(n4650), .C(n4651) );
  CKBD0 U4534 ( .CLK(n4651), .C(n4652) );
  BUFFD0 U4535 ( .I(n4652), .Z(n4653) );
  CKBD0 U4536 ( .CLK(n4653), .C(n4654) );
  CKBD0 U4537 ( .CLK(n4654), .C(n4655) );
  CKBD0 U4538 ( .CLK(n4655), .C(n4656) );
  CKBD0 U4539 ( .CLK(n4656), .C(n4657) );
  CKBD0 U4540 ( .CLK(n4657), .C(n4658) );
  CKBD0 U4541 ( .CLK(n4658), .C(n4659) );
  BUFFD0 U4542 ( .I(n4659), .Z(n4660) );
  CKBD0 U4543 ( .CLK(n4660), .C(n4661) );
  BUFFD0 U4544 ( .I(n4661), .Z(n4662) );
  CKBD0 U4545 ( .CLK(n4662), .C(n4663) );
  BUFFD0 U4546 ( .I(n4663), .Z(n4664) );
  CKBD0 U4547 ( .CLK(n4664), .C(n4665) );
  BUFFD0 U4548 ( .I(n4665), .Z(n4666) );
  CKBD0 U4549 ( .CLK(n4666), .C(n4667) );
  BUFFD0 U4550 ( .I(n4667), .Z(n4668) );
  CKBD0 U4551 ( .CLK(n4668), .C(n4669) );
  BUFFD0 U4552 ( .I(n4669), .Z(n4670) );
  CKBD0 U4553 ( .CLK(n4670), .C(n4671) );
  BUFFD0 U4554 ( .I(n4671), .Z(n4672) );
  CKBD0 U4555 ( .CLK(n4672), .C(n4673) );
  BUFFD0 U4556 ( .I(n4673), .Z(n4674) );
  BUFFD0 U4557 ( .I(n4676), .Z(n4675) );
  BUFFD0 U4558 ( .I(n4677), .Z(n4676) );
  BUFFD0 U4559 ( .I(n147), .Z(n4677) );
  CKBD0 U4560 ( .CLK(n1063), .C(n4678) );
  CKBD0 U4561 ( .CLK(n4678), .C(n4679) );
  CKBD0 U4562 ( .CLK(n4679), .C(n4680) );
  BUFFD0 U4563 ( .I(n4680), .Z(n4681) );
  CKBD0 U4564 ( .CLK(n4681), .C(n4682) );
  CKBD0 U4565 ( .CLK(n4682), .C(n4683) );
  CKBD0 U4566 ( .CLK(n4683), .C(n4684) );
  CKBD0 U4567 ( .CLK(n4684), .C(n4685) );
  CKBD0 U4568 ( .CLK(n4685), .C(n4686) );
  CKBD0 U4569 ( .CLK(n4686), .C(n4687) );
  CKBD0 U4570 ( .CLK(n4687), .C(n4688) );
  CKBD0 U4571 ( .CLK(n4688), .C(n4689) );
  CKBD0 U4572 ( .CLK(n4689), .C(n4690) );
  CKBD0 U4573 ( .CLK(n4690), .C(n4691) );
  BUFFD0 U4574 ( .I(n4691), .Z(n4692) );
  CKBD0 U4575 ( .CLK(n4692), .C(n4693) );
  CKBD0 U4576 ( .CLK(n4693), .C(n4694) );
  CKBD0 U4577 ( .CLK(n4694), .C(n4695) );
  CKBD0 U4578 ( .CLK(n4695), .C(n4696) );
  CKBD0 U4579 ( .CLK(n4696), .C(n4697) );
  CKBD0 U4580 ( .CLK(n4697), .C(n4698) );
  CKBD0 U4581 ( .CLK(n4698), .C(n4699) );
  CKBD0 U4582 ( .CLK(n4699), .C(n4700) );
  CKBD0 U4583 ( .CLK(n4700), .C(n4701) );
  CKBD0 U4584 ( .CLK(n4701), .C(n4702) );
  BUFFD0 U4585 ( .I(n4702), .Z(n4703) );
  CKBD0 U4586 ( .CLK(n4703), .C(n4704) );
  CKBD0 U4587 ( .CLK(n4704), .C(n4705) );
  CKBD0 U4588 ( .CLK(n4705), .C(n4706) );
  CKBD0 U4589 ( .CLK(n4706), .C(n4707) );
  CKBD0 U4590 ( .CLK(n4707), .C(n4708) );
  CKBD0 U4591 ( .CLK(n4708), .C(n4709) );
  CKBD0 U4592 ( .CLK(n4709), .C(n4710) );
  CKBD0 U4593 ( .CLK(n4710), .C(n4711) );
  CKBD0 U4594 ( .CLK(n4711), .C(n4712) );
  CKBD0 U4595 ( .CLK(n4712), .C(n4713) );
  BUFFD0 U4596 ( .I(n4713), .Z(n4714) );
  CKBD0 U4597 ( .CLK(n4714), .C(n4715) );
  CKBD0 U4598 ( .CLK(n4715), .C(n4716) );
  CKBD0 U4599 ( .CLK(n4716), .C(n4717) );
  CKBD0 U4600 ( .CLK(n4717), .C(n4718) );
  CKBD0 U4601 ( .CLK(n4718), .C(n4719) );
  CKBD0 U4602 ( .CLK(n4719), .C(n4720) );
  CKBD0 U4603 ( .CLK(n4720), .C(n4721) );
  CKBD0 U4604 ( .CLK(n4721), .C(n4722) );
  CKBD0 U4605 ( .CLK(n4722), .C(n4723) );
  BUFFD0 U4606 ( .I(n4723), .Z(n4724) );
  CKBD0 U4607 ( .CLK(n4724), .C(n4725) );
  CKBD0 U4608 ( .CLK(n4725), .C(n4726) );
  CKBD0 U4609 ( .CLK(n4726), .C(n4727) );
  CKBD0 U4610 ( .CLK(n4727), .C(n4728) );
  CKBD0 U4611 ( .CLK(n4728), .C(n4729) );
  CKBD0 U4612 ( .CLK(n4729), .C(n4730) );
  CKBD0 U4613 ( .CLK(n4730), .C(n4731) );
  CKBD0 U4614 ( .CLK(n4731), .C(n4732) );
  CKBD0 U4615 ( .CLK(n4732), .C(n4733) );
  CKBD0 U4616 ( .CLK(n4733), .C(n4734) );
  CKBD0 U4617 ( .CLK(n4734), .C(n4735) );
  BUFFD0 U4618 ( .I(n4735), .Z(n4736) );
  CKBD0 U4619 ( .CLK(n4736), .C(n4737) );
  CKBD0 U4620 ( .CLK(n4737), .C(n4738) );
  CKBD0 U4621 ( .CLK(n4738), .C(n4739) );
  CKBD0 U4622 ( .CLK(n4739), .C(n4740) );
  CKBD0 U4623 ( .CLK(n4740), .C(n4741) );
  CKBD0 U4624 ( .CLK(n4741), .C(n4742) );
  CKBD0 U4625 ( .CLK(n4742), .C(n4743) );
  CKBD0 U4626 ( .CLK(n4743), .C(n4744) );
  CKBD0 U4627 ( .CLK(n4744), .C(n4745) );
  BUFFD0 U4628 ( .I(n4745), .Z(n4746) );
  CKBD0 U4629 ( .CLK(n4746), .C(n4747) );
  CKBD0 U4630 ( .CLK(n4747), .C(n4748) );
  CKBD0 U4631 ( .CLK(n4748), .C(n4749) );
  CKBD0 U4632 ( .CLK(n4749), .C(n4750) );
  CKBD0 U4633 ( .CLK(n4750), .C(n4751) );
  CKBD0 U4634 ( .CLK(n4751), .C(n4752) );
  CKBD0 U4635 ( .CLK(n4752), .C(n4753) );
  CKBD0 U4636 ( .CLK(n4753), .C(n4754) );
  CKBD0 U4637 ( .CLK(n4754), .C(n4755) );
  CKBD0 U4638 ( .CLK(n4755), .C(n4756) );
  BUFFD0 U4639 ( .I(n4756), .Z(n4757) );
  CKBD0 U4640 ( .CLK(n4757), .C(n4758) );
  CKBD0 U4641 ( .CLK(n4758), .C(n4759) );
  CKBD0 U4642 ( .CLK(n4759), .C(n4760) );
  CKBD0 U4643 ( .CLK(n4760), .C(n4761) );
  CKBD0 U4644 ( .CLK(n4761), .C(n4762) );
  CKBD0 U4645 ( .CLK(n4762), .C(n4763) );
  CKBD0 U4646 ( .CLK(n4763), .C(n4764) );
  CKBD0 U4647 ( .CLK(n4764), .C(n4765) );
  CKBD0 U4648 ( .CLK(n4765), .C(n4766) );
  CKBD0 U4649 ( .CLK(n4766), .C(n4767) );
  BUFFD0 U4650 ( .I(n4767), .Z(n4768) );
  CKBD0 U4651 ( .CLK(n4768), .C(n4769) );
  CKBD0 U4652 ( .CLK(n4769), .C(n4770) );
  CKBD0 U4653 ( .CLK(n4770), .C(n4771) );
  CKBD0 U4654 ( .CLK(n4771), .C(n4772) );
  CKBD0 U4655 ( .CLK(n4772), .C(n4773) );
  CKBD0 U4656 ( .CLK(n4773), .C(n4774) );
  CKBD0 U4657 ( .CLK(n4774), .C(n4775) );
  CKBD0 U4658 ( .CLK(n4775), .C(n4776) );
  CKBD0 U4659 ( .CLK(n4776), .C(n4777) );
  CKBD0 U4660 ( .CLK(n4777), .C(n4778) );
  BUFFD0 U4661 ( .I(n4778), .Z(n4779) );
  CKBD0 U4662 ( .CLK(n4779), .C(n4780) );
  CKBD0 U4663 ( .CLK(n4780), .C(n4781) );
  CKBD0 U4664 ( .CLK(n4781), .C(n4782) );
  CKBD0 U4665 ( .CLK(n4782), .C(n4783) );
  CKBD0 U4666 ( .CLK(n4783), .C(n4784) );
  CKBD0 U4667 ( .CLK(n4784), .C(n4785) );
  CKBD0 U4668 ( .CLK(n4785), .C(n4786) );
  CKBD0 U4669 ( .CLK(n4786), .C(n4787) );
  CKBD0 U4670 ( .CLK(n4787), .C(n4788) );
  CKBD0 U4671 ( .CLK(n4788), .C(n4789) );
  BUFFD0 U4672 ( .I(n4789), .Z(n4790) );
  CKBD0 U4673 ( .CLK(n4790), .C(n4791) );
  CKBD0 U4674 ( .CLK(n4791), .C(n4792) );
  CKBD0 U4675 ( .CLK(n4792), .C(n4793) );
  CKBD0 U4676 ( .CLK(n4793), .C(n4794) );
  CKBD0 U4677 ( .CLK(n4794), .C(n4795) );
  BUFFD0 U4678 ( .I(n4795), .Z(n4796) );
  CKBD0 U4679 ( .CLK(n4796), .C(n4797) );
  BUFFD0 U4680 ( .I(n4797), .Z(n4798) );
  CKBD0 U4681 ( .CLK(n4798), .C(n4799) );
  BUFFD0 U4682 ( .I(n4799), .Z(n4800) );
  CKBD0 U4683 ( .CLK(n4800), .C(n4801) );
  BUFFD0 U4684 ( .I(n4801), .Z(n4802) );
  CKBD0 U4685 ( .CLK(n4802), .C(n4803) );
  BUFFD0 U4686 ( .I(n4803), .Z(n4804) );
  CKBD0 U4687 ( .CLK(n4804), .C(n4805) );
  BUFFD0 U4688 ( .I(n4805), .Z(n4806) );
  CKBD0 U4689 ( .CLK(n4806), .C(n4807) );
  BUFFD0 U4690 ( .I(n4807), .Z(n4808) );
  CKBD0 U4691 ( .CLK(n4808), .C(n4809) );
  BUFFD0 U4692 ( .I(n4809), .Z(n4810) );
  BUFFD0 U4693 ( .I(n4812), .Z(n4811) );
  BUFFD0 U4694 ( .I(n4813), .Z(n4812) );
  BUFFD0 U4695 ( .I(n146), .Z(n4813) );
  CKBD0 U4696 ( .CLK(n1061), .C(n4814) );
  CKBD0 U4697 ( .CLK(n4814), .C(n4815) );
  CKBD0 U4698 ( .CLK(n4815), .C(n4816) );
  BUFFD0 U4699 ( .I(n4816), .Z(n4817) );
  CKBD0 U4700 ( .CLK(n4817), .C(n4818) );
  CKBD0 U4701 ( .CLK(n4818), .C(n4819) );
  CKBD0 U4702 ( .CLK(n4819), .C(n4820) );
  CKBD0 U4703 ( .CLK(n4820), .C(n4821) );
  CKBD0 U4704 ( .CLK(n4821), .C(n4822) );
  CKBD0 U4705 ( .CLK(n4822), .C(n4823) );
  CKBD0 U4706 ( .CLK(n4823), .C(n4824) );
  CKBD0 U4707 ( .CLK(n4824), .C(n4825) );
  CKBD0 U4708 ( .CLK(n4825), .C(n4826) );
  CKBD0 U4709 ( .CLK(n4826), .C(n4827) );
  BUFFD0 U4710 ( .I(n4827), .Z(n4828) );
  CKBD0 U4711 ( .CLK(n4828), .C(n4829) );
  CKBD0 U4712 ( .CLK(n4829), .C(n4830) );
  CKBD0 U4713 ( .CLK(n4830), .C(n4831) );
  CKBD0 U4714 ( .CLK(n4831), .C(n4832) );
  CKBD0 U4715 ( .CLK(n4832), .C(n4833) );
  CKBD0 U4716 ( .CLK(n4833), .C(n4834) );
  CKBD0 U4717 ( .CLK(n4834), .C(n4835) );
  CKBD0 U4718 ( .CLK(n4835), .C(n4836) );
  CKBD0 U4719 ( .CLK(n4836), .C(n4837) );
  CKBD0 U4720 ( .CLK(n4837), .C(n4838) );
  BUFFD0 U4721 ( .I(n4838), .Z(n4839) );
  CKBD0 U4722 ( .CLK(n4839), .C(n4840) );
  CKBD0 U4723 ( .CLK(n4840), .C(n4841) );
  CKBD0 U4724 ( .CLK(n4841), .C(n4842) );
  CKBD0 U4725 ( .CLK(n4842), .C(n4843) );
  CKBD0 U4726 ( .CLK(n4843), .C(n4844) );
  CKBD0 U4727 ( .CLK(n4844), .C(n4845) );
  CKBD0 U4728 ( .CLK(n4845), .C(n4846) );
  CKBD0 U4729 ( .CLK(n4846), .C(n4847) );
  CKBD0 U4730 ( .CLK(n4847), .C(n4848) );
  CKBD0 U4731 ( .CLK(n4848), .C(n4849) );
  BUFFD0 U4732 ( .I(n4849), .Z(n4850) );
  CKBD0 U4733 ( .CLK(n4850), .C(n4851) );
  CKBD0 U4734 ( .CLK(n4851), .C(n4852) );
  CKBD0 U4735 ( .CLK(n4852), .C(n4853) );
  CKBD0 U4736 ( .CLK(n4853), .C(n4854) );
  CKBD0 U4737 ( .CLK(n4854), .C(n4855) );
  CKBD0 U4738 ( .CLK(n4855), .C(n4856) );
  CKBD0 U4739 ( .CLK(n4856), .C(n4857) );
  CKBD0 U4740 ( .CLK(n4857), .C(n4858) );
  CKBD0 U4741 ( .CLK(n4858), .C(n4859) );
  CKBD0 U4742 ( .CLK(n4859), .C(n4860) );
  BUFFD0 U4743 ( .I(n4860), .Z(n4861) );
  CKBD0 U4744 ( .CLK(n4861), .C(n4862) );
  CKBD0 U4745 ( .CLK(n4862), .C(n4863) );
  CKBD0 U4746 ( .CLK(n4863), .C(n4864) );
  CKBD0 U4747 ( .CLK(n4864), .C(n4865) );
  CKBD0 U4748 ( .CLK(n4865), .C(n4866) );
  CKBD0 U4749 ( .CLK(n4866), .C(n4867) );
  CKBD0 U4750 ( .CLK(n4867), .C(n4868) );
  CKBD0 U4751 ( .CLK(n4868), .C(n4869) );
  CKBD0 U4752 ( .CLK(n4869), .C(n4870) );
  CKBD0 U4753 ( .CLK(n4870), .C(n4871) );
  BUFFD0 U4754 ( .I(n4871), .Z(n4872) );
  CKBD0 U4755 ( .CLK(n4872), .C(n4873) );
  CKBD0 U4756 ( .CLK(n4873), .C(n4874) );
  CKBD0 U4757 ( .CLK(n4874), .C(n4875) );
  CKBD0 U4758 ( .CLK(n4875), .C(n4876) );
  CKBD0 U4759 ( .CLK(n4876), .C(n4877) );
  CKBD0 U4760 ( .CLK(n4877), .C(n4878) );
  CKBD0 U4761 ( .CLK(n4878), .C(n4879) );
  CKBD0 U4762 ( .CLK(n4879), .C(n4880) );
  CKBD0 U4763 ( .CLK(n4880), .C(n4881) );
  BUFFD0 U4764 ( .I(n4881), .Z(n4882) );
  CKBD0 U4765 ( .CLK(n4882), .C(n4883) );
  CKBD0 U4766 ( .CLK(n4883), .C(n4884) );
  CKBD0 U4767 ( .CLK(n4884), .C(n4885) );
  CKBD0 U4768 ( .CLK(n4885), .C(n4886) );
  CKBD0 U4769 ( .CLK(n4886), .C(n4887) );
  CKBD0 U4770 ( .CLK(n4887), .C(n4888) );
  CKBD0 U4771 ( .CLK(n4888), .C(n4889) );
  CKBD0 U4772 ( .CLK(n4889), .C(n4890) );
  CKBD0 U4773 ( .CLK(n4890), .C(n4891) );
  CKBD0 U4774 ( .CLK(n4891), .C(n4892) );
  CKBD0 U4775 ( .CLK(n4892), .C(n4893) );
  BUFFD0 U4776 ( .I(n4893), .Z(n4894) );
  CKBD0 U4777 ( .CLK(n4894), .C(n4895) );
  CKBD0 U4778 ( .CLK(n4895), .C(n4896) );
  CKBD0 U4779 ( .CLK(n4896), .C(n4897) );
  CKBD0 U4780 ( .CLK(n4897), .C(n4898) );
  CKBD0 U4781 ( .CLK(n4898), .C(n4899) );
  CKBD0 U4782 ( .CLK(n4899), .C(n4900) );
  CKBD0 U4783 ( .CLK(n4900), .C(n4901) );
  CKBD0 U4784 ( .CLK(n4901), .C(n4902) );
  CKBD0 U4785 ( .CLK(n4902), .C(n4903) );
  BUFFD0 U4786 ( .I(n4903), .Z(n4904) );
  CKBD0 U4787 ( .CLK(n4904), .C(n4905) );
  CKBD0 U4788 ( .CLK(n4905), .C(n4906) );
  CKBD0 U4789 ( .CLK(n4906), .C(n4907) );
  CKBD0 U4790 ( .CLK(n4907), .C(n4908) );
  CKBD0 U4791 ( .CLK(n4908), .C(n4909) );
  CKBD0 U4792 ( .CLK(n4909), .C(n4910) );
  CKBD0 U4793 ( .CLK(n4910), .C(n4911) );
  CKBD0 U4794 ( .CLK(n4911), .C(n4912) );
  CKBD0 U4795 ( .CLK(n4912), .C(n4913) );
  BUFFD0 U4796 ( .I(n4913), .Z(n4914) );
  CKBD0 U4797 ( .CLK(n4914), .C(n4915) );
  CKBD0 U4798 ( .CLK(n4915), .C(n4916) );
  CKBD0 U4799 ( .CLK(n4916), .C(n4917) );
  CKBD0 U4800 ( .CLK(n4917), .C(n4918) );
  CKBD0 U4801 ( .CLK(n4918), .C(n4919) );
  CKBD0 U4802 ( .CLK(n4919), .C(n4920) );
  CKBD0 U4803 ( .CLK(n4920), .C(n4921) );
  CKBD0 U4804 ( .CLK(n4921), .C(n4922) );
  CKBD0 U4805 ( .CLK(n4922), .C(n4923) );
  CKBD0 U4806 ( .CLK(n4923), .C(n4924) );
  CKBD0 U4807 ( .CLK(n4924), .C(n4925) );
  BUFFD0 U4808 ( .I(n4925), .Z(n4926) );
  CKBD0 U4809 ( .CLK(n4926), .C(n4927) );
  CKBD0 U4810 ( .CLK(n4927), .C(n4928) );
  CKBD0 U4811 ( .CLK(n4928), .C(n4929) );
  CKBD0 U4812 ( .CLK(n4929), .C(n4930) );
  CKBD0 U4813 ( .CLK(n4930), .C(n4931) );
  BUFFD0 U4814 ( .I(n4931), .Z(n4932) );
  CKBD0 U4815 ( .CLK(n4932), .C(n4933) );
  BUFFD0 U4816 ( .I(n4933), .Z(n4934) );
  CKBD0 U4817 ( .CLK(n4934), .C(n4935) );
  BUFFD0 U4818 ( .I(n4935), .Z(n4936) );
  CKBD0 U4819 ( .CLK(n4936), .C(n4937) );
  BUFFD0 U4820 ( .I(n4937), .Z(n4938) );
  CKBD0 U4821 ( .CLK(n4938), .C(n4939) );
  BUFFD0 U4822 ( .I(n4939), .Z(n4940) );
  CKBD0 U4823 ( .CLK(n4940), .C(n4941) );
  BUFFD0 U4824 ( .I(n4941), .Z(n4942) );
  CKBD0 U4825 ( .CLK(n4942), .C(n4943) );
  BUFFD0 U4826 ( .I(n4943), .Z(n4944) );
  CKBD0 U4827 ( .CLK(n4944), .C(n4945) );
  BUFFD0 U4828 ( .I(n4945), .Z(n4946) );
  BUFFD0 U4829 ( .I(n4948), .Z(n4947) );
  BUFFD0 U4830 ( .I(n4949), .Z(n4948) );
  BUFFD0 U4831 ( .I(n145), .Z(n4949) );
  CKBD0 U4832 ( .CLK(n1059), .C(n4950) );
  CKBD0 U4833 ( .CLK(n4950), .C(n4951) );
  CKBD0 U4834 ( .CLK(n4951), .C(n4952) );
  BUFFD0 U4835 ( .I(n4952), .Z(n4953) );
  CKBD0 U4836 ( .CLK(n4953), .C(n4954) );
  CKBD0 U4837 ( .CLK(n4954), .C(n4955) );
  CKBD0 U4838 ( .CLK(n4955), .C(n4956) );
  CKBD0 U4839 ( .CLK(n4956), .C(n4957) );
  CKBD0 U4840 ( .CLK(n4957), .C(n4958) );
  CKBD0 U4841 ( .CLK(n4958), .C(n4959) );
  CKBD0 U4842 ( .CLK(n4959), .C(n4960) );
  CKBD0 U4843 ( .CLK(n4960), .C(n4961) );
  CKBD0 U4844 ( .CLK(n4961), .C(n4962) );
  CKBD0 U4845 ( .CLK(n4962), .C(n4963) );
  CKBD0 U4846 ( .CLK(n4963), .C(n4964) );
  BUFFD0 U4847 ( .I(n4964), .Z(n4965) );
  CKBD0 U4848 ( .CLK(n4965), .C(n4966) );
  CKBD0 U4849 ( .CLK(n4966), .C(n4967) );
  CKBD0 U4850 ( .CLK(n4967), .C(n4968) );
  CKBD0 U4851 ( .CLK(n4968), .C(n4969) );
  CKBD0 U4852 ( .CLK(n4969), .C(n4970) );
  CKBD0 U4853 ( .CLK(n4970), .C(n4971) );
  CKBD0 U4854 ( .CLK(n4971), .C(n4972) );
  CKBD0 U4855 ( .CLK(n4972), .C(n4973) );
  CKBD0 U4856 ( .CLK(n4973), .C(n4974) );
  BUFFD0 U4857 ( .I(n4974), .Z(n4975) );
  CKBD0 U4858 ( .CLK(n4975), .C(n4976) );
  CKBD0 U4859 ( .CLK(n4976), .C(n4977) );
  CKBD0 U4860 ( .CLK(n4977), .C(n4978) );
  CKBD0 U4861 ( .CLK(n4978), .C(n4979) );
  CKBD0 U4862 ( .CLK(n4979), .C(n4980) );
  CKBD0 U4863 ( .CLK(n4980), .C(n4981) );
  CKBD0 U4864 ( .CLK(n4981), .C(n4982) );
  CKBD0 U4865 ( .CLK(n4982), .C(n4983) );
  CKBD0 U4866 ( .CLK(n4983), .C(n4984) );
  BUFFD0 U4867 ( .I(n4984), .Z(n4985) );
  CKBD0 U4868 ( .CLK(n4985), .C(n4986) );
  CKBD0 U4869 ( .CLK(n4986), .C(n4987) );
  CKBD0 U4870 ( .CLK(n4987), .C(n4988) );
  CKBD0 U4871 ( .CLK(n4988), .C(n4989) );
  CKBD0 U4872 ( .CLK(n4989), .C(n4990) );
  CKBD0 U4873 ( .CLK(n4990), .C(n4991) );
  CKBD0 U4874 ( .CLK(n4991), .C(n4992) );
  CKBD0 U4875 ( .CLK(n4992), .C(n4993) );
  CKBD0 U4876 ( .CLK(n4993), .C(n4994) );
  CKBD0 U4877 ( .CLK(n4994), .C(n4995) );
  CKBD0 U4878 ( .CLK(n4995), .C(n4996) );
  BUFFD0 U4879 ( .I(n4996), .Z(n4997) );
  CKBD0 U4880 ( .CLK(n4997), .C(n4998) );
  CKBD0 U4881 ( .CLK(n4998), .C(n4999) );
  CKBD0 U4882 ( .CLK(n4999), .C(n5000) );
  CKBD0 U4883 ( .CLK(n5000), .C(n5001) );
  CKBD0 U4884 ( .CLK(n5001), .C(n5002) );
  CKBD0 U4885 ( .CLK(n5002), .C(n5003) );
  CKBD0 U4886 ( .CLK(n5003), .C(n5004) );
  CKBD0 U4887 ( .CLK(n5004), .C(n5005) );
  CKBD0 U4888 ( .CLK(n5005), .C(n5006) );
  BUFFD0 U4889 ( .I(n5006), .Z(n5007) );
  CKBD0 U4890 ( .CLK(n5007), .C(n5008) );
  CKBD0 U4891 ( .CLK(n5008), .C(n5009) );
  CKBD0 U4892 ( .CLK(n5009), .C(n5010) );
  CKBD0 U4893 ( .CLK(n5010), .C(n5011) );
  CKBD0 U4894 ( .CLK(n5011), .C(n5012) );
  CKBD0 U4895 ( .CLK(n5012), .C(n5013) );
  CKBD0 U4896 ( .CLK(n5013), .C(n5014) );
  CKBD0 U4897 ( .CLK(n5014), .C(n5015) );
  CKBD0 U4898 ( .CLK(n5015), .C(n5016) );
  CKBD0 U4899 ( .CLK(n5016), .C(n5017) );
  BUFFD0 U4900 ( .I(n5017), .Z(n5018) );
  CKBD0 U4901 ( .CLK(n5018), .C(n5019) );
  CKBD0 U4902 ( .CLK(n5019), .C(n5020) );
  CKBD0 U4903 ( .CLK(n5020), .C(n5021) );
  CKBD0 U4904 ( .CLK(n5021), .C(n5022) );
  CKBD0 U4905 ( .CLK(n5022), .C(n5023) );
  CKBD0 U4906 ( .CLK(n5023), .C(n5024) );
  CKBD0 U4907 ( .CLK(n5024), .C(n5025) );
  CKBD0 U4908 ( .CLK(n5025), .C(n5026) );
  CKBD0 U4909 ( .CLK(n5026), .C(n5027) );
  CKBD0 U4910 ( .CLK(n5027), .C(n5028) );
  BUFFD0 U4911 ( .I(n5028), .Z(n5029) );
  CKBD0 U4912 ( .CLK(n5029), .C(n5030) );
  CKBD0 U4913 ( .CLK(n5030), .C(n5031) );
  CKBD0 U4914 ( .CLK(n5031), .C(n5032) );
  CKBD0 U4915 ( .CLK(n5032), .C(n5033) );
  CKBD0 U4916 ( .CLK(n5033), .C(n5034) );
  CKBD0 U4917 ( .CLK(n5034), .C(n5035) );
  CKBD0 U4918 ( .CLK(n5035), .C(n5036) );
  CKBD0 U4919 ( .CLK(n5036), .C(n5037) );
  CKBD0 U4920 ( .CLK(n5037), .C(n5038) );
  CKBD0 U4921 ( .CLK(n5038), .C(n5039) );
  BUFFD0 U4922 ( .I(n5039), .Z(n5040) );
  CKBD0 U4923 ( .CLK(n5040), .C(n5041) );
  CKBD0 U4924 ( .CLK(n5041), .C(n5042) );
  CKBD0 U4925 ( .CLK(n5042), .C(n5043) );
  CKBD0 U4926 ( .CLK(n5043), .C(n5044) );
  CKBD0 U4927 ( .CLK(n5044), .C(n5045) );
  CKBD0 U4928 ( .CLK(n5045), .C(n5046) );
  CKBD0 U4929 ( .CLK(n5046), .C(n5047) );
  CKBD0 U4930 ( .CLK(n5047), .C(n5048) );
  CKBD0 U4931 ( .CLK(n5048), .C(n5049) );
  BUFFD0 U4932 ( .I(n5049), .Z(n5050) );
  CKBD0 U4933 ( .CLK(n5050), .C(n5051) );
  CKBD0 U4934 ( .CLK(n5051), .C(n5052) );
  CKBD0 U4935 ( .CLK(n5052), .C(n5053) );
  CKBD0 U4936 ( .CLK(n5053), .C(n5054) );
  CKBD0 U4937 ( .CLK(n5054), .C(n5055) );
  CKBD0 U4938 ( .CLK(n5055), .C(n5056) );
  CKBD0 U4939 ( .CLK(n5056), .C(n5057) );
  CKBD0 U4940 ( .CLK(n5057), .C(n5058) );
  CKBD0 U4941 ( .CLK(n5058), .C(n5059) );
  CKBD0 U4942 ( .CLK(n5059), .C(n5060) );
  CKBD0 U4943 ( .CLK(n5060), .C(n5061) );
  BUFFD0 U4944 ( .I(n5061), .Z(n5062) );
  CKBD0 U4945 ( .CLK(n5062), .C(n5063) );
  CKBD0 U4946 ( .CLK(n5063), .C(n5064) );
  CKBD0 U4947 ( .CLK(n5064), .C(n5065) );
  CKBD0 U4948 ( .CLK(n5065), .C(n5066) );
  CKBD0 U4949 ( .CLK(n5066), .C(n5067) );
  BUFFD0 U4950 ( .I(n5067), .Z(n5068) );
  CKBD0 U4951 ( .CLK(n5068), .C(n5069) );
  BUFFD0 U4952 ( .I(n5069), .Z(n5070) );
  CKBD0 U4953 ( .CLK(n5070), .C(n5071) );
  BUFFD0 U4954 ( .I(n5071), .Z(n5072) );
  CKBD0 U4955 ( .CLK(n5072), .C(n5073) );
  BUFFD0 U4956 ( .I(n5073), .Z(n5074) );
  CKBD0 U4957 ( .CLK(n5074), .C(n5075) );
  BUFFD0 U4958 ( .I(n5075), .Z(n5076) );
  CKBD0 U4959 ( .CLK(n5076), .C(n5077) );
  BUFFD0 U4960 ( .I(n5077), .Z(n5078) );
  CKBD0 U4961 ( .CLK(n5078), .C(n5079) );
  BUFFD0 U4962 ( .I(n5079), .Z(n5080) );
  CKBD0 U4963 ( .CLK(n5080), .C(n5081) );
  BUFFD0 U4964 ( .I(n5081), .Z(n5082) );
  BUFFD0 U4965 ( .I(n5084), .Z(n5083) );
  BUFFD0 U4966 ( .I(n5085), .Z(n5084) );
  BUFFD0 U4967 ( .I(n144), .Z(n5085) );
  CKBD0 U4968 ( .CLK(n1057), .C(n5086) );
  CKBD0 U4969 ( .CLK(n5086), .C(n5087) );
  CKBD0 U4970 ( .CLK(n5087), .C(n5088) );
  BUFFD0 U4971 ( .I(n5088), .Z(n5089) );
  CKBD0 U4972 ( .CLK(n5089), .C(n5090) );
  CKBD0 U4973 ( .CLK(n5090), .C(n5091) );
  CKBD0 U4974 ( .CLK(n5091), .C(n5092) );
  CKBD0 U4975 ( .CLK(n5092), .C(n5093) );
  CKBD0 U4976 ( .CLK(n5093), .C(n5094) );
  CKBD0 U4977 ( .CLK(n5094), .C(n5095) );
  CKBD0 U4978 ( .CLK(n5095), .C(n5096) );
  CKBD0 U4979 ( .CLK(n5096), .C(n5097) );
  CKBD0 U4980 ( .CLK(n5097), .C(n5098) );
  CKBD0 U4981 ( .CLK(n5098), .C(n5099) );
  BUFFD0 U4982 ( .I(n5099), .Z(n5100) );
  CKBD0 U4983 ( .CLK(n5100), .C(n5101) );
  CKBD0 U4984 ( .CLK(n5101), .C(n5102) );
  CKBD0 U4985 ( .CLK(n5102), .C(n5103) );
  CKBD0 U4986 ( .CLK(n5103), .C(n5104) );
  CKBD0 U4987 ( .CLK(n5104), .C(n5105) );
  CKBD0 U4988 ( .CLK(n5105), .C(n5106) );
  CKBD0 U4989 ( .CLK(n5106), .C(n5107) );
  CKBD0 U4990 ( .CLK(n5107), .C(n5108) );
  CKBD0 U4991 ( .CLK(n5108), .C(n5109) );
  CKBD0 U4992 ( .CLK(n5109), .C(n5110) );
  BUFFD0 U4993 ( .I(n5110), .Z(n5111) );
  CKBD0 U4994 ( .CLK(n5111), .C(n5112) );
  CKBD0 U4995 ( .CLK(n5112), .C(n5113) );
  CKBD0 U4996 ( .CLK(n5113), .C(n5114) );
  CKBD0 U4997 ( .CLK(n5114), .C(n5115) );
  CKBD0 U4998 ( .CLK(n5115), .C(n5116) );
  CKBD0 U4999 ( .CLK(n5116), .C(n5117) );
  CKBD0 U5000 ( .CLK(n5117), .C(n5118) );
  CKBD0 U5001 ( .CLK(n5118), .C(n5119) );
  CKBD0 U5002 ( .CLK(n5119), .C(n5120) );
  BUFFD0 U5003 ( .I(n5120), .Z(n5121) );
  CKBD0 U5004 ( .CLK(n5121), .C(n5122) );
  CKBD0 U5005 ( .CLK(n5122), .C(n5123) );
  CKBD0 U5006 ( .CLK(n5123), .C(n5124) );
  CKBD0 U5007 ( .CLK(n5124), .C(n5125) );
  CKBD0 U5008 ( .CLK(n5125), .C(n5126) );
  CKBD0 U5009 ( .CLK(n5126), .C(n5127) );
  CKBD0 U5010 ( .CLK(n5127), .C(n5128) );
  CKBD0 U5011 ( .CLK(n5128), .C(n5129) );
  CKBD0 U5012 ( .CLK(n5129), .C(n5130) );
  CKBD0 U5013 ( .CLK(n5130), .C(n5131) );
  CKBD0 U5014 ( .CLK(n5131), .C(n5132) );
  BUFFD0 U5015 ( .I(n5132), .Z(n5133) );
  CKBD0 U5016 ( .CLK(n5133), .C(n5134) );
  CKBD0 U5017 ( .CLK(n5134), .C(n5135) );
  CKBD0 U5018 ( .CLK(n5135), .C(n5136) );
  CKBD0 U5019 ( .CLK(n5136), .C(n5137) );
  CKBD0 U5020 ( .CLK(n5137), .C(n5138) );
  CKBD0 U5021 ( .CLK(n5138), .C(n5139) );
  CKBD0 U5022 ( .CLK(n5139), .C(n5140) );
  CKBD0 U5023 ( .CLK(n5140), .C(n5141) );
  CKBD0 U5024 ( .CLK(n5141), .C(n5142) );
  BUFFD0 U5025 ( .I(n5142), .Z(n5143) );
  CKBD0 U5026 ( .CLK(n5143), .C(n5144) );
  CKBD0 U5027 ( .CLK(n5144), .C(n5145) );
  CKBD0 U5028 ( .CLK(n5145), .C(n5146) );
  CKBD0 U5029 ( .CLK(n5146), .C(n5147) );
  CKBD0 U5030 ( .CLK(n5147), .C(n5148) );
  CKBD0 U5031 ( .CLK(n5148), .C(n5149) );
  CKBD0 U5032 ( .CLK(n5149), .C(n5150) );
  CKBD0 U5033 ( .CLK(n5150), .C(n5151) );
  CKBD0 U5034 ( .CLK(n5151), .C(n5152) );
  CKBD0 U5035 ( .CLK(n5152), .C(n5153) );
  CKBD0 U5036 ( .CLK(n5153), .C(n5154) );
  BUFFD0 U5037 ( .I(n5154), .Z(n5155) );
  CKBD0 U5038 ( .CLK(n5155), .C(n5156) );
  CKBD0 U5039 ( .CLK(n5156), .C(n5157) );
  CKBD0 U5040 ( .CLK(n5157), .C(n5158) );
  CKBD0 U5041 ( .CLK(n5158), .C(n5159) );
  CKBD0 U5042 ( .CLK(n5159), .C(n5160) );
  CKBD0 U5043 ( .CLK(n5160), .C(n5161) );
  CKBD0 U5044 ( .CLK(n5161), .C(n5162) );
  CKBD0 U5045 ( .CLK(n5162), .C(n5163) );
  CKBD0 U5046 ( .CLK(n5163), .C(n5164) );
  BUFFD0 U5047 ( .I(n5164), .Z(n5165) );
  CKBD0 U5048 ( .CLK(n5165), .C(n5166) );
  CKBD0 U5049 ( .CLK(n5166), .C(n5167) );
  CKBD0 U5050 ( .CLK(n5167), .C(n5168) );
  CKBD0 U5051 ( .CLK(n5168), .C(n5169) );
  CKBD0 U5052 ( .CLK(n5169), .C(n5170) );
  CKBD0 U5053 ( .CLK(n5170), .C(n5171) );
  CKBD0 U5054 ( .CLK(n5171), .C(n5172) );
  CKBD0 U5055 ( .CLK(n5172), .C(n5173) );
  CKBD0 U5056 ( .CLK(n5173), .C(n5174) );
  CKBD0 U5057 ( .CLK(n5174), .C(n5175) );
  BUFFD0 U5058 ( .I(n5175), .Z(n5176) );
  CKBD0 U5059 ( .CLK(n5176), .C(n5177) );
  CKBD0 U5060 ( .CLK(n5177), .C(n5178) );
  CKBD0 U5061 ( .CLK(n5178), .C(n5179) );
  CKBD0 U5062 ( .CLK(n5179), .C(n5180) );
  CKBD0 U5063 ( .CLK(n5180), .C(n5181) );
  CKBD0 U5064 ( .CLK(n5181), .C(n5182) );
  CKBD0 U5065 ( .CLK(n5182), .C(n5183) );
  CKBD0 U5066 ( .CLK(n5183), .C(n5184) );
  CKBD0 U5067 ( .CLK(n5184), .C(n5185) );
  CKBD0 U5068 ( .CLK(n5185), .C(n5186) );
  BUFFD0 U5069 ( .I(n5186), .Z(n5187) );
  CKBD0 U5070 ( .CLK(n5187), .C(n5188) );
  CKBD0 U5071 ( .CLK(n5188), .C(n5189) );
  CKBD0 U5072 ( .CLK(n5189), .C(n5190) );
  CKBD0 U5073 ( .CLK(n5190), .C(n5191) );
  CKBD0 U5074 ( .CLK(n5191), .C(n5192) );
  CKBD0 U5075 ( .CLK(n5192), .C(n5193) );
  CKBD0 U5076 ( .CLK(n5193), .C(n5194) );
  CKBD0 U5077 ( .CLK(n5194), .C(n5195) );
  CKBD0 U5078 ( .CLK(n5195), .C(n5196) );
  CKBD0 U5079 ( .CLK(n5196), .C(n5197) );
  BUFFD0 U5080 ( .I(n5197), .Z(n5198) );
  CKBD0 U5081 ( .CLK(n5198), .C(n5199) );
  CKBD0 U5082 ( .CLK(n5199), .C(n5200) );
  CKBD0 U5083 ( .CLK(n5200), .C(n5201) );
  CKBD0 U5084 ( .CLK(n5201), .C(n5202) );
  CKBD0 U5085 ( .CLK(n5202), .C(n5203) );
  BUFFD0 U5086 ( .I(n5203), .Z(n5204) );
  CKBD0 U5087 ( .CLK(n5204), .C(n5205) );
  BUFFD0 U5088 ( .I(n5205), .Z(n5206) );
  CKBD0 U5089 ( .CLK(n5206), .C(n5207) );
  BUFFD0 U5090 ( .I(n5207), .Z(n5208) );
  CKBD0 U5091 ( .CLK(n5208), .C(n5209) );
  BUFFD0 U5092 ( .I(n5209), .Z(n5210) );
  CKBD0 U5093 ( .CLK(n5210), .C(n5211) );
  BUFFD0 U5094 ( .I(n5211), .Z(n5212) );
  CKBD0 U5095 ( .CLK(n5212), .C(n5213) );
  BUFFD0 U5096 ( .I(n5213), .Z(n5214) );
  CKBD0 U5097 ( .CLK(n5214), .C(n5215) );
  BUFFD0 U5098 ( .I(n5215), .Z(n5216) );
  CKBD0 U5099 ( .CLK(n5216), .C(n5217) );
  BUFFD0 U5100 ( .I(n5217), .Z(n5218) );
  BUFFD0 U5101 ( .I(n5220), .Z(n5219) );
  BUFFD0 U5102 ( .I(n5221), .Z(n5220) );
  BUFFD0 U5103 ( .I(n143), .Z(n5221) );
  CKBD0 U5104 ( .CLK(n1055), .C(n5222) );
  CKBD0 U5105 ( .CLK(n5222), .C(n5223) );
  CKBD0 U5106 ( .CLK(n5223), .C(n5224) );
  CKBD0 U5107 ( .CLK(n5224), .C(n5225) );
  BUFFD0 U5108 ( .I(n5225), .Z(n5226) );
  CKBD0 U5109 ( .CLK(n5226), .C(n5227) );
  CKBD0 U5110 ( .CLK(n5227), .C(n5228) );
  CKBD0 U5111 ( .CLK(n5228), .C(n5229) );
  CKBD0 U5112 ( .CLK(n5229), .C(n5230) );
  CKBD0 U5113 ( .CLK(n5230), .C(n5231) );
  CKBD0 U5114 ( .CLK(n5231), .C(n5232) );
  CKBD0 U5115 ( .CLK(n5232), .C(n5233) );
  CKBD0 U5116 ( .CLK(n5233), .C(n5234) );
  CKBD0 U5117 ( .CLK(n5234), .C(n5235) );
  BUFFD0 U5118 ( .I(n5235), .Z(n5236) );
  CKBD0 U5119 ( .CLK(n5236), .C(n5237) );
  CKBD0 U5120 ( .CLK(n5237), .C(n5238) );
  CKBD0 U5121 ( .CLK(n5238), .C(n5239) );
  CKBD0 U5122 ( .CLK(n5239), .C(n5240) );
  CKBD0 U5123 ( .CLK(n5240), .C(n5241) );
  CKBD0 U5124 ( .CLK(n5241), .C(n5242) );
  CKBD0 U5125 ( .CLK(n5242), .C(n5243) );
  CKBD0 U5126 ( .CLK(n5243), .C(n5244) );
  CKBD0 U5127 ( .CLK(n5244), .C(n5245) );
  CKBD0 U5128 ( .CLK(n5245), .C(n5246) );
  BUFFD0 U5129 ( .I(n5246), .Z(n5247) );
  CKBD0 U5130 ( .CLK(n5247), .C(n5248) );
  CKBD0 U5131 ( .CLK(n5248), .C(n5249) );
  CKBD0 U5132 ( .CLK(n5249), .C(n5250) );
  CKBD0 U5133 ( .CLK(n5250), .C(n5251) );
  CKBD0 U5134 ( .CLK(n5251), .C(n5252) );
  CKBD0 U5135 ( .CLK(n5252), .C(n5253) );
  CKBD0 U5136 ( .CLK(n5253), .C(n5254) );
  CKBD0 U5137 ( .CLK(n5254), .C(n5255) );
  CKBD0 U5138 ( .CLK(n5255), .C(n5256) );
  CKBD0 U5139 ( .CLK(n5256), .C(n5257) );
  BUFFD0 U5140 ( .I(n5257), .Z(n5258) );
  CKBD0 U5141 ( .CLK(n5258), .C(n5259) );
  CKBD0 U5142 ( .CLK(n5259), .C(n5260) );
  CKBD0 U5143 ( .CLK(n5260), .C(n5261) );
  CKBD0 U5144 ( .CLK(n5261), .C(n5262) );
  CKBD0 U5145 ( .CLK(n5262), .C(n5263) );
  CKBD0 U5146 ( .CLK(n5263), .C(n5264) );
  CKBD0 U5147 ( .CLK(n5264), .C(n5265) );
  CKBD0 U5148 ( .CLK(n5265), .C(n5266) );
  CKBD0 U5149 ( .CLK(n5266), .C(n5267) );
  CKBD0 U5150 ( .CLK(n5267), .C(n5268) );
  BUFFD0 U5151 ( .I(n5268), .Z(n5269) );
  CKBD0 U5152 ( .CLK(n5269), .C(n5270) );
  CKBD0 U5153 ( .CLK(n5270), .C(n5271) );
  CKBD0 U5154 ( .CLK(n5271), .C(n5272) );
  CKBD0 U5155 ( .CLK(n5272), .C(n5273) );
  CKBD0 U5156 ( .CLK(n5273), .C(n5274) );
  CKBD0 U5157 ( .CLK(n5274), .C(n5275) );
  CKBD0 U5158 ( .CLK(n5275), .C(n5276) );
  CKBD0 U5159 ( .CLK(n5276), .C(n5277) );
  CKBD0 U5160 ( .CLK(n5277), .C(n5278) );
  BUFFD0 U5161 ( .I(n5278), .Z(n5279) );
  CKBD0 U5162 ( .CLK(n5279), .C(n5280) );
  CKBD0 U5163 ( .CLK(n5280), .C(n5281) );
  CKBD0 U5164 ( .CLK(n5281), .C(n5282) );
  CKBD0 U5165 ( .CLK(n5282), .C(n5283) );
  CKBD0 U5166 ( .CLK(n5283), .C(n5284) );
  CKBD0 U5167 ( .CLK(n5284), .C(n5285) );
  CKBD0 U5168 ( .CLK(n5285), .C(n5286) );
  CKBD0 U5169 ( .CLK(n5286), .C(n5287) );
  CKBD0 U5170 ( .CLK(n5287), .C(n5288) );
  CKBD0 U5171 ( .CLK(n5288), .C(n5289) );
  CKBD0 U5172 ( .CLK(n5289), .C(n5290) );
  BUFFD0 U5173 ( .I(n5290), .Z(n5291) );
  CKBD0 U5174 ( .CLK(n5291), .C(n5292) );
  CKBD0 U5175 ( .CLK(n5292), .C(n5293) );
  CKBD0 U5176 ( .CLK(n5293), .C(n5294) );
  CKBD0 U5177 ( .CLK(n5294), .C(n5295) );
  CKBD0 U5178 ( .CLK(n5295), .C(n5296) );
  CKBD0 U5179 ( .CLK(n5296), .C(n5297) );
  CKBD0 U5180 ( .CLK(n5297), .C(n5298) );
  CKBD0 U5181 ( .CLK(n5298), .C(n5299) );
  CKBD0 U5182 ( .CLK(n5299), .C(n5300) );
  BUFFD0 U5183 ( .I(n5300), .Z(n5301) );
  CKBD0 U5184 ( .CLK(n5301), .C(n5302) );
  CKBD0 U5185 ( .CLK(n5302), .C(n5303) );
  CKBD0 U5186 ( .CLK(n5303), .C(n5304) );
  CKBD0 U5187 ( .CLK(n5304), .C(n5305) );
  CKBD0 U5188 ( .CLK(n5305), .C(n5306) );
  CKBD0 U5189 ( .CLK(n5306), .C(n5307) );
  CKBD0 U5190 ( .CLK(n5307), .C(n5308) );
  CKBD0 U5191 ( .CLK(n5308), .C(n5309) );
  CKBD0 U5192 ( .CLK(n5309), .C(n5310) );
  BUFFD0 U5193 ( .I(n5310), .Z(n5311) );
  CKBD0 U5194 ( .CLK(n5311), .C(n5312) );
  CKBD0 U5195 ( .CLK(n5312), .C(n5313) );
  CKBD0 U5196 ( .CLK(n5313), .C(n5314) );
  CKBD0 U5197 ( .CLK(n5314), .C(n5315) );
  CKBD0 U5198 ( .CLK(n5315), .C(n5316) );
  CKBD0 U5199 ( .CLK(n5316), .C(n5317) );
  CKBD0 U5200 ( .CLK(n5317), .C(n5318) );
  CKBD0 U5201 ( .CLK(n5318), .C(n5319) );
  CKBD0 U5202 ( .CLK(n5319), .C(n5320) );
  CKBD0 U5203 ( .CLK(n5320), .C(n5321) );
  CKBD0 U5204 ( .CLK(n5321), .C(n5322) );
  BUFFD0 U5205 ( .I(n5322), .Z(n5323) );
  CKBD0 U5206 ( .CLK(n5323), .C(n5324) );
  CKBD0 U5207 ( .CLK(n5324), .C(n5325) );
  CKBD0 U5208 ( .CLK(n5325), .C(n5326) );
  CKBD0 U5209 ( .CLK(n5326), .C(n5327) );
  CKBD0 U5210 ( .CLK(n5327), .C(n5328) );
  CKBD0 U5211 ( .CLK(n5328), .C(n5329) );
  CKBD0 U5212 ( .CLK(n5329), .C(n5330) );
  CKBD0 U5213 ( .CLK(n5330), .C(n5331) );
  CKBD0 U5214 ( .CLK(n5331), .C(n5332) );
  CKBD0 U5215 ( .CLK(n5332), .C(n5333) );
  BUFFD0 U5216 ( .I(n5333), .Z(n5334) );
  CKBD0 U5217 ( .CLK(n5334), .C(n5335) );
  CKBD0 U5218 ( .CLK(n5335), .C(n5336) );
  CKBD0 U5219 ( .CLK(n5336), .C(n5337) );
  CKBD0 U5220 ( .CLK(n5337), .C(n5338) );
  CKBD0 U5221 ( .CLK(n5338), .C(n5339) );
  BUFFD0 U5222 ( .I(n5339), .Z(n5340) );
  CKBD0 U5223 ( .CLK(n5340), .C(n5341) );
  BUFFD0 U5224 ( .I(n5341), .Z(n5342) );
  CKBD0 U5225 ( .CLK(n5342), .C(n5343) );
  BUFFD0 U5226 ( .I(n5343), .Z(n5344) );
  CKBD0 U5227 ( .CLK(n5344), .C(n5345) );
  BUFFD0 U5228 ( .I(n5345), .Z(n5346) );
  CKBD0 U5229 ( .CLK(n5346), .C(n5347) );
  BUFFD0 U5230 ( .I(n5347), .Z(n5348) );
  CKBD0 U5231 ( .CLK(n5348), .C(n5349) );
  BUFFD0 U5232 ( .I(n5349), .Z(n5350) );
  CKBD0 U5233 ( .CLK(n5350), .C(n5351) );
  BUFFD0 U5234 ( .I(n5351), .Z(n5352) );
  CKBD0 U5235 ( .CLK(n5352), .C(n5353) );
  BUFFD0 U5236 ( .I(n5353), .Z(n5354) );
  BUFFD0 U5237 ( .I(n5356), .Z(n5355) );
  BUFFD0 U5238 ( .I(n5357), .Z(n5356) );
  BUFFD0 U5239 ( .I(n5358), .Z(n5357) );
  BUFFD0 U5240 ( .I(n142), .Z(n5358) );
  CKBD0 U5241 ( .CLK(n1053), .C(n5359) );
  CKBD0 U5242 ( .CLK(n5359), .C(n5360) );
  CKBD0 U5243 ( .CLK(n5360), .C(n5361) );
  CKBD0 U5244 ( .CLK(n5361), .C(n5362) );
  BUFFD0 U5245 ( .I(n5362), .Z(n5363) );
  CKBD0 U5246 ( .CLK(n5363), .C(n5364) );
  CKBD0 U5247 ( .CLK(n5364), .C(n5365) );
  CKBD0 U5248 ( .CLK(n5365), .C(n5366) );
  CKBD0 U5249 ( .CLK(n5366), .C(n5367) );
  CKBD0 U5250 ( .CLK(n5367), .C(n5368) );
  CKBD0 U5251 ( .CLK(n5368), .C(n5369) );
  CKBD0 U5252 ( .CLK(n5369), .C(n5370) );
  CKBD0 U5253 ( .CLK(n5370), .C(n5371) );
  CKBD0 U5254 ( .CLK(n5371), .C(n5372) );
  BUFFD0 U5255 ( .I(n5372), .Z(n5373) );
  CKBD0 U5256 ( .CLK(n5373), .C(n5374) );
  CKBD0 U5257 ( .CLK(n5374), .C(n5375) );
  CKBD0 U5258 ( .CLK(n5375), .C(n5376) );
  CKBD0 U5259 ( .CLK(n5376), .C(n5377) );
  CKBD0 U5260 ( .CLK(n5377), .C(n5378) );
  CKBD0 U5261 ( .CLK(n5378), .C(n5379) );
  CKBD0 U5262 ( .CLK(n5379), .C(n5380) );
  CKBD0 U5263 ( .CLK(n5380), .C(n5381) );
  CKBD0 U5264 ( .CLK(n5381), .C(n5382) );
  CKBD0 U5265 ( .CLK(n5382), .C(n5383) );
  BUFFD0 U5266 ( .I(n5383), .Z(n5384) );
  CKBD0 U5267 ( .CLK(n5384), .C(n5385) );
  CKBD0 U5268 ( .CLK(n5385), .C(n5386) );
  CKBD0 U5269 ( .CLK(n5386), .C(n5387) );
  CKBD0 U5270 ( .CLK(n5387), .C(n5388) );
  CKBD0 U5271 ( .CLK(n5388), .C(n5389) );
  CKBD0 U5272 ( .CLK(n5389), .C(n5390) );
  CKBD0 U5273 ( .CLK(n5390), .C(n5391) );
  CKBD0 U5274 ( .CLK(n5391), .C(n5392) );
  CKBD0 U5275 ( .CLK(n5392), .C(n5393) );
  CKBD0 U5276 ( .CLK(n5393), .C(n5394) );
  BUFFD0 U5277 ( .I(n5394), .Z(n5395) );
  CKBD0 U5278 ( .CLK(n5395), .C(n5396) );
  CKBD0 U5279 ( .CLK(n5396), .C(n5397) );
  CKBD0 U5280 ( .CLK(n5397), .C(n5398) );
  CKBD0 U5281 ( .CLK(n5398), .C(n5399) );
  CKBD0 U5282 ( .CLK(n5399), .C(n5400) );
  CKBD0 U5283 ( .CLK(n5400), .C(n5401) );
  CKBD0 U5284 ( .CLK(n5401), .C(n5402) );
  CKBD0 U5285 ( .CLK(n5402), .C(n5403) );
  CKBD0 U5286 ( .CLK(n5403), .C(n5404) );
  CKBD0 U5287 ( .CLK(n5404), .C(n5405) );
  BUFFD0 U5288 ( .I(n5405), .Z(n5406) );
  CKBD0 U5289 ( .CLK(n5406), .C(n5407) );
  CKBD0 U5290 ( .CLK(n5407), .C(n5408) );
  CKBD0 U5291 ( .CLK(n5408), .C(n5409) );
  CKBD0 U5292 ( .CLK(n5409), .C(n5410) );
  CKBD0 U5293 ( .CLK(n5410), .C(n5411) );
  CKBD0 U5294 ( .CLK(n5411), .C(n5412) );
  CKBD0 U5295 ( .CLK(n5412), .C(n5413) );
  CKBD0 U5296 ( .CLK(n5413), .C(n5414) );
  CKBD0 U5297 ( .CLK(n5414), .C(n5415) );
  BUFFD0 U5298 ( .I(n5415), .Z(n5416) );
  CKBD0 U5299 ( .CLK(n5416), .C(n5417) );
  CKBD0 U5300 ( .CLK(n5417), .C(n5418) );
  CKBD0 U5301 ( .CLK(n5418), .C(n5419) );
  CKBD0 U5302 ( .CLK(n5419), .C(n5420) );
  CKBD0 U5303 ( .CLK(n5420), .C(n5421) );
  CKBD0 U5304 ( .CLK(n5421), .C(n5422) );
  CKBD0 U5305 ( .CLK(n5422), .C(n5423) );
  CKBD0 U5306 ( .CLK(n5423), .C(n5424) );
  CKBD0 U5307 ( .CLK(n5424), .C(n5425) );
  CKBD0 U5308 ( .CLK(n5425), .C(n5426) );
  CKBD0 U5309 ( .CLK(n5426), .C(n5427) );
  BUFFD0 U5310 ( .I(n5427), .Z(n5428) );
  CKBD0 U5311 ( .CLK(n5428), .C(n5429) );
  CKBD0 U5312 ( .CLK(n5429), .C(n5430) );
  CKBD0 U5313 ( .CLK(n5430), .C(n5431) );
  CKBD0 U5314 ( .CLK(n5431), .C(n5432) );
  CKBD0 U5315 ( .CLK(n5432), .C(n5433) );
  CKBD0 U5316 ( .CLK(n5433), .C(n5434) );
  CKBD0 U5317 ( .CLK(n5434), .C(n5435) );
  CKBD0 U5318 ( .CLK(n5435), .C(n5436) );
  CKBD0 U5319 ( .CLK(n5436), .C(n5437) );
  BUFFD0 U5320 ( .I(n5437), .Z(n5438) );
  CKBD0 U5321 ( .CLK(n5438), .C(n5439) );
  CKBD0 U5322 ( .CLK(n5439), .C(n5440) );
  CKBD0 U5323 ( .CLK(n5440), .C(n5441) );
  CKBD0 U5324 ( .CLK(n5441), .C(n5442) );
  CKBD0 U5325 ( .CLK(n5442), .C(n5443) );
  CKBD0 U5326 ( .CLK(n5443), .C(n5444) );
  CKBD0 U5327 ( .CLK(n5444), .C(n5445) );
  CKBD0 U5328 ( .CLK(n5445), .C(n5446) );
  CKBD0 U5329 ( .CLK(n5446), .C(n5447) );
  CKBD0 U5330 ( .CLK(n5447), .C(n5448) );
  BUFFD0 U5331 ( .I(n5448), .Z(n5449) );
  CKBD0 U5332 ( .CLK(n5449), .C(n5450) );
  CKBD0 U5333 ( .CLK(n5450), .C(n5451) );
  CKBD0 U5334 ( .CLK(n5451), .C(n5452) );
  CKBD0 U5335 ( .CLK(n5452), .C(n5453) );
  CKBD0 U5336 ( .CLK(n5453), .C(n5454) );
  CKBD0 U5337 ( .CLK(n5454), .C(n5455) );
  CKBD0 U5338 ( .CLK(n5455), .C(n5456) );
  CKBD0 U5339 ( .CLK(n5456), .C(n5457) );
  CKBD0 U5340 ( .CLK(n5457), .C(n5458) );
  CKBD0 U5341 ( .CLK(n5458), .C(n5459) );
  BUFFD0 U5342 ( .I(n5459), .Z(n5460) );
  CKBD0 U5343 ( .CLK(n5460), .C(n5461) );
  CKBD0 U5344 ( .CLK(n5461), .C(n5462) );
  CKBD0 U5345 ( .CLK(n5462), .C(n5463) );
  CKBD0 U5346 ( .CLK(n5463), .C(n5464) );
  CKBD0 U5347 ( .CLK(n5464), .C(n5465) );
  CKBD0 U5348 ( .CLK(n5465), .C(n5466) );
  CKBD0 U5349 ( .CLK(n5466), .C(n5467) );
  CKBD0 U5350 ( .CLK(n5467), .C(n5468) );
  CKBD0 U5351 ( .CLK(n5468), .C(n5469) );
  CKBD0 U5352 ( .CLK(n5469), .C(n5470) );
  BUFFD0 U5353 ( .I(n5470), .Z(n5471) );
  CKBD0 U5354 ( .CLK(n5471), .C(n5472) );
  CKBD0 U5355 ( .CLK(n5472), .C(n5473) );
  CKBD0 U5356 ( .CLK(n5473), .C(n5474) );
  CKBD0 U5357 ( .CLK(n5474), .C(n5475) );
  CKBD0 U5358 ( .CLK(n5475), .C(n5476) );
  BUFFD0 U5359 ( .I(n5476), .Z(n5477) );
  CKBD0 U5360 ( .CLK(n5477), .C(n5478) );
  BUFFD0 U5361 ( .I(n5478), .Z(n5479) );
  CKBD0 U5362 ( .CLK(n5479), .C(n5480) );
  BUFFD0 U5363 ( .I(n5480), .Z(n5481) );
  CKBD0 U5364 ( .CLK(n5481), .C(n5482) );
  BUFFD0 U5365 ( .I(n5482), .Z(n5483) );
  CKBD0 U5366 ( .CLK(n5483), .C(n5484) );
  BUFFD0 U5367 ( .I(n5484), .Z(n5485) );
  CKBD0 U5368 ( .CLK(n5485), .C(n5486) );
  BUFFD0 U5369 ( .I(n5486), .Z(n5487) );
  CKBD0 U5370 ( .CLK(n5487), .C(n5488) );
  BUFFD0 U5371 ( .I(n5488), .Z(n5489) );
  CKBD0 U5372 ( .CLK(n5489), .C(n5490) );
  BUFFD0 U5373 ( .I(n5490), .Z(n5491) );
  BUFFD0 U5374 ( .I(n5493), .Z(n5492) );
  BUFFD0 U5375 ( .I(n5494), .Z(n5493) );
  BUFFD0 U5376 ( .I(n5495), .Z(n5494) );
  BUFFD0 U5377 ( .I(n141), .Z(n5495) );
  CKBD0 U5378 ( .CLK(n1051), .C(n5496) );
  CKBD0 U5379 ( .CLK(n5496), .C(n5497) );
  CKBD0 U5380 ( .CLK(n5497), .C(n5498) );
  BUFFD0 U5381 ( .I(n5498), .Z(n5499) );
  CKBD0 U5382 ( .CLK(n5499), .C(n5500) );
  CKBD0 U5383 ( .CLK(n5500), .C(n5501) );
  CKBD0 U5384 ( .CLK(n5501), .C(n5502) );
  CKBD0 U5385 ( .CLK(n5502), .C(n5503) );
  CKBD0 U5386 ( .CLK(n5503), .C(n5504) );
  CKBD0 U5387 ( .CLK(n5504), .C(n5505) );
  CKBD0 U5388 ( .CLK(n5505), .C(n5506) );
  CKBD0 U5389 ( .CLK(n5506), .C(n5507) );
  CKBD0 U5390 ( .CLK(n5507), .C(n5508) );
  CKBD0 U5391 ( .CLK(n5508), .C(n5509) );
  BUFFD0 U5392 ( .I(n5509), .Z(n5510) );
  CKBD0 U5393 ( .CLK(n5510), .C(n5511) );
  CKBD0 U5394 ( .CLK(n5511), .C(n5512) );
  CKBD0 U5395 ( .CLK(n5512), .C(n5513) );
  CKBD0 U5396 ( .CLK(n5513), .C(n5514) );
  CKBD0 U5397 ( .CLK(n5514), .C(n5515) );
  CKBD0 U5398 ( .CLK(n5515), .C(n5516) );
  CKBD0 U5399 ( .CLK(n5516), .C(n5517) );
  CKBD0 U5400 ( .CLK(n5517), .C(n5518) );
  CKBD0 U5401 ( .CLK(n5518), .C(n5519) );
  CKBD0 U5402 ( .CLK(n5519), .C(n5520) );
  BUFFD0 U5403 ( .I(n5520), .Z(n5521) );
  CKBD0 U5404 ( .CLK(n5521), .C(n5522) );
  CKBD0 U5405 ( .CLK(n5522), .C(n5523) );
  CKBD0 U5406 ( .CLK(n5523), .C(n5524) );
  CKBD0 U5407 ( .CLK(n5524), .C(n5525) );
  CKBD0 U5408 ( .CLK(n5525), .C(n5526) );
  CKBD0 U5409 ( .CLK(n5526), .C(n5527) );
  CKBD0 U5410 ( .CLK(n5527), .C(n5528) );
  CKBD0 U5411 ( .CLK(n5528), .C(n5529) );
  CKBD0 U5412 ( .CLK(n5529), .C(n5530) );
  BUFFD0 U5413 ( .I(n5530), .Z(n5531) );
  CKBD0 U5414 ( .CLK(n5531), .C(n5532) );
  CKBD0 U5415 ( .CLK(n5532), .C(n5533) );
  CKBD0 U5416 ( .CLK(n5533), .C(n5534) );
  CKBD0 U5417 ( .CLK(n5534), .C(n5535) );
  CKBD0 U5418 ( .CLK(n5535), .C(n5536) );
  CKBD0 U5419 ( .CLK(n5536), .C(n5537) );
  CKBD0 U5420 ( .CLK(n5537), .C(n5538) );
  CKBD0 U5421 ( .CLK(n5538), .C(n5539) );
  CKBD0 U5422 ( .CLK(n5539), .C(n5540) );
  CKBD0 U5423 ( .CLK(n5540), .C(n5541) );
  CKBD0 U5424 ( .CLK(n5541), .C(n5542) );
  BUFFD0 U5425 ( .I(n5542), .Z(n5543) );
  CKBD0 U5426 ( .CLK(n5543), .C(n5544) );
  CKBD0 U5427 ( .CLK(n5544), .C(n5545) );
  CKBD0 U5428 ( .CLK(n5545), .C(n5546) );
  CKBD0 U5429 ( .CLK(n5546), .C(n5547) );
  CKBD0 U5430 ( .CLK(n5547), .C(n5548) );
  CKBD0 U5431 ( .CLK(n5548), .C(n5549) );
  CKBD0 U5432 ( .CLK(n5549), .C(n5550) );
  CKBD0 U5433 ( .CLK(n5550), .C(n5551) );
  CKBD0 U5434 ( .CLK(n5551), .C(n5552) );
  CKBD0 U5435 ( .CLK(n5552), .C(n5553) );
  BUFFD0 U5436 ( .I(n5553), .Z(n5554) );
  CKBD0 U5437 ( .CLK(n5554), .C(n5555) );
  CKBD0 U5438 ( .CLK(n5555), .C(n5556) );
  CKBD0 U5439 ( .CLK(n5556), .C(n5557) );
  CKBD0 U5440 ( .CLK(n5557), .C(n5558) );
  CKBD0 U5441 ( .CLK(n5558), .C(n5559) );
  CKBD0 U5442 ( .CLK(n5559), .C(n5560) );
  CKBD0 U5443 ( .CLK(n5560), .C(n5561) );
  CKBD0 U5444 ( .CLK(n5561), .C(n5562) );
  CKBD0 U5445 ( .CLK(n5562), .C(n5563) );
  BUFFD0 U5446 ( .I(n5563), .Z(n5564) );
  CKBD0 U5447 ( .CLK(n5564), .C(n5565) );
  CKBD0 U5448 ( .CLK(n5565), .C(n5566) );
  CKBD0 U5449 ( .CLK(n5566), .C(n5567) );
  CKBD0 U5450 ( .CLK(n5567), .C(n5568) );
  CKBD0 U5451 ( .CLK(n5568), .C(n5569) );
  CKBD0 U5452 ( .CLK(n5569), .C(n5570) );
  CKBD0 U5453 ( .CLK(n5570), .C(n5571) );
  CKBD0 U5454 ( .CLK(n5571), .C(n5572) );
  CKBD0 U5455 ( .CLK(n5572), .C(n5573) );
  CKBD0 U5456 ( .CLK(n5573), .C(n5574) );
  CKBD0 U5457 ( .CLK(n5574), .C(n5575) );
  BUFFD0 U5458 ( .I(n5575), .Z(n5576) );
  CKBD0 U5459 ( .CLK(n5576), .C(n5577) );
  CKBD0 U5460 ( .CLK(n5577), .C(n5578) );
  CKBD0 U5461 ( .CLK(n5578), .C(n5579) );
  CKBD0 U5462 ( .CLK(n5579), .C(n5580) );
  CKBD0 U5463 ( .CLK(n5580), .C(n5581) );
  CKBD0 U5464 ( .CLK(n5581), .C(n5582) );
  CKBD0 U5465 ( .CLK(n5582), .C(n5583) );
  CKBD0 U5466 ( .CLK(n5583), .C(n5584) );
  CKBD0 U5467 ( .CLK(n5584), .C(n5585) );
  BUFFD0 U5468 ( .I(n5585), .Z(n5586) );
  CKBD0 U5469 ( .CLK(n5586), .C(n5587) );
  CKBD0 U5470 ( .CLK(n5587), .C(n5588) );
  CKBD0 U5471 ( .CLK(n5588), .C(n5589) );
  CKBD0 U5472 ( .CLK(n5589), .C(n5590) );
  CKBD0 U5473 ( .CLK(n5590), .C(n5591) );
  CKBD0 U5474 ( .CLK(n5591), .C(n5592) );
  CKBD0 U5475 ( .CLK(n5592), .C(n5593) );
  CKBD0 U5476 ( .CLK(n5593), .C(n5594) );
  CKBD0 U5477 ( .CLK(n5594), .C(n5595) );
  BUFFD0 U5478 ( .I(n5595), .Z(n5596) );
  CKBD0 U5479 ( .CLK(n5596), .C(n5597) );
  CKBD0 U5480 ( .CLK(n5597), .C(n5598) );
  CKBD0 U5481 ( .CLK(n5598), .C(n5599) );
  CKBD0 U5482 ( .CLK(n5599), .C(n5600) );
  CKBD0 U5483 ( .CLK(n5600), .C(n5601) );
  CKBD0 U5484 ( .CLK(n5601), .C(n5602) );
  CKBD0 U5485 ( .CLK(n5602), .C(n5603) );
  CKBD0 U5486 ( .CLK(n5603), .C(n5604) );
  CKBD0 U5487 ( .CLK(n5604), .C(n5605) );
  CKBD0 U5488 ( .CLK(n5605), .C(n5606) );
  CKBD0 U5489 ( .CLK(n5606), .C(n5607) );
  BUFFD0 U5490 ( .I(n5607), .Z(n5608) );
  CKBD0 U5491 ( .CLK(n5608), .C(n5609) );
  CKBD0 U5492 ( .CLK(n5609), .C(n5610) );
  CKBD0 U5493 ( .CLK(n5610), .C(n5611) );
  CKBD0 U5494 ( .CLK(n5611), .C(n5612) );
  CKBD0 U5495 ( .CLK(n5612), .C(n5613) );
  BUFFD0 U5496 ( .I(n5613), .Z(n5614) );
  CKBD0 U5497 ( .CLK(n5614), .C(n5615) );
  BUFFD0 U5498 ( .I(n5615), .Z(n5616) );
  CKBD0 U5499 ( .CLK(n5616), .C(n5617) );
  BUFFD0 U5500 ( .I(n5617), .Z(n5618) );
  CKBD0 U5501 ( .CLK(n5618), .C(n5619) );
  BUFFD0 U5502 ( .I(n5619), .Z(n5620) );
  CKBD0 U5503 ( .CLK(n5620), .C(n5621) );
  BUFFD0 U5504 ( .I(n5621), .Z(n5622) );
  CKBD0 U5505 ( .CLK(n5622), .C(n5623) );
  BUFFD0 U5506 ( .I(n5623), .Z(n5624) );
  CKBD0 U5507 ( .CLK(n5624), .C(n5625) );
  BUFFD0 U5508 ( .I(n5625), .Z(n5626) );
  CKBD0 U5509 ( .CLK(n5626), .C(n5627) );
  BUFFD0 U5510 ( .I(n5627), .Z(n5628) );
  BUFFD0 U5511 ( .I(n5630), .Z(n5629) );
  BUFFD0 U5512 ( .I(n5631), .Z(n5630) );
  BUFFD0 U5513 ( .I(n140), .Z(n5631) );
  CKBD0 U5514 ( .CLK(n2363), .C(n5632) );
  CKBD0 U5515 ( .CLK(n5632), .C(n5633) );
  CKBD0 U5516 ( .CLK(n5633), .C(n5634) );
  BUFFD0 U5517 ( .I(n5634), .Z(n5635) );
  CKBD0 U5518 ( .CLK(n5635), .C(n5636) );
  CKBD0 U5519 ( .CLK(n5636), .C(n5637) );
  CKBD0 U5520 ( .CLK(n5637), .C(n5638) );
  CKBD0 U5521 ( .CLK(n5638), .C(n5639) );
  CKBD0 U5522 ( .CLK(n5639), .C(n5640) );
  CKBD0 U5523 ( .CLK(n5640), .C(n5641) );
  CKBD0 U5524 ( .CLK(n5641), .C(n5642) );
  CKBD0 U5525 ( .CLK(n5642), .C(n5643) );
  CKBD0 U5526 ( .CLK(n5643), .C(n5644) );
  CKBD0 U5527 ( .CLK(n5644), .C(n5645) );
  BUFFD0 U5528 ( .I(n5645), .Z(n5646) );
  CKBD0 U5529 ( .CLK(n5646), .C(n5647) );
  CKBD0 U5530 ( .CLK(n5647), .C(n5648) );
  CKBD0 U5531 ( .CLK(n5648), .C(n5649) );
  CKBD0 U5532 ( .CLK(n5649), .C(n5650) );
  CKBD0 U5533 ( .CLK(n5650), .C(n5651) );
  CKBD0 U5534 ( .CLK(n5651), .C(n5652) );
  CKBD0 U5535 ( .CLK(n5652), .C(n5653) );
  CKBD0 U5536 ( .CLK(n5653), .C(n5654) );
  CKBD0 U5537 ( .CLK(n5654), .C(n5655) );
  CKBD0 U5538 ( .CLK(n5655), .C(n5656) );
  BUFFD0 U5539 ( .I(n5656), .Z(n5657) );
  CKBD0 U5540 ( .CLK(n5657), .C(n5658) );
  CKBD0 U5541 ( .CLK(n5658), .C(n5659) );
  CKBD0 U5542 ( .CLK(n5659), .C(n5660) );
  CKBD0 U5543 ( .CLK(n5660), .C(n5661) );
  CKBD0 U5544 ( .CLK(n5661), .C(n5662) );
  CKBD0 U5545 ( .CLK(n5662), .C(n5663) );
  CKBD0 U5546 ( .CLK(n5663), .C(n5664) );
  CKBD0 U5547 ( .CLK(n5664), .C(n5665) );
  CKBD0 U5548 ( .CLK(n5665), .C(n5666) );
  BUFFD0 U5549 ( .I(n5666), .Z(n5667) );
  CKBD0 U5550 ( .CLK(n5667), .C(n5668) );
  CKBD0 U5551 ( .CLK(n5668), .C(n5669) );
  CKBD0 U5552 ( .CLK(n5669), .C(n5670) );
  CKBD0 U5553 ( .CLK(n5670), .C(n5671) );
  CKBD0 U5554 ( .CLK(n5671), .C(n5672) );
  CKBD0 U5555 ( .CLK(n5672), .C(n5673) );
  CKBD0 U5556 ( .CLK(n5673), .C(n5674) );
  CKBD0 U5557 ( .CLK(n5674), .C(n5675) );
  CKBD0 U5558 ( .CLK(n5675), .C(n5676) );
  CKBD0 U5559 ( .CLK(n5676), .C(n5677) );
  CKBD0 U5560 ( .CLK(n5677), .C(n5678) );
  BUFFD0 U5561 ( .I(n5678), .Z(n5679) );
  CKBD0 U5562 ( .CLK(n5679), .C(n5680) );
  CKBD0 U5563 ( .CLK(n5680), .C(n5681) );
  CKBD0 U5564 ( .CLK(n5681), .C(n5682) );
  CKBD0 U5565 ( .CLK(n5682), .C(n5683) );
  CKBD0 U5566 ( .CLK(n5683), .C(n5684) );
  CKBD0 U5567 ( .CLK(n5684), .C(n5685) );
  CKBD0 U5568 ( .CLK(n5685), .C(n5686) );
  CKBD0 U5569 ( .CLK(n5686), .C(n5687) );
  CKBD0 U5570 ( .CLK(n5687), .C(n5688) );
  BUFFD0 U5571 ( .I(n5688), .Z(n5689) );
  CKBD0 U5572 ( .CLK(n5689), .C(n5690) );
  CKBD0 U5573 ( .CLK(n5690), .C(n5691) );
  CKBD0 U5574 ( .CLK(n5691), .C(n5692) );
  CKBD0 U5575 ( .CLK(n5692), .C(n5693) );
  CKBD0 U5576 ( .CLK(n5693), .C(n5694) );
  CKBD0 U5577 ( .CLK(n5694), .C(n5695) );
  CKBD0 U5578 ( .CLK(n5695), .C(n5696) );
  CKBD0 U5579 ( .CLK(n5696), .C(n5697) );
  CKBD0 U5580 ( .CLK(n5697), .C(n5698) );
  CKBD0 U5581 ( .CLK(n5698), .C(n5699) );
  BUFFD0 U5582 ( .I(n5699), .Z(n5700) );
  CKBD0 U5583 ( .CLK(n5700), .C(n5701) );
  CKBD0 U5584 ( .CLK(n5701), .C(n5702) );
  CKBD0 U5585 ( .CLK(n5702), .C(n5703) );
  CKBD0 U5586 ( .CLK(n5703), .C(n5704) );
  CKBD0 U5587 ( .CLK(n5704), .C(n5705) );
  CKBD0 U5588 ( .CLK(n5705), .C(n5706) );
  CKBD0 U5589 ( .CLK(n5706), .C(n5707) );
  CKBD0 U5590 ( .CLK(n5707), .C(n5708) );
  CKBD0 U5591 ( .CLK(n5708), .C(n5709) );
  CKBD0 U5592 ( .CLK(n5709), .C(n5710) );
  BUFFD0 U5593 ( .I(n5710), .Z(n5711) );
  CKBD0 U5594 ( .CLK(n5711), .C(n5712) );
  CKBD0 U5595 ( .CLK(n5712), .C(n5713) );
  CKBD0 U5596 ( .CLK(n5713), .C(n5714) );
  CKBD0 U5597 ( .CLK(n5714), .C(n5715) );
  CKBD0 U5598 ( .CLK(n5715), .C(n5716) );
  CKBD0 U5599 ( .CLK(n5716), .C(n5717) );
  CKBD0 U5600 ( .CLK(n5717), .C(n5718) );
  CKBD0 U5601 ( .CLK(n5718), .C(n5719) );
  CKBD0 U5602 ( .CLK(n5719), .C(n5720) );
  CKBD0 U5603 ( .CLK(n5720), .C(n5721) );
  BUFFD0 U5604 ( .I(n5721), .Z(n5722) );
  CKBD0 U5605 ( .CLK(n5722), .C(n5723) );
  CKBD0 U5606 ( .CLK(n5723), .C(n5724) );
  CKBD0 U5607 ( .CLK(n5724), .C(n5725) );
  CKBD0 U5608 ( .CLK(n5725), .C(n5726) );
  CKBD0 U5609 ( .CLK(n5726), .C(n5727) );
  CKBD0 U5610 ( .CLK(n5727), .C(n5728) );
  CKBD0 U5611 ( .CLK(n5728), .C(n5729) );
  CKBD0 U5612 ( .CLK(n5729), .C(n5730) );
  CKBD0 U5613 ( .CLK(n5730), .C(n5731) );
  CKBD0 U5614 ( .CLK(n5731), .C(n5732) );
  BUFFD0 U5615 ( .I(n5732), .Z(n5733) );
  CKBD0 U5616 ( .CLK(n5733), .C(n5734) );
  CKBD0 U5617 ( .CLK(n5734), .C(n5735) );
  CKBD0 U5618 ( .CLK(n5735), .C(n5736) );
  CKBD0 U5619 ( .CLK(n5736), .C(n5737) );
  CKBD0 U5620 ( .CLK(n5737), .C(n5738) );
  CKBD0 U5621 ( .CLK(n5738), .C(n5739) );
  CKBD0 U5622 ( .CLK(n5739), .C(n5740) );
  CKBD0 U5623 ( .CLK(n5740), .C(n5741) );
  CKBD0 U5624 ( .CLK(n5741), .C(n5742) );
  CKBD0 U5625 ( .CLK(n5742), .C(n5743) );
  BUFFD0 U5626 ( .I(n5743), .Z(n5744) );
  CKBD0 U5627 ( .CLK(n5744), .C(n5745) );
  CKBD0 U5628 ( .CLK(n5745), .C(n5746) );
  CKBD0 U5629 ( .CLK(n5746), .C(n5747) );
  CKBD0 U5630 ( .CLK(n5747), .C(n5748) );
  CKBD0 U5631 ( .CLK(n5748), .C(n5749) );
  BUFFD0 U5632 ( .I(n5749), .Z(n5750) );
  CKBD0 U5633 ( .CLK(n5750), .C(n5751) );
  BUFFD0 U5634 ( .I(n5751), .Z(n5752) );
  CKBD0 U5635 ( .CLK(n5752), .C(n5753) );
  BUFFD0 U5636 ( .I(n5753), .Z(n5754) );
  CKBD0 U5637 ( .CLK(n5754), .C(n5755) );
  BUFFD0 U5638 ( .I(n5755), .Z(n5756) );
  CKBD0 U5639 ( .CLK(n5756), .C(n5757) );
  BUFFD0 U5640 ( .I(n5757), .Z(n5758) );
  CKBD0 U5641 ( .CLK(n5758), .C(n5759) );
  BUFFD0 U5642 ( .I(n5759), .Z(n5760) );
  CKBD0 U5643 ( .CLK(n5760), .C(n5761) );
  BUFFD0 U5644 ( .I(n5761), .Z(n5762) );
  CKBD0 U5645 ( .CLK(n5762), .C(n5763) );
  BUFFD0 U5646 ( .I(n5763), .Z(n5764) );
  BUFFD0 U5647 ( .I(n5766), .Z(n5765) );
  BUFFD0 U5648 ( .I(n5767), .Z(n5766) );
  BUFFD0 U5649 ( .I(n5768), .Z(n5767) );
  BUFFD0 U5650 ( .I(n139), .Z(n5768) );
  CKBD0 U5651 ( .CLK(n870), .C(n5769) );
  CKBD0 U5652 ( .CLK(n5769), .C(n5770) );
  CKBD0 U5653 ( .CLK(n5770), .C(n5771) );
  BUFFD0 U5654 ( .I(n5771), .Z(n5772) );
  CKBD0 U5655 ( .CLK(n5772), .C(n5773) );
  CKBD0 U5656 ( .CLK(n5773), .C(n5774) );
  CKBD0 U5657 ( .CLK(n5774), .C(n5775) );
  CKBD0 U5658 ( .CLK(n5775), .C(n5776) );
  CKBD0 U5659 ( .CLK(n5776), .C(n5777) );
  CKBD0 U5660 ( .CLK(n5777), .C(n5778) );
  CKBD0 U5661 ( .CLK(n5778), .C(n5779) );
  CKBD0 U5662 ( .CLK(n5779), .C(n5780) );
  CKBD0 U5663 ( .CLK(n5780), .C(n5781) );
  CKBD0 U5664 ( .CLK(n5781), .C(n5782) );
  BUFFD0 U5665 ( .I(n5782), .Z(n5783) );
  CKBD0 U5666 ( .CLK(n5783), .C(n5784) );
  CKBD0 U5667 ( .CLK(n5784), .C(n5785) );
  CKBD0 U5668 ( .CLK(n5785), .C(n5786) );
  CKBD0 U5669 ( .CLK(n5786), .C(n5787) );
  CKBD0 U5670 ( .CLK(n5787), .C(n5788) );
  CKBD0 U5671 ( .CLK(n5788), .C(n5789) );
  CKBD0 U5672 ( .CLK(n5789), .C(n5790) );
  CKBD0 U5673 ( .CLK(n5790), .C(n5791) );
  CKBD0 U5674 ( .CLK(n5791), .C(n5792) );
  CKBD0 U5675 ( .CLK(n5792), .C(n5793) );
  BUFFD0 U5676 ( .I(n5793), .Z(n5794) );
  CKBD0 U5677 ( .CLK(n5794), .C(n5795) );
  CKBD0 U5678 ( .CLK(n5795), .C(n5796) );
  CKBD0 U5679 ( .CLK(n5796), .C(n5797) );
  CKBD0 U5680 ( .CLK(n5797), .C(n5798) );
  CKBD0 U5681 ( .CLK(n5798), .C(n5799) );
  CKBD0 U5682 ( .CLK(n5799), .C(n5800) );
  CKBD0 U5683 ( .CLK(n5800), .C(n5801) );
  CKBD0 U5684 ( .CLK(n5801), .C(n5802) );
  CKBD0 U5685 ( .CLK(n5802), .C(n5803) );
  CKBD0 U5686 ( .CLK(n5803), .C(n5804) );
  BUFFD0 U5687 ( .I(n5804), .Z(n5805) );
  CKBD0 U5688 ( .CLK(n5805), .C(n5806) );
  CKBD0 U5689 ( .CLK(n5806), .C(n5807) );
  CKBD0 U5690 ( .CLK(n5807), .C(n5808) );
  CKBD0 U5691 ( .CLK(n5808), .C(n5809) );
  CKBD0 U5692 ( .CLK(n5809), .C(n5810) );
  CKBD0 U5693 ( .CLK(n5810), .C(n5811) );
  CKBD0 U5694 ( .CLK(n5811), .C(n5812) );
  CKBD0 U5695 ( .CLK(n5812), .C(n5813) );
  CKBD0 U5696 ( .CLK(n5813), .C(n5814) );
  BUFFD0 U5697 ( .I(n5814), .Z(n5815) );
  CKBD0 U5698 ( .CLK(n5815), .C(n5816) );
  CKBD0 U5699 ( .CLK(n5816), .C(n5817) );
  CKBD0 U5700 ( .CLK(n5817), .C(n5818) );
  CKBD0 U5701 ( .CLK(n5818), .C(n5819) );
  CKBD0 U5702 ( .CLK(n5819), .C(n5820) );
  CKBD0 U5703 ( .CLK(n5820), .C(n5821) );
  CKBD0 U5704 ( .CLK(n5821), .C(n5822) );
  CKBD0 U5705 ( .CLK(n5822), .C(n5823) );
  CKBD0 U5706 ( .CLK(n5823), .C(n5824) );
  CKBD0 U5707 ( .CLK(n5824), .C(n5825) );
  CKBD0 U5708 ( .CLK(n5825), .C(n5826) );
  BUFFD0 U5709 ( .I(n5826), .Z(n5827) );
  CKBD0 U5710 ( .CLK(n5827), .C(n5828) );
  CKBD0 U5711 ( .CLK(n5828), .C(n5829) );
  CKBD0 U5712 ( .CLK(n5829), .C(n5830) );
  CKBD0 U5713 ( .CLK(n5830), .C(n5831) );
  CKBD0 U5714 ( .CLK(n5831), .C(n5832) );
  CKBD0 U5715 ( .CLK(n5832), .C(n5833) );
  CKBD0 U5716 ( .CLK(n5833), .C(n5834) );
  CKBD0 U5717 ( .CLK(n5834), .C(n5835) );
  CKBD0 U5718 ( .CLK(n5835), .C(n5836) );
  BUFFD0 U5719 ( .I(n5836), .Z(n5837) );
  CKBD0 U5720 ( .CLK(n5837), .C(n5838) );
  CKBD0 U5721 ( .CLK(n5838), .C(n5839) );
  CKBD0 U5722 ( .CLK(n5839), .C(n5840) );
  CKBD0 U5723 ( .CLK(n5840), .C(n5841) );
  CKBD0 U5724 ( .CLK(n5841), .C(n5842) );
  CKBD0 U5725 ( .CLK(n5842), .C(n5843) );
  CKBD0 U5726 ( .CLK(n5843), .C(n5844) );
  CKBD0 U5727 ( .CLK(n5844), .C(n5845) );
  CKBD0 U5728 ( .CLK(n5845), .C(n5846) );
  CKBD0 U5729 ( .CLK(n5846), .C(n5847) );
  BUFFD0 U5730 ( .I(n5847), .Z(n5848) );
  CKBD0 U5731 ( .CLK(n5848), .C(n5849) );
  CKBD0 U5732 ( .CLK(n5849), .C(n5850) );
  CKBD0 U5733 ( .CLK(n5850), .C(n5851) );
  CKBD0 U5734 ( .CLK(n5851), .C(n5852) );
  CKBD0 U5735 ( .CLK(n5852), .C(n5853) );
  CKBD0 U5736 ( .CLK(n5853), .C(n5854) );
  CKBD0 U5737 ( .CLK(n5854), .C(n5855) );
  CKBD0 U5738 ( .CLK(n5855), .C(n5856) );
  CKBD0 U5739 ( .CLK(n5856), .C(n5857) );
  CKBD0 U5740 ( .CLK(n5857), .C(n5858) );
  BUFFD0 U5741 ( .I(n5858), .Z(n5859) );
  CKBD0 U5742 ( .CLK(n5859), .C(n5860) );
  CKBD0 U5743 ( .CLK(n5860), .C(n5861) );
  CKBD0 U5744 ( .CLK(n5861), .C(n5862) );
  CKBD0 U5745 ( .CLK(n5862), .C(n5863) );
  CKBD0 U5746 ( .CLK(n5863), .C(n5864) );
  CKBD0 U5747 ( .CLK(n5864), .C(n5865) );
  CKBD0 U5748 ( .CLK(n5865), .C(n5866) );
  CKBD0 U5749 ( .CLK(n5866), .C(n5867) );
  CKBD0 U5750 ( .CLK(n5867), .C(n5868) );
  CKBD0 U5751 ( .CLK(n5868), .C(n5869) );
  BUFFD0 U5752 ( .I(n5869), .Z(n5870) );
  CKBD0 U5753 ( .CLK(n5870), .C(n5871) );
  CKBD0 U5754 ( .CLK(n5871), .C(n5872) );
  CKBD0 U5755 ( .CLK(n5872), .C(n5873) );
  CKBD0 U5756 ( .CLK(n5873), .C(n5874) );
  CKBD0 U5757 ( .CLK(n5874), .C(n5875) );
  CKBD0 U5758 ( .CLK(n5875), .C(n5876) );
  CKBD0 U5759 ( .CLK(n5876), .C(n5877) );
  CKBD0 U5760 ( .CLK(n5877), .C(n5878) );
  CKBD0 U5761 ( .CLK(n5878), .C(n5879) );
  CKBD0 U5762 ( .CLK(n5879), .C(n5880) );
  BUFFD0 U5763 ( .I(n5880), .Z(n5881) );
  CKBD0 U5764 ( .CLK(n5881), .C(n5882) );
  CKBD0 U5765 ( .CLK(n5882), .C(n5883) );
  CKBD0 U5766 ( .CLK(n5883), .C(n5884) );
  CKBD0 U5767 ( .CLK(n5884), .C(n5885) );
  CKBD0 U5768 ( .CLK(n5885), .C(n5886) );
  BUFFD0 U5769 ( .I(n5886), .Z(n5887) );
  CKBD0 U5770 ( .CLK(n5887), .C(n5888) );
  BUFFD0 U5771 ( .I(n5888), .Z(n5889) );
  CKBD0 U5772 ( .CLK(n5889), .C(n5890) );
  BUFFD0 U5773 ( .I(n5890), .Z(n5891) );
  CKBD0 U5774 ( .CLK(n5891), .C(n5892) );
  BUFFD0 U5775 ( .I(n5892), .Z(n5893) );
  CKBD0 U5776 ( .CLK(n5893), .C(n5894) );
  BUFFD0 U5777 ( .I(n5894), .Z(n5895) );
  CKBD0 U5778 ( .CLK(n5895), .C(n5896) );
  BUFFD0 U5779 ( .I(n5896), .Z(n5897) );
  CKBD0 U5780 ( .CLK(n5897), .C(n5898) );
  BUFFD0 U5781 ( .I(n5898), .Z(n5899) );
  CKBD0 U5782 ( .CLK(n5899), .C(n5900) );
  BUFFD0 U5783 ( .I(n5900), .Z(n5901) );
  BUFFD0 U5784 ( .I(n138), .Z(n5902) );
  BUFFD0 U5785 ( .I(n5904), .Z(n5903) );
  BUFFD0 U5786 ( .I(n5905), .Z(n5904) );
  BUFFD0 U5787 ( .I(Decoder[5]), .Z(n5905) );
  CKBD0 U5788 ( .CLK(n868), .C(n5906) );
  CKBD0 U5789 ( .CLK(n5906), .C(n5907) );
  CKBD0 U5790 ( .CLK(n5907), .C(n5908) );
  CKBD0 U5791 ( .CLK(n5908), .C(n5909) );
  BUFFD0 U5792 ( .I(n5909), .Z(n5910) );
  CKBD0 U5793 ( .CLK(n5910), .C(n5911) );
  CKBD0 U5794 ( .CLK(n5911), .C(n5912) );
  CKBD0 U5795 ( .CLK(n5912), .C(n5913) );
  CKBD0 U5796 ( .CLK(n5913), .C(n5914) );
  CKBD0 U5797 ( .CLK(n5914), .C(n5915) );
  CKBD0 U5798 ( .CLK(n5915), .C(n5916) );
  CKBD0 U5799 ( .CLK(n5916), .C(n5917) );
  CKBD0 U5800 ( .CLK(n5917), .C(n5918) );
  CKBD0 U5801 ( .CLK(n5918), .C(n5919) );
  BUFFD0 U5802 ( .I(n5919), .Z(n5920) );
  CKBD0 U5803 ( .CLK(n5920), .C(n5921) );
  CKBD0 U5804 ( .CLK(n5921), .C(n5922) );
  CKBD0 U5805 ( .CLK(n5922), .C(n5923) );
  CKBD0 U5806 ( .CLK(n5923), .C(n5924) );
  CKBD0 U5807 ( .CLK(n5924), .C(n5925) );
  CKBD0 U5808 ( .CLK(n5925), .C(n5926) );
  CKBD0 U5809 ( .CLK(n5926), .C(n5927) );
  CKBD0 U5810 ( .CLK(n5927), .C(n5928) );
  CKBD0 U5811 ( .CLK(n5928), .C(n5929) );
  CKBD0 U5812 ( .CLK(n5929), .C(n5930) );
  BUFFD0 U5813 ( .I(n5930), .Z(n5931) );
  CKBD0 U5814 ( .CLK(n5931), .C(n5932) );
  CKBD0 U5815 ( .CLK(n5932), .C(n5933) );
  CKBD0 U5816 ( .CLK(n5933), .C(n5934) );
  CKBD0 U5817 ( .CLK(n5934), .C(n5935) );
  CKBD0 U5818 ( .CLK(n5935), .C(n5936) );
  CKBD0 U5819 ( .CLK(n5936), .C(n5937) );
  CKBD0 U5820 ( .CLK(n5937), .C(n5938) );
  CKBD0 U5821 ( .CLK(n5938), .C(n5939) );
  CKBD0 U5822 ( .CLK(n5939), .C(n5940) );
  CKBD0 U5823 ( .CLK(n5940), .C(n5941) );
  BUFFD0 U5824 ( .I(n5941), .Z(n5942) );
  CKBD0 U5825 ( .CLK(n5942), .C(n5943) );
  CKBD0 U5826 ( .CLK(n5943), .C(n5944) );
  CKBD0 U5827 ( .CLK(n5944), .C(n5945) );
  CKBD0 U5828 ( .CLK(n5945), .C(n5946) );
  CKBD0 U5829 ( .CLK(n5946), .C(n5947) );
  CKBD0 U5830 ( .CLK(n5947), .C(n5948) );
  CKBD0 U5831 ( .CLK(n5948), .C(n5949) );
  CKBD0 U5832 ( .CLK(n5949), .C(n5950) );
  CKBD0 U5833 ( .CLK(n5950), .C(n5951) );
  CKBD0 U5834 ( .CLK(n5951), .C(n5952) );
  BUFFD0 U5835 ( .I(n5952), .Z(n5953) );
  CKBD0 U5836 ( .CLK(n5953), .C(n5954) );
  CKBD0 U5837 ( .CLK(n5954), .C(n5955) );
  CKBD0 U5838 ( .CLK(n5955), .C(n5956) );
  CKBD0 U5839 ( .CLK(n5956), .C(n5957) );
  CKBD0 U5840 ( .CLK(n5957), .C(n5958) );
  CKBD0 U5841 ( .CLK(n5958), .C(n5959) );
  CKBD0 U5842 ( .CLK(n5959), .C(n5960) );
  CKBD0 U5843 ( .CLK(n5960), .C(n5961) );
  CKBD0 U5844 ( .CLK(n5961), .C(n5962) );
  BUFFD0 U5845 ( .I(n5962), .Z(n5963) );
  CKBD0 U5846 ( .CLK(n5963), .C(n5964) );
  CKBD0 U5847 ( .CLK(n5964), .C(n5965) );
  CKBD0 U5848 ( .CLK(n5965), .C(n5966) );
  CKBD0 U5849 ( .CLK(n5966), .C(n5967) );
  CKBD0 U5850 ( .CLK(n5967), .C(n5968) );
  CKBD0 U5851 ( .CLK(n5968), .C(n5969) );
  CKBD0 U5852 ( .CLK(n5969), .C(n5970) );
  CKBD0 U5853 ( .CLK(n5970), .C(n5971) );
  CKBD0 U5854 ( .CLK(n5971), .C(n5972) );
  CKBD0 U5855 ( .CLK(n5972), .C(n5973) );
  CKBD0 U5856 ( .CLK(n5973), .C(n5974) );
  BUFFD0 U5857 ( .I(n5974), .Z(n5975) );
  CKBD0 U5858 ( .CLK(n5975), .C(n5976) );
  CKBD0 U5859 ( .CLK(n5976), .C(n5977) );
  CKBD0 U5860 ( .CLK(n5977), .C(n5978) );
  CKBD0 U5861 ( .CLK(n5978), .C(n5979) );
  CKBD0 U5862 ( .CLK(n5979), .C(n5980) );
  CKBD0 U5863 ( .CLK(n5980), .C(n5981) );
  CKBD0 U5864 ( .CLK(n5981), .C(n5982) );
  CKBD0 U5865 ( .CLK(n5982), .C(n5983) );
  CKBD0 U5866 ( .CLK(n5983), .C(n5984) );
  BUFFD0 U5867 ( .I(n5984), .Z(n5985) );
  CKBD0 U5868 ( .CLK(n5985), .C(n5986) );
  CKBD0 U5869 ( .CLK(n5986), .C(n5987) );
  CKBD0 U5870 ( .CLK(n5987), .C(n5988) );
  CKBD0 U5871 ( .CLK(n5988), .C(n5989) );
  CKBD0 U5872 ( .CLK(n5989), .C(n5990) );
  CKBD0 U5873 ( .CLK(n5990), .C(n5991) );
  CKBD0 U5874 ( .CLK(n5991), .C(n5992) );
  CKBD0 U5875 ( .CLK(n5992), .C(n5993) );
  CKBD0 U5876 ( .CLK(n5993), .C(n5994) );
  BUFFD0 U5877 ( .I(n5994), .Z(n5995) );
  CKBD0 U5878 ( .CLK(n5995), .C(n5996) );
  CKBD0 U5879 ( .CLK(n5996), .C(n5997) );
  CKBD0 U5880 ( .CLK(n5997), .C(n5998) );
  CKBD0 U5881 ( .CLK(n5998), .C(n5999) );
  CKBD0 U5882 ( .CLK(n5999), .C(n6000) );
  CKBD0 U5883 ( .CLK(n6000), .C(n6001) );
  CKBD0 U5884 ( .CLK(n6001), .C(n6002) );
  CKBD0 U5885 ( .CLK(n6002), .C(n6003) );
  CKBD0 U5886 ( .CLK(n6003), .C(n6004) );
  CKBD0 U5887 ( .CLK(n6004), .C(n6005) );
  CKBD0 U5888 ( .CLK(n6005), .C(n6006) );
  BUFFD0 U5889 ( .I(n6006), .Z(n6007) );
  CKBD0 U5890 ( .CLK(n6007), .C(n6008) );
  CKBD0 U5891 ( .CLK(n6008), .C(n6009) );
  CKBD0 U5892 ( .CLK(n6009), .C(n6010) );
  CKBD0 U5893 ( .CLK(n6010), .C(n6011) );
  CKBD0 U5894 ( .CLK(n6011), .C(n6012) );
  CKBD0 U5895 ( .CLK(n6012), .C(n6013) );
  CKBD0 U5896 ( .CLK(n6013), .C(n6014) );
  CKBD0 U5897 ( .CLK(n6014), .C(n6015) );
  CKBD0 U5898 ( .CLK(n6015), .C(n6016) );
  CKBD0 U5899 ( .CLK(n6016), .C(n6017) );
  BUFFD0 U5900 ( .I(n6017), .Z(n6018) );
  CKBD0 U5901 ( .CLK(n6018), .C(n6019) );
  CKBD0 U5902 ( .CLK(n6019), .C(n6020) );
  CKBD0 U5903 ( .CLK(n6020), .C(n6021) );
  CKBD0 U5904 ( .CLK(n6021), .C(n6022) );
  CKBD0 U5905 ( .CLK(n6022), .C(n6023) );
  BUFFD0 U5906 ( .I(n6023), .Z(n6024) );
  CKBD0 U5907 ( .CLK(n6024), .C(n6025) );
  BUFFD0 U5908 ( .I(n6025), .Z(n6026) );
  CKBD0 U5909 ( .CLK(n6026), .C(n6027) );
  BUFFD0 U5910 ( .I(n6027), .Z(n6028) );
  CKBD0 U5911 ( .CLK(n6028), .C(n6029) );
  BUFFD0 U5912 ( .I(n6029), .Z(n6030) );
  CKBD0 U5913 ( .CLK(n6030), .C(n6031) );
  BUFFD0 U5914 ( .I(n6031), .Z(n6032) );
  CKBD0 U5915 ( .CLK(n6032), .C(n6033) );
  BUFFD0 U5916 ( .I(n6033), .Z(n6034) );
  CKBD0 U5917 ( .CLK(n6034), .C(n6035) );
  BUFFD0 U5918 ( .I(n6035), .Z(n6036) );
  CKBD0 U5919 ( .CLK(n6036), .C(n6037) );
  BUFFD0 U5920 ( .I(n6037), .Z(n6038) );
  BUFFD0 U5921 ( .I(n137), .Z(n6039) );
  BUFFD0 U5922 ( .I(n6041), .Z(n6040) );
  BUFFD0 U5923 ( .I(n6042), .Z(n6041) );
  BUFFD0 U5924 ( .I(Decoder[4]), .Z(n6042) );
  CKBD0 U5925 ( .CLK(n866), .C(n6043) );
  CKBD0 U5926 ( .CLK(n6043), .C(n6044) );
  CKBD0 U5927 ( .CLK(n6044), .C(n6045) );
  BUFFD0 U5928 ( .I(n6045), .Z(n6046) );
  CKBD0 U5929 ( .CLK(n6046), .C(n6047) );
  CKBD0 U5930 ( .CLK(n6047), .C(n6048) );
  CKBD0 U5931 ( .CLK(n6048), .C(n6049) );
  CKBD0 U5932 ( .CLK(n6049), .C(n6050) );
  CKBD0 U5933 ( .CLK(n6050), .C(n6051) );
  CKBD0 U5934 ( .CLK(n6051), .C(n6052) );
  CKBD0 U5935 ( .CLK(n6052), .C(n6053) );
  CKBD0 U5936 ( .CLK(n6053), .C(n6054) );
  CKBD0 U5937 ( .CLK(n6054), .C(n6055) );
  CKBD0 U5938 ( .CLK(n6055), .C(n6056) );
  BUFFD0 U5939 ( .I(n6056), .Z(n6057) );
  CKBD0 U5940 ( .CLK(n6057), .C(n6058) );
  CKBD0 U5941 ( .CLK(n6058), .C(n6059) );
  CKBD0 U5942 ( .CLK(n6059), .C(n6060) );
  CKBD0 U5943 ( .CLK(n6060), .C(n6061) );
  CKBD0 U5944 ( .CLK(n6061), .C(n6062) );
  CKBD0 U5945 ( .CLK(n6062), .C(n6063) );
  CKBD0 U5946 ( .CLK(n6063), .C(n6064) );
  CKBD0 U5947 ( .CLK(n6064), .C(n6065) );
  CKBD0 U5948 ( .CLK(n6065), .C(n6066) );
  CKBD0 U5949 ( .CLK(n6066), .C(n6067) );
  BUFFD0 U5950 ( .I(n6067), .Z(n6068) );
  CKBD0 U5951 ( .CLK(n6068), .C(n6069) );
  CKBD0 U5952 ( .CLK(n6069), .C(n6070) );
  CKBD0 U5953 ( .CLK(n6070), .C(n6071) );
  CKBD0 U5954 ( .CLK(n6071), .C(n6072) );
  CKBD0 U5955 ( .CLK(n6072), .C(n6073) );
  CKBD0 U5956 ( .CLK(n6073), .C(n6074) );
  CKBD0 U5957 ( .CLK(n6074), .C(n6075) );
  CKBD0 U5958 ( .CLK(n6075), .C(n6076) );
  CKBD0 U5959 ( .CLK(n6076), .C(n6077) );
  BUFFD0 U5960 ( .I(n6077), .Z(n6078) );
  CKBD0 U5961 ( .CLK(n6078), .C(n6079) );
  CKBD0 U5962 ( .CLK(n6079), .C(n6080) );
  CKBD0 U5963 ( .CLK(n6080), .C(n6081) );
  CKBD0 U5964 ( .CLK(n6081), .C(n6082) );
  CKBD0 U5965 ( .CLK(n6082), .C(n6083) );
  CKBD0 U5966 ( .CLK(n6083), .C(n6084) );
  CKBD0 U5967 ( .CLK(n6084), .C(n6085) );
  CKBD0 U5968 ( .CLK(n6085), .C(n6086) );
  CKBD0 U5969 ( .CLK(n6086), .C(n6087) );
  CKBD0 U5970 ( .CLK(n6087), .C(n6088) );
  CKBD0 U5971 ( .CLK(n6088), .C(n6089) );
  BUFFD0 U5972 ( .I(n6089), .Z(n6090) );
  CKBD0 U5973 ( .CLK(n6090), .C(n6091) );
  CKBD0 U5974 ( .CLK(n6091), .C(n6092) );
  CKBD0 U5975 ( .CLK(n6092), .C(n6093) );
  CKBD0 U5976 ( .CLK(n6093), .C(n6094) );
  CKBD0 U5977 ( .CLK(n6094), .C(n6095) );
  CKBD0 U5978 ( .CLK(n6095), .C(n6096) );
  CKBD0 U5979 ( .CLK(n6096), .C(n6097) );
  CKBD0 U5980 ( .CLK(n6097), .C(n6098) );
  CKBD0 U5981 ( .CLK(n6098), .C(n6099) );
  CKBD0 U5982 ( .CLK(n6099), .C(n6100) );
  BUFFD0 U5983 ( .I(n6100), .Z(n6101) );
  CKBD0 U5984 ( .CLK(n6101), .C(n6102) );
  CKBD0 U5985 ( .CLK(n6102), .C(n6103) );
  CKBD0 U5986 ( .CLK(n6103), .C(n6104) );
  CKBD0 U5987 ( .CLK(n6104), .C(n6105) );
  CKBD0 U5988 ( .CLK(n6105), .C(n6106) );
  CKBD0 U5989 ( .CLK(n6106), .C(n6107) );
  CKBD0 U5990 ( .CLK(n6107), .C(n6108) );
  CKBD0 U5991 ( .CLK(n6108), .C(n6109) );
  CKBD0 U5992 ( .CLK(n6109), .C(n6110) );
  BUFFD0 U5993 ( .I(n6110), .Z(n6111) );
  CKBD0 U5994 ( .CLK(n6111), .C(n6112) );
  CKBD0 U5995 ( .CLK(n6112), .C(n6113) );
  CKBD0 U5996 ( .CLK(n6113), .C(n6114) );
  CKBD0 U5997 ( .CLK(n6114), .C(n6115) );
  CKBD0 U5998 ( .CLK(n6115), .C(n6116) );
  CKBD0 U5999 ( .CLK(n6116), .C(n6117) );
  CKBD0 U6000 ( .CLK(n6117), .C(n6118) );
  CKBD0 U6001 ( .CLK(n6118), .C(n6119) );
  CKBD0 U6002 ( .CLK(n6119), .C(n6120) );
  CKBD0 U6003 ( .CLK(n6120), .C(n6121) );
  CKBD0 U6004 ( .CLK(n6121), .C(n6122) );
  BUFFD0 U6005 ( .I(n6122), .Z(n6123) );
  CKBD0 U6006 ( .CLK(n6123), .C(n6124) );
  CKBD0 U6007 ( .CLK(n6124), .C(n6125) );
  CKBD0 U6008 ( .CLK(n6125), .C(n6126) );
  CKBD0 U6009 ( .CLK(n6126), .C(n6127) );
  CKBD0 U6010 ( .CLK(n6127), .C(n6128) );
  CKBD0 U6011 ( .CLK(n6128), .C(n6129) );
  CKBD0 U6012 ( .CLK(n6129), .C(n6130) );
  CKBD0 U6013 ( .CLK(n6130), .C(n6131) );
  CKBD0 U6014 ( .CLK(n6131), .C(n6132) );
  BUFFD0 U6015 ( .I(n6132), .Z(n6133) );
  CKBD0 U6016 ( .CLK(n6133), .C(n6134) );
  CKBD0 U6017 ( .CLK(n6134), .C(n6135) );
  CKBD0 U6018 ( .CLK(n6135), .C(n6136) );
  CKBD0 U6019 ( .CLK(n6136), .C(n6137) );
  CKBD0 U6020 ( .CLK(n6137), .C(n6138) );
  CKBD0 U6021 ( .CLK(n6138), .C(n6139) );
  CKBD0 U6022 ( .CLK(n6139), .C(n6140) );
  CKBD0 U6023 ( .CLK(n6140), .C(n6141) );
  CKBD0 U6024 ( .CLK(n6141), .C(n6142) );
  BUFFD0 U6025 ( .I(n6142), .Z(n6143) );
  CKBD0 U6026 ( .CLK(n6143), .C(n6144) );
  CKBD0 U6027 ( .CLK(n6144), .C(n6145) );
  CKBD0 U6028 ( .CLK(n6145), .C(n6146) );
  CKBD0 U6029 ( .CLK(n6146), .C(n6147) );
  CKBD0 U6030 ( .CLK(n6147), .C(n6148) );
  CKBD0 U6031 ( .CLK(n6148), .C(n6149) );
  CKBD0 U6032 ( .CLK(n6149), .C(n6150) );
  CKBD0 U6033 ( .CLK(n6150), .C(n6151) );
  CKBD0 U6034 ( .CLK(n6151), .C(n6152) );
  CKBD0 U6035 ( .CLK(n6152), .C(n6153) );
  CKBD0 U6036 ( .CLK(n6153), .C(n6154) );
  BUFFD0 U6037 ( .I(n6154), .Z(n6155) );
  CKBD0 U6038 ( .CLK(n6155), .C(n6156) );
  CKBD0 U6039 ( .CLK(n6156), .C(n6157) );
  CKBD0 U6040 ( .CLK(n6157), .C(n6158) );
  CKBD0 U6041 ( .CLK(n6158), .C(n6159) );
  CKBD0 U6042 ( .CLK(n6159), .C(n6160) );
  BUFFD0 U6043 ( .I(n6160), .Z(n6161) );
  CKBD0 U6044 ( .CLK(n6161), .C(n6162) );
  BUFFD0 U6045 ( .I(n6162), .Z(n6163) );
  CKBD0 U6046 ( .CLK(n6163), .C(n6164) );
  BUFFD0 U6047 ( .I(n6164), .Z(n6165) );
  CKBD0 U6048 ( .CLK(n6165), .C(n6166) );
  BUFFD0 U6049 ( .I(n6166), .Z(n6167) );
  CKBD0 U6050 ( .CLK(n6167), .C(n6168) );
  BUFFD0 U6051 ( .I(n6168), .Z(n6169) );
  CKBD0 U6052 ( .CLK(n6169), .C(n6170) );
  BUFFD0 U6053 ( .I(n6170), .Z(n6171) );
  CKBD0 U6054 ( .CLK(n6171), .C(n6172) );
  BUFFD0 U6055 ( .I(n6172), .Z(n6173) );
  CKBD0 U6056 ( .CLK(n6173), .C(n6174) );
  BUFFD0 U6057 ( .I(n6174), .Z(n6175) );
  BUFFD0 U6058 ( .I(n136), .Z(n6176) );
  BUFFD0 U6059 ( .I(n6178), .Z(n6177) );
  BUFFD0 U6060 ( .I(n6179), .Z(n6178) );
  BUFFD0 U6061 ( .I(Decoder[3]), .Z(n6179) );
  CKBD0 U6062 ( .CLK(n864), .C(n6180) );
  CKBD0 U6063 ( .CLK(n6180), .C(n6181) );
  CKBD0 U6064 ( .CLK(n6181), .C(n6182) );
  BUFFD0 U6065 ( .I(n6182), .Z(n6183) );
  CKBD0 U6066 ( .CLK(n6183), .C(n6184) );
  CKBD0 U6067 ( .CLK(n6184), .C(n6185) );
  CKBD0 U6068 ( .CLK(n6185), .C(n6186) );
  CKBD0 U6069 ( .CLK(n6186), .C(n6187) );
  CKBD0 U6070 ( .CLK(n6187), .C(n6188) );
  CKBD0 U6071 ( .CLK(n6188), .C(n6189) );
  CKBD0 U6072 ( .CLK(n6189), .C(n6190) );
  CKBD0 U6073 ( .CLK(n6190), .C(n6191) );
  CKBD0 U6074 ( .CLK(n6191), .C(n6192) );
  CKBD0 U6075 ( .CLK(n6192), .C(n6193) );
  BUFFD0 U6076 ( .I(n6193), .Z(n6194) );
  CKBD0 U6077 ( .CLK(n6194), .C(n6195) );
  CKBD0 U6078 ( .CLK(n6195), .C(n6196) );
  CKBD0 U6079 ( .CLK(n6196), .C(n6197) );
  CKBD0 U6080 ( .CLK(n6197), .C(n6198) );
  CKBD0 U6081 ( .CLK(n6198), .C(n6199) );
  CKBD0 U6082 ( .CLK(n6199), .C(n6200) );
  CKBD0 U6083 ( .CLK(n6200), .C(n6201) );
  CKBD0 U6084 ( .CLK(n6201), .C(n6202) );
  CKBD0 U6085 ( .CLK(n6202), .C(n6203) );
  CKBD0 U6086 ( .CLK(n6203), .C(n6204) );
  BUFFD0 U6087 ( .I(n6204), .Z(n6205) );
  CKBD0 U6088 ( .CLK(n6205), .C(n6206) );
  CKBD0 U6089 ( .CLK(n6206), .C(n6207) );
  CKBD0 U6090 ( .CLK(n6207), .C(n6208) );
  CKBD0 U6091 ( .CLK(n6208), .C(n6209) );
  CKBD0 U6092 ( .CLK(n6209), .C(n6210) );
  CKBD0 U6093 ( .CLK(n6210), .C(n6211) );
  CKBD0 U6094 ( .CLK(n6211), .C(n6212) );
  CKBD0 U6095 ( .CLK(n6212), .C(n6213) );
  CKBD0 U6096 ( .CLK(n6213), .C(n6214) );
  CKBD0 U6097 ( .CLK(n6214), .C(n6215) );
  BUFFD0 U6098 ( .I(n6215), .Z(n6216) );
  CKBD0 U6099 ( .CLK(n6216), .C(n6217) );
  CKBD0 U6100 ( .CLK(n6217), .C(n6218) );
  CKBD0 U6101 ( .CLK(n6218), .C(n6219) );
  CKBD0 U6102 ( .CLK(n6219), .C(n6220) );
  CKBD0 U6103 ( .CLK(n6220), .C(n6221) );
  CKBD0 U6104 ( .CLK(n6221), .C(n6222) );
  CKBD0 U6105 ( .CLK(n6222), .C(n6223) );
  CKBD0 U6106 ( .CLK(n6223), .C(n6224) );
  CKBD0 U6107 ( .CLK(n6224), .C(n6225) );
  BUFFD0 U6108 ( .I(n6225), .Z(n6226) );
  CKBD0 U6109 ( .CLK(n6226), .C(n6227) );
  CKBD0 U6110 ( .CLK(n6227), .C(n6228) );
  CKBD0 U6111 ( .CLK(n6228), .C(n6229) );
  CKBD0 U6112 ( .CLK(n6229), .C(n6230) );
  CKBD0 U6113 ( .CLK(n6230), .C(n6231) );
  CKBD0 U6114 ( .CLK(n6231), .C(n6232) );
  CKBD0 U6115 ( .CLK(n6232), .C(n6233) );
  CKBD0 U6116 ( .CLK(n6233), .C(n6234) );
  CKBD0 U6117 ( .CLK(n6234), .C(n6235) );
  CKBD0 U6118 ( .CLK(n6235), .C(n6236) );
  CKBD0 U6119 ( .CLK(n6236), .C(n6237) );
  BUFFD0 U6120 ( .I(n6237), .Z(n6238) );
  CKBD0 U6121 ( .CLK(n6238), .C(n6239) );
  CKBD0 U6122 ( .CLK(n6239), .C(n6240) );
  CKBD0 U6123 ( .CLK(n6240), .C(n6241) );
  CKBD0 U6124 ( .CLK(n6241), .C(n6242) );
  CKBD0 U6125 ( .CLK(n6242), .C(n6243) );
  CKBD0 U6126 ( .CLK(n6243), .C(n6244) );
  CKBD0 U6127 ( .CLK(n6244), .C(n6245) );
  CKBD0 U6128 ( .CLK(n6245), .C(n6246) );
  CKBD0 U6129 ( .CLK(n6246), .C(n6247) );
  BUFFD0 U6130 ( .I(n6247), .Z(n6248) );
  CKBD0 U6131 ( .CLK(n6248), .C(n6249) );
  CKBD0 U6132 ( .CLK(n6249), .C(n6250) );
  CKBD0 U6133 ( .CLK(n6250), .C(n6251) );
  CKBD0 U6134 ( .CLK(n6251), .C(n6252) );
  CKBD0 U6135 ( .CLK(n6252), .C(n6253) );
  CKBD0 U6136 ( .CLK(n6253), .C(n6254) );
  CKBD0 U6137 ( .CLK(n6254), .C(n6255) );
  CKBD0 U6138 ( .CLK(n6255), .C(n6256) );
  CKBD0 U6139 ( .CLK(n6256), .C(n6257) );
  CKBD0 U6140 ( .CLK(n6257), .C(n6258) );
  BUFFD0 U6141 ( .I(n6258), .Z(n6259) );
  CKBD0 U6142 ( .CLK(n6259), .C(n6260) );
  CKBD0 U6143 ( .CLK(n6260), .C(n6261) );
  CKBD0 U6144 ( .CLK(n6261), .C(n6262) );
  CKBD0 U6145 ( .CLK(n6262), .C(n6263) );
  CKBD0 U6146 ( .CLK(n6263), .C(n6264) );
  CKBD0 U6147 ( .CLK(n6264), .C(n6265) );
  CKBD0 U6148 ( .CLK(n6265), .C(n6266) );
  CKBD0 U6149 ( .CLK(n6266), .C(n6267) );
  CKBD0 U6150 ( .CLK(n6267), .C(n6268) );
  CKBD0 U6151 ( .CLK(n6268), .C(n6269) );
  CKBD0 U6152 ( .CLK(n6269), .C(n6270) );
  BUFFD0 U6153 ( .I(n6270), .Z(n6271) );
  CKBD0 U6154 ( .CLK(n6271), .C(n6272) );
  CKBD0 U6155 ( .CLK(n6272), .C(n6273) );
  CKBD0 U6156 ( .CLK(n6273), .C(n6274) );
  CKBD0 U6157 ( .CLK(n6274), .C(n6275) );
  CKBD0 U6158 ( .CLK(n6275), .C(n6276) );
  CKBD0 U6159 ( .CLK(n6276), .C(n6277) );
  CKBD0 U6160 ( .CLK(n6277), .C(n6278) );
  CKBD0 U6161 ( .CLK(n6278), .C(n6279) );
  CKBD0 U6162 ( .CLK(n6279), .C(n6280) );
  BUFFD0 U6163 ( .I(n6280), .Z(n6281) );
  CKBD0 U6164 ( .CLK(n6281), .C(n6282) );
  CKBD0 U6165 ( .CLK(n6282), .C(n6283) );
  CKBD0 U6166 ( .CLK(n6283), .C(n6284) );
  CKBD0 U6167 ( .CLK(n6284), .C(n6285) );
  CKBD0 U6168 ( .CLK(n6285), .C(n6286) );
  CKBD0 U6169 ( .CLK(n6286), .C(n6287) );
  CKBD0 U6170 ( .CLK(n6287), .C(n6288) );
  CKBD0 U6171 ( .CLK(n6288), .C(n6289) );
  CKBD0 U6172 ( .CLK(n6289), .C(n6290) );
  BUFFD0 U6173 ( .I(n6290), .Z(n6291) );
  CKBD0 U6174 ( .CLK(n6291), .C(n6292) );
  CKBD0 U6175 ( .CLK(n6292), .C(n6293) );
  CKBD0 U6176 ( .CLK(n6293), .C(n6294) );
  CKBD0 U6177 ( .CLK(n6294), .C(n6295) );
  CKBD0 U6178 ( .CLK(n6295), .C(n6296) );
  CKBD0 U6179 ( .CLK(n6296), .C(n6297) );
  BUFFD0 U6180 ( .I(n6297), .Z(n6298) );
  CKBD0 U6181 ( .CLK(n6298), .C(n6299) );
  BUFFD0 U6182 ( .I(n6299), .Z(n6300) );
  CKBD0 U6183 ( .CLK(n6300), .C(n6301) );
  BUFFD0 U6184 ( .I(n6301), .Z(n6302) );
  CKBD0 U6185 ( .CLK(n6302), .C(n6303) );
  BUFFD0 U6186 ( .I(n6303), .Z(n6304) );
  CKBD0 U6187 ( .CLK(n6304), .C(n6305) );
  BUFFD0 U6188 ( .I(n6305), .Z(n6306) );
  CKBD0 U6189 ( .CLK(n6306), .C(n6307) );
  BUFFD0 U6190 ( .I(n6307), .Z(n6308) );
  CKBD0 U6191 ( .CLK(n6308), .C(n6309) );
  BUFFD0 U6192 ( .I(n6309), .Z(n6310) );
  CKBD0 U6193 ( .CLK(n6310), .C(n6311) );
  BUFFD0 U6194 ( .I(n6311), .Z(n6312) );
  BUFFD0 U6195 ( .I(n135), .Z(n6313) );
  BUFFD0 U6196 ( .I(n6315), .Z(n6314) );
  BUFFD0 U6197 ( .I(n6316), .Z(n6315) );
  BUFFD0 U6198 ( .I(Decoder[2]), .Z(n6316) );
  CKBD0 U6199 ( .CLK(n862), .C(n6317) );
  CKBD0 U6200 ( .CLK(n6317), .C(n6318) );
  CKBD0 U6201 ( .CLK(n6318), .C(n6319) );
  BUFFD0 U6202 ( .I(n6319), .Z(n6320) );
  CKBD0 U6203 ( .CLK(n6320), .C(n6321) );
  CKBD0 U6204 ( .CLK(n6321), .C(n6322) );
  CKBD0 U6205 ( .CLK(n6322), .C(n6323) );
  CKBD0 U6206 ( .CLK(n6323), .C(n6324) );
  CKBD0 U6207 ( .CLK(n6324), .C(n6325) );
  CKBD0 U6208 ( .CLK(n6325), .C(n6326) );
  CKBD0 U6209 ( .CLK(n6326), .C(n6327) );
  CKBD0 U6210 ( .CLK(n6327), .C(n6328) );
  CKBD0 U6211 ( .CLK(n6328), .C(n6329) );
  CKBD0 U6212 ( .CLK(n6329), .C(n6330) );
  BUFFD0 U6213 ( .I(n6330), .Z(n6331) );
  CKBD0 U6214 ( .CLK(n6331), .C(n6332) );
  CKBD0 U6215 ( .CLK(n6332), .C(n6333) );
  CKBD0 U6216 ( .CLK(n6333), .C(n6334) );
  CKBD0 U6217 ( .CLK(n6334), .C(n6335) );
  CKBD0 U6218 ( .CLK(n6335), .C(n6336) );
  CKBD0 U6219 ( .CLK(n6336), .C(n6337) );
  CKBD0 U6220 ( .CLK(n6337), .C(n6338) );
  CKBD0 U6221 ( .CLK(n6338), .C(n6339) );
  CKBD0 U6222 ( .CLK(n6339), .C(n6340) );
  CKBD0 U6223 ( .CLK(n6340), .C(n6341) );
  BUFFD0 U6224 ( .I(n6341), .Z(n6342) );
  CKBD0 U6225 ( .CLK(n6342), .C(n6343) );
  CKBD0 U6226 ( .CLK(n6343), .C(n6344) );
  CKBD0 U6227 ( .CLK(n6344), .C(n6345) );
  CKBD0 U6228 ( .CLK(n6345), .C(n6346) );
  CKBD0 U6229 ( .CLK(n6346), .C(n6347) );
  CKBD0 U6230 ( .CLK(n6347), .C(n6348) );
  CKBD0 U6231 ( .CLK(n6348), .C(n6349) );
  CKBD0 U6232 ( .CLK(n6349), .C(n6350) );
  CKBD0 U6233 ( .CLK(n6350), .C(n6351) );
  BUFFD0 U6234 ( .I(n6351), .Z(n6352) );
  CKBD0 U6235 ( .CLK(n6352), .C(n6353) );
  CKBD0 U6236 ( .CLK(n6353), .C(n6354) );
  CKBD0 U6237 ( .CLK(n6354), .C(n6355) );
  CKBD0 U6238 ( .CLK(n6355), .C(n6356) );
  CKBD0 U6239 ( .CLK(n6356), .C(n6357) );
  CKBD0 U6240 ( .CLK(n6357), .C(n6358) );
  CKBD0 U6241 ( .CLK(n6358), .C(n6359) );
  CKBD0 U6242 ( .CLK(n6359), .C(n6360) );
  CKBD0 U6243 ( .CLK(n6360), .C(n6361) );
  CKBD0 U6244 ( .CLK(n6361), .C(n6362) );
  CKBD0 U6245 ( .CLK(n6362), .C(n6363) );
  BUFFD0 U6246 ( .I(n6363), .Z(n6364) );
  CKBD0 U6247 ( .CLK(n6364), .C(n6365) );
  CKBD0 U6248 ( .CLK(n6365), .C(n6366) );
  CKBD0 U6249 ( .CLK(n6366), .C(n6367) );
  CKBD0 U6250 ( .CLK(n6367), .C(n6368) );
  CKBD0 U6251 ( .CLK(n6368), .C(n6369) );
  CKBD0 U6252 ( .CLK(n6369), .C(n6370) );
  CKBD0 U6253 ( .CLK(n6370), .C(n6371) );
  CKBD0 U6254 ( .CLK(n6371), .C(n6372) );
  CKBD0 U6255 ( .CLK(n6372), .C(n6373) );
  BUFFD0 U6256 ( .I(n6373), .Z(n6374) );
  CKBD0 U6257 ( .CLK(n6374), .C(n6375) );
  CKBD0 U6258 ( .CLK(n6375), .C(n6376) );
  CKBD0 U6259 ( .CLK(n6376), .C(n6377) );
  CKBD0 U6260 ( .CLK(n6377), .C(n6378) );
  CKBD0 U6261 ( .CLK(n6378), .C(n6379) );
  CKBD0 U6262 ( .CLK(n6379), .C(n6380) );
  CKBD0 U6263 ( .CLK(n6380), .C(n6381) );
  CKBD0 U6264 ( .CLK(n6381), .C(n6382) );
  CKBD0 U6265 ( .CLK(n6382), .C(n6383) );
  CKBD0 U6266 ( .CLK(n6383), .C(n6384) );
  BUFFD0 U6267 ( .I(n6384), .Z(n6385) );
  CKBD0 U6268 ( .CLK(n6385), .C(n6386) );
  CKBD0 U6269 ( .CLK(n6386), .C(n6387) );
  CKBD0 U6270 ( .CLK(n6387), .C(n6388) );
  CKBD0 U6271 ( .CLK(n6388), .C(n6389) );
  CKBD0 U6272 ( .CLK(n6389), .C(n6390) );
  CKBD0 U6273 ( .CLK(n6390), .C(n6391) );
  CKBD0 U6274 ( .CLK(n6391), .C(n6392) );
  CKBD0 U6275 ( .CLK(n6392), .C(n6393) );
  CKBD0 U6276 ( .CLK(n6393), .C(n6394) );
  CKBD0 U6277 ( .CLK(n6394), .C(n6395) );
  BUFFD0 U6278 ( .I(n6395), .Z(n6396) );
  CKBD0 U6279 ( .CLK(n6396), .C(n6397) );
  CKBD0 U6280 ( .CLK(n6397), .C(n6398) );
  CKBD0 U6281 ( .CLK(n6398), .C(n6399) );
  CKBD0 U6282 ( .CLK(n6399), .C(n6400) );
  CKBD0 U6283 ( .CLK(n6400), .C(n6401) );
  CKBD0 U6284 ( .CLK(n6401), .C(n6402) );
  CKBD0 U6285 ( .CLK(n6402), .C(n6403) );
  CKBD0 U6286 ( .CLK(n6403), .C(n6404) );
  CKBD0 U6287 ( .CLK(n6404), .C(n6405) );
  CKBD0 U6288 ( .CLK(n6405), .C(n6406) );
  BUFFD0 U6289 ( .I(n6406), .Z(n6407) );
  CKBD0 U6290 ( .CLK(n6407), .C(n6408) );
  CKBD0 U6291 ( .CLK(n6408), .C(n6409) );
  CKBD0 U6292 ( .CLK(n6409), .C(n6410) );
  CKBD0 U6293 ( .CLK(n6410), .C(n6411) );
  CKBD0 U6294 ( .CLK(n6411), .C(n6412) );
  CKBD0 U6295 ( .CLK(n6412), .C(n6413) );
  CKBD0 U6296 ( .CLK(n6413), .C(n6414) );
  CKBD0 U6297 ( .CLK(n6414), .C(n6415) );
  CKBD0 U6298 ( .CLK(n6415), .C(n6416) );
  CKBD0 U6299 ( .CLK(n6416), .C(n6417) );
  BUFFD0 U6300 ( .I(n6417), .Z(n6418) );
  CKBD0 U6301 ( .CLK(n6418), .C(n6419) );
  CKBD0 U6302 ( .CLK(n6419), .C(n6420) );
  CKBD0 U6303 ( .CLK(n6420), .C(n6421) );
  CKBD0 U6304 ( .CLK(n6421), .C(n6422) );
  CKBD0 U6305 ( .CLK(n6422), .C(n6423) );
  CKBD0 U6306 ( .CLK(n6423), .C(n6424) );
  CKBD0 U6307 ( .CLK(n6424), .C(n6425) );
  CKBD0 U6308 ( .CLK(n6425), .C(n6426) );
  CKBD0 U6309 ( .CLK(n6426), .C(n6427) );
  CKBD0 U6310 ( .CLK(n6427), .C(n6428) );
  BUFFD0 U6311 ( .I(n6428), .Z(n6429) );
  CKBD0 U6312 ( .CLK(n6429), .C(n6430) );
  CKBD0 U6313 ( .CLK(n6430), .C(n6431) );
  CKBD0 U6314 ( .CLK(n6431), .C(n6432) );
  CKBD0 U6315 ( .CLK(n6432), .C(n6433) );
  CKBD0 U6316 ( .CLK(n6433), .C(n6434) );
  BUFFD0 U6317 ( .I(n6434), .Z(n6435) );
  CKBD0 U6318 ( .CLK(n6435), .C(n6436) );
  BUFFD0 U6319 ( .I(n6436), .Z(n6437) );
  CKBD0 U6320 ( .CLK(n6437), .C(n6438) );
  BUFFD0 U6321 ( .I(n6438), .Z(n6439) );
  CKBD0 U6322 ( .CLK(n6439), .C(n6440) );
  BUFFD0 U6323 ( .I(n6440), .Z(n6441) );
  CKBD0 U6324 ( .CLK(n6441), .C(n6442) );
  BUFFD0 U6325 ( .I(n6442), .Z(n6443) );
  CKBD0 U6326 ( .CLK(n6443), .C(n6444) );
  BUFFD0 U6327 ( .I(n6444), .Z(n6445) );
  CKBD0 U6328 ( .CLK(n6445), .C(n6446) );
  BUFFD0 U6329 ( .I(n6446), .Z(n6447) );
  CKBD0 U6330 ( .CLK(n6447), .C(n6448) );
  BUFFD0 U6331 ( .I(n6448), .Z(n6449) );
  BUFFD0 U6332 ( .I(n134), .Z(n6450) );
  BUFFD0 U6333 ( .I(n6452), .Z(n6451) );
  BUFFD0 U6334 ( .I(n6453), .Z(n6452) );
  BUFFD0 U6335 ( .I(Decoder[1]), .Z(n6453) );
  CKBD0 U6336 ( .CLK(n860), .C(n6454) );
  CKBD0 U6337 ( .CLK(n6454), .C(n6455) );
  CKBD0 U6338 ( .CLK(n6455), .C(n6456) );
  BUFFD0 U6339 ( .I(n6456), .Z(n6457) );
  CKBD0 U6340 ( .CLK(n6457), .C(n6458) );
  CKBD0 U6341 ( .CLK(n6458), .C(n6459) );
  CKBD0 U6342 ( .CLK(n6459), .C(n6460) );
  CKBD0 U6343 ( .CLK(n6460), .C(n6461) );
  CKBD0 U6344 ( .CLK(n6461), .C(n6462) );
  CKBD0 U6345 ( .CLK(n6462), .C(n6463) );
  CKBD0 U6346 ( .CLK(n6463), .C(n6464) );
  CKBD0 U6347 ( .CLK(n6464), .C(n6465) );
  CKBD0 U6348 ( .CLK(n6465), .C(n6466) );
  CKBD0 U6349 ( .CLK(n6466), .C(n6467) );
  BUFFD0 U6350 ( .I(n6467), .Z(n6468) );
  CKBD0 U6351 ( .CLK(n6468), .C(n6469) );
  CKBD0 U6352 ( .CLK(n6469), .C(n6470) );
  CKBD0 U6353 ( .CLK(n6470), .C(n6471) );
  CKBD0 U6354 ( .CLK(n6471), .C(n6472) );
  CKBD0 U6355 ( .CLK(n6472), .C(n6473) );
  CKBD0 U6356 ( .CLK(n6473), .C(n6474) );
  CKBD0 U6357 ( .CLK(n6474), .C(n6475) );
  CKBD0 U6358 ( .CLK(n6475), .C(n6476) );
  CKBD0 U6359 ( .CLK(n6476), .C(n6477) );
  CKBD0 U6360 ( .CLK(n6477), .C(n6478) );
  BUFFD0 U6361 ( .I(n6478), .Z(n6479) );
  CKBD0 U6362 ( .CLK(n6479), .C(n6480) );
  CKBD0 U6363 ( .CLK(n6480), .C(n6481) );
  CKBD0 U6364 ( .CLK(n6481), .C(n6482) );
  CKBD0 U6365 ( .CLK(n6482), .C(n6483) );
  CKBD0 U6366 ( .CLK(n6483), .C(n6484) );
  CKBD0 U6367 ( .CLK(n6484), .C(n6485) );
  CKBD0 U6368 ( .CLK(n6485), .C(n6486) );
  CKBD0 U6369 ( .CLK(n6486), .C(n6487) );
  CKBD0 U6370 ( .CLK(n6487), .C(n6488) );
  CKBD0 U6371 ( .CLK(n6488), .C(n6489) );
  BUFFD0 U6372 ( .I(n6489), .Z(n6490) );
  CKBD0 U6373 ( .CLK(n6490), .C(n6491) );
  CKBD0 U6374 ( .CLK(n6491), .C(n6492) );
  CKBD0 U6375 ( .CLK(n6492), .C(n6493) );
  CKBD0 U6376 ( .CLK(n6493), .C(n6494) );
  CKBD0 U6377 ( .CLK(n6494), .C(n6495) );
  CKBD0 U6378 ( .CLK(n6495), .C(n6496) );
  CKBD0 U6379 ( .CLK(n6496), .C(n6497) );
  CKBD0 U6380 ( .CLK(n6497), .C(n6498) );
  CKBD0 U6381 ( .CLK(n6498), .C(n6499) );
  BUFFD0 U6382 ( .I(n6499), .Z(n6500) );
  CKBD0 U6383 ( .CLK(n6500), .C(n6501) );
  CKBD0 U6384 ( .CLK(n6501), .C(n6502) );
  CKBD0 U6385 ( .CLK(n6502), .C(n6503) );
  CKBD0 U6386 ( .CLK(n6503), .C(n6504) );
  CKBD0 U6387 ( .CLK(n6504), .C(n6505) );
  CKBD0 U6388 ( .CLK(n6505), .C(n6506) );
  CKBD0 U6389 ( .CLK(n6506), .C(n6507) );
  CKBD0 U6390 ( .CLK(n6507), .C(n6508) );
  CKBD0 U6391 ( .CLK(n6508), .C(n6509) );
  CKBD0 U6392 ( .CLK(n6509), .C(n6510) );
  CKBD0 U6393 ( .CLK(n6510), .C(n6511) );
  BUFFD0 U6394 ( .I(n6511), .Z(n6512) );
  CKBD0 U6395 ( .CLK(n6512), .C(n6513) );
  CKBD0 U6396 ( .CLK(n6513), .C(n6514) );
  CKBD0 U6397 ( .CLK(n6514), .C(n6515) );
  CKBD0 U6398 ( .CLK(n6515), .C(n6516) );
  CKBD0 U6399 ( .CLK(n6516), .C(n6517) );
  CKBD0 U6400 ( .CLK(n6517), .C(n6518) );
  CKBD0 U6401 ( .CLK(n6518), .C(n6519) );
  CKBD0 U6402 ( .CLK(n6519), .C(n6520) );
  CKBD0 U6403 ( .CLK(n6520), .C(n6521) );
  BUFFD0 U6404 ( .I(n6521), .Z(n6522) );
  CKBD0 U6405 ( .CLK(n6522), .C(n6523) );
  CKBD0 U6406 ( .CLK(n6523), .C(n6524) );
  CKBD0 U6407 ( .CLK(n6524), .C(n6525) );
  CKBD0 U6408 ( .CLK(n6525), .C(n6526) );
  CKBD0 U6409 ( .CLK(n6526), .C(n6527) );
  CKBD0 U6410 ( .CLK(n6527), .C(n6528) );
  CKBD0 U6411 ( .CLK(n6528), .C(n6529) );
  CKBD0 U6412 ( .CLK(n6529), .C(n6530) );
  CKBD0 U6413 ( .CLK(n6530), .C(n6531) );
  CKBD0 U6414 ( .CLK(n6531), .C(n6532) );
  BUFFD0 U6415 ( .I(n6532), .Z(n6533) );
  CKBD0 U6416 ( .CLK(n6533), .C(n6534) );
  CKBD0 U6417 ( .CLK(n6534), .C(n6535) );
  CKBD0 U6418 ( .CLK(n6535), .C(n6536) );
  CKBD0 U6419 ( .CLK(n6536), .C(n6537) );
  CKBD0 U6420 ( .CLK(n6537), .C(n6538) );
  CKBD0 U6421 ( .CLK(n6538), .C(n6539) );
  CKBD0 U6422 ( .CLK(n6539), .C(n6540) );
  CKBD0 U6423 ( .CLK(n6540), .C(n6541) );
  CKBD0 U6424 ( .CLK(n6541), .C(n6542) );
  CKBD0 U6425 ( .CLK(n6542), .C(n6543) );
  BUFFD0 U6426 ( .I(n6543), .Z(n6544) );
  CKBD0 U6427 ( .CLK(n6544), .C(n6545) );
  CKBD0 U6428 ( .CLK(n6545), .C(n6546) );
  CKBD0 U6429 ( .CLK(n6546), .C(n6547) );
  CKBD0 U6430 ( .CLK(n6547), .C(n6548) );
  CKBD0 U6431 ( .CLK(n6548), .C(n6549) );
  CKBD0 U6432 ( .CLK(n6549), .C(n6550) );
  CKBD0 U6433 ( .CLK(n6550), .C(n6551) );
  CKBD0 U6434 ( .CLK(n6551), .C(n6552) );
  CKBD0 U6435 ( .CLK(n6552), .C(n6553) );
  CKBD0 U6436 ( .CLK(n6553), .C(n6554) );
  BUFFD0 U6437 ( .I(n6554), .Z(n6555) );
  CKBD0 U6438 ( .CLK(n6555), .C(n6556) );
  CKBD0 U6439 ( .CLK(n6556), .C(n6557) );
  CKBD0 U6440 ( .CLK(n6557), .C(n6558) );
  CKBD0 U6441 ( .CLK(n6558), .C(n6559) );
  CKBD0 U6442 ( .CLK(n6559), .C(n6560) );
  CKBD0 U6443 ( .CLK(n6560), .C(n6561) );
  CKBD0 U6444 ( .CLK(n6561), .C(n6562) );
  CKBD0 U6445 ( .CLK(n6562), .C(n6563) );
  CKBD0 U6446 ( .CLK(n6563), .C(n6564) );
  CKBD0 U6447 ( .CLK(n6564), .C(n6565) );
  BUFFD0 U6448 ( .I(n6565), .Z(n6566) );
  CKBD0 U6449 ( .CLK(n6566), .C(n6567) );
  CKBD0 U6450 ( .CLK(n6567), .C(n6568) );
  CKBD0 U6451 ( .CLK(n6568), .C(n6569) );
  CKBD0 U6452 ( .CLK(n6569), .C(n6570) );
  CKBD0 U6453 ( .CLK(n6570), .C(n6571) );
  BUFFD0 U6454 ( .I(n6571), .Z(n6572) );
  CKBD0 U6455 ( .CLK(n6572), .C(n6573) );
  BUFFD0 U6456 ( .I(n6573), .Z(n6574) );
  CKBD0 U6457 ( .CLK(n6574), .C(n6575) );
  BUFFD0 U6458 ( .I(n6575), .Z(n6576) );
  CKBD0 U6459 ( .CLK(n6576), .C(n6577) );
  BUFFD0 U6460 ( .I(n6577), .Z(n6578) );
  CKBD0 U6461 ( .CLK(n6578), .C(n6579) );
  BUFFD0 U6462 ( .I(n6579), .Z(n6580) );
  CKBD0 U6463 ( .CLK(n6580), .C(n6581) );
  BUFFD0 U6464 ( .I(n6581), .Z(n6582) );
  CKBD0 U6465 ( .CLK(n6582), .C(n6583) );
  BUFFD0 U6466 ( .I(n6583), .Z(n6584) );
  CKBD0 U6467 ( .CLK(n6584), .C(n6585) );
  BUFFD0 U6468 ( .I(n6585), .Z(n6586) );
  BUFFD0 U6469 ( .I(n133), .Z(n6587) );
  BUFFD0 U6470 ( .I(n6589), .Z(n6588) );
  BUFFD0 U6471 ( .I(n6590), .Z(n6589) );
  BUFFD0 U6472 ( .I(Decoder[0]), .Z(n6590) );
  CKBD0 U6473 ( .CLK(n858), .C(n6591) );
  CKBD0 U6474 ( .CLK(n6591), .C(n6592) );
  CKBD0 U6475 ( .CLK(n6592), .C(n6593) );
  CKBD0 U6476 ( .CLK(n6593), .C(n6594) );
  BUFFD0 U6477 ( .I(n6594), .Z(n6595) );
  CKBD0 U6478 ( .CLK(n6595), .C(n6596) );
  CKBD0 U6479 ( .CLK(n6596), .C(n6597) );
  CKBD0 U6480 ( .CLK(n6597), .C(n6598) );
  CKBD0 U6481 ( .CLK(n6598), .C(n6599) );
  CKBD0 U6482 ( .CLK(n6599), .C(n6600) );
  CKBD0 U6483 ( .CLK(n6600), .C(n6601) );
  CKBD0 U6484 ( .CLK(n6601), .C(n6602) );
  CKBD0 U6485 ( .CLK(n6602), .C(n6603) );
  CKBD0 U6486 ( .CLK(n6603), .C(n6604) );
  BUFFD0 U6487 ( .I(n6604), .Z(n6605) );
  CKBD0 U6488 ( .CLK(n6605), .C(n6606) );
  CKBD0 U6489 ( .CLK(n6606), .C(n6607) );
  CKBD0 U6490 ( .CLK(n6607), .C(n6608) );
  CKBD0 U6491 ( .CLK(n6608), .C(n6609) );
  CKBD0 U6492 ( .CLK(n6609), .C(n6610) );
  CKBD0 U6493 ( .CLK(n6610), .C(n6611) );
  CKBD0 U6494 ( .CLK(n6611), .C(n6612) );
  CKBD0 U6495 ( .CLK(n6612), .C(n6613) );
  CKBD0 U6496 ( .CLK(n6613), .C(n6614) );
  CKBD0 U6497 ( .CLK(n6614), .C(n6615) );
  BUFFD0 U6498 ( .I(n6615), .Z(n6616) );
  CKBD0 U6499 ( .CLK(n6616), .C(n6617) );
  CKBD0 U6500 ( .CLK(n6617), .C(n6618) );
  CKBD0 U6501 ( .CLK(n6618), .C(n6619) );
  CKBD0 U6502 ( .CLK(n6619), .C(n6620) );
  CKBD0 U6503 ( .CLK(n6620), .C(n6621) );
  CKBD0 U6504 ( .CLK(n6621), .C(n6622) );
  CKBD0 U6505 ( .CLK(n6622), .C(n6623) );
  CKBD0 U6506 ( .CLK(n6623), .C(n6624) );
  CKBD0 U6507 ( .CLK(n6624), .C(n6625) );
  CKBD0 U6508 ( .CLK(n6625), .C(n6626) );
  BUFFD0 U6509 ( .I(n6626), .Z(n6627) );
  CKBD0 U6510 ( .CLK(n6627), .C(n6628) );
  CKBD0 U6511 ( .CLK(n6628), .C(n6629) );
  CKBD0 U6512 ( .CLK(n6629), .C(n6630) );
  CKBD0 U6513 ( .CLK(n6630), .C(n6631) );
  CKBD0 U6514 ( .CLK(n6631), .C(n6632) );
  CKBD0 U6515 ( .CLK(n6632), .C(n6633) );
  CKBD0 U6516 ( .CLK(n6633), .C(n6634) );
  CKBD0 U6517 ( .CLK(n6634), .C(n6635) );
  CKBD0 U6518 ( .CLK(n6635), .C(n6636) );
  CKBD0 U6519 ( .CLK(n6636), .C(n6637) );
  BUFFD0 U6520 ( .I(n6637), .Z(n6638) );
  CKBD0 U6521 ( .CLK(n6638), .C(n6639) );
  CKBD0 U6522 ( .CLK(n6639), .C(n6640) );
  CKBD0 U6523 ( .CLK(n6640), .C(n6641) );
  CKBD0 U6524 ( .CLK(n6641), .C(n6642) );
  CKBD0 U6525 ( .CLK(n6642), .C(n6643) );
  CKBD0 U6526 ( .CLK(n6643), .C(n6644) );
  CKBD0 U6527 ( .CLK(n6644), .C(n6645) );
  CKBD0 U6528 ( .CLK(n6645), .C(n6646) );
  CKBD0 U6529 ( .CLK(n6646), .C(n6647) );
  BUFFD0 U6530 ( .I(n6647), .Z(n6648) );
  CKBD0 U6531 ( .CLK(n6648), .C(n6649) );
  CKBD0 U6532 ( .CLK(n6649), .C(n6650) );
  CKBD0 U6533 ( .CLK(n6650), .C(n6651) );
  CKBD0 U6534 ( .CLK(n6651), .C(n6652) );
  CKBD0 U6535 ( .CLK(n6652), .C(n6653) );
  CKBD0 U6536 ( .CLK(n6653), .C(n6654) );
  CKBD0 U6537 ( .CLK(n6654), .C(n6655) );
  CKBD0 U6538 ( .CLK(n6655), .C(n6656) );
  CKBD0 U6539 ( .CLK(n6656), .C(n6657) );
  CKBD0 U6540 ( .CLK(n6657), .C(n6658) );
  CKBD0 U6541 ( .CLK(n6658), .C(n6659) );
  BUFFD0 U6542 ( .I(n6659), .Z(n6660) );
  CKBD0 U6543 ( .CLK(n6660), .C(n6661) );
  CKBD0 U6544 ( .CLK(n6661), .C(n6662) );
  CKBD0 U6545 ( .CLK(n6662), .C(n6663) );
  CKBD0 U6546 ( .CLK(n6663), .C(n6664) );
  CKBD0 U6547 ( .CLK(n6664), .C(n6665) );
  CKBD0 U6548 ( .CLK(n6665), .C(n6666) );
  CKBD0 U6549 ( .CLK(n6666), .C(n6667) );
  CKBD0 U6550 ( .CLK(n6667), .C(n6668) );
  CKBD0 U6551 ( .CLK(n6668), .C(n6669) );
  BUFFD0 U6552 ( .I(n6669), .Z(n6670) );
  CKBD0 U6553 ( .CLK(n6670), .C(n6671) );
  CKBD0 U6554 ( .CLK(n6671), .C(n6672) );
  CKBD0 U6555 ( .CLK(n6672), .C(n6673) );
  CKBD0 U6556 ( .CLK(n6673), .C(n6674) );
  CKBD0 U6557 ( .CLK(n6674), .C(n6675) );
  CKBD0 U6558 ( .CLK(n6675), .C(n6676) );
  CKBD0 U6559 ( .CLK(n6676), .C(n6677) );
  CKBD0 U6560 ( .CLK(n6677), .C(n6678) );
  CKBD0 U6561 ( .CLK(n6678), .C(n6679) );
  BUFFD0 U6562 ( .I(n6679), .Z(n6680) );
  CKBD0 U6563 ( .CLK(n6680), .C(n6681) );
  CKBD0 U6564 ( .CLK(n6681), .C(n6682) );
  CKBD0 U6565 ( .CLK(n6682), .C(n6683) );
  CKBD0 U6566 ( .CLK(n6683), .C(n6684) );
  CKBD0 U6567 ( .CLK(n6684), .C(n6685) );
  CKBD0 U6568 ( .CLK(n6685), .C(n6686) );
  CKBD0 U6569 ( .CLK(n6686), .C(n6687) );
  CKBD0 U6570 ( .CLK(n6687), .C(n6688) );
  CKBD0 U6571 ( .CLK(n6688), .C(n6689) );
  CKBD0 U6572 ( .CLK(n6689), .C(n6690) );
  CKBD0 U6573 ( .CLK(n6690), .C(n6691) );
  BUFFD0 U6574 ( .I(n6691), .Z(n6692) );
  CKBD0 U6575 ( .CLK(n6692), .C(n6693) );
  CKBD0 U6576 ( .CLK(n6693), .C(n6694) );
  CKBD0 U6577 ( .CLK(n6694), .C(n6695) );
  CKBD0 U6578 ( .CLK(n6695), .C(n6696) );
  CKBD0 U6579 ( .CLK(n6696), .C(n6697) );
  CKBD0 U6580 ( .CLK(n6697), .C(n6698) );
  CKBD0 U6581 ( .CLK(n6698), .C(n6699) );
  CKBD0 U6582 ( .CLK(n6699), .C(n6700) );
  CKBD0 U6583 ( .CLK(n6700), .C(n6701) );
  CKBD0 U6584 ( .CLK(n6701), .C(n6702) );
  BUFFD0 U6585 ( .I(n6702), .Z(n6703) );
  CKBD0 U6586 ( .CLK(n6703), .C(n6704) );
  CKBD0 U6587 ( .CLK(n6704), .C(n6705) );
  CKBD0 U6588 ( .CLK(n6705), .C(n6706) );
  CKBD0 U6589 ( .CLK(n6706), .C(n6707) );
  CKBD0 U6590 ( .CLK(n6707), .C(n6708) );
  BUFFD0 U6591 ( .I(n6708), .Z(n6709) );
  CKBD0 U6592 ( .CLK(n6709), .C(n6710) );
  BUFFD0 U6593 ( .I(n6710), .Z(n6711) );
  CKBD0 U6594 ( .CLK(n6711), .C(n6712) );
  BUFFD0 U6595 ( .I(n6712), .Z(n6713) );
  CKBD0 U6596 ( .CLK(n6713), .C(n6714) );
  BUFFD0 U6597 ( .I(n6714), .Z(n6715) );
  CKBD0 U6598 ( .CLK(n6715), .C(n6716) );
  BUFFD0 U6599 ( .I(n6716), .Z(n6717) );
  CKBD0 U6600 ( .CLK(n6717), .C(n6718) );
  BUFFD0 U6601 ( .I(n6718), .Z(n6719) );
  CKBD0 U6602 ( .CLK(n6719), .C(n6720) );
  BUFFD0 U6603 ( .I(n6720), .Z(n6721) );
  CKBD0 U6604 ( .CLK(n6721), .C(n6722) );
  BUFFD0 U6605 ( .I(n6722), .Z(n6723) );
  BUFFD0 U6606 ( .I(n6725), .Z(n6724) );
  BUFFD0 U6607 ( .I(n99), .Z(n6725) );
  CKND2D0 U6608 ( .A1(n232), .A2(ParValidTimer[0]), .ZN(n10) );
  XOR2D0 U6609 ( .A1(n9020), .A2(n10), .Z(n11) );
  BUFFD0 U6610 ( .I(N39), .Z(n6726) );
  CKBD0 U6611 ( .CLK(Count32[0]), .C(n6735) );
  BUFFD0 U6612 ( .I(Count32[1]), .Z(n6727) );
  BUFFD0 U6613 ( .I(n100), .Z(n6728) );
  BUFFD0 U6614 ( .I(n12), .Z(n6729) );
  CKXOR2D0 U6615 ( .A1(n232), .A2(n6), .Z(n12) );
  BUFFD0 U6616 ( .I(n6731), .Z(n6730) );
  BUFFD0 U6617 ( .I(N41), .Z(n6731) );
  BUFFD0 U6618 ( .I(n6733), .Z(n6732) );
  BUFFD0 U6619 ( .I(N40), .Z(n6733) );
  BUFFD0 U6620 ( .I(N38), .Z(n6734) );
  BUFFD0 U6621 ( .I(n6737), .Z(n6736) );
  BUFFD0 U6622 ( .I(n6738), .Z(n6737) );
  BUFFD0 U6623 ( .I(n6739), .Z(n6738) );
  BUFFD0 U6624 ( .I(n132), .Z(n6739) );
  IOA22D0 U6625 ( .B1(n9128), .B2(n63), .A1(n1), .A2(Decoder[0]), .ZN(n132) );
  BUFFD0 U6626 ( .I(n6741), .Z(n6740) );
  BUFFD0 U6627 ( .I(n6742), .Z(n6741) );
  BUFFD0 U6628 ( .I(n6743), .Z(n6742) );
  BUFFD0 U6629 ( .I(n131), .Z(n6743) );
  IOA22D0 U6630 ( .B1(n9127), .B2(n62), .A1(n1), .A2(Decoder[1]), .ZN(n131) );
  BUFFD0 U6631 ( .I(n6745), .Z(n6744) );
  BUFFD0 U6632 ( .I(n6746), .Z(n6745) );
  BUFFD0 U6633 ( .I(n6747), .Z(n6746) );
  BUFFD0 U6634 ( .I(n130), .Z(n6747) );
  IOA22D0 U6635 ( .B1(n9127), .B2(n61), .A1(n1), .A2(Decoder[2]), .ZN(n130) );
  BUFFD0 U6636 ( .I(n6749), .Z(n6748) );
  BUFFD0 U6637 ( .I(n6750), .Z(n6749) );
  BUFFD0 U6638 ( .I(n6751), .Z(n6750) );
  BUFFD0 U6639 ( .I(n129), .Z(n6751) );
  IOA22D0 U6640 ( .B1(n9127), .B2(n60), .A1(n1), .A2(Decoder[3]), .ZN(n129) );
  BUFFD0 U6641 ( .I(n6753), .Z(n6752) );
  BUFFD0 U6642 ( .I(n6754), .Z(n6753) );
  BUFFD0 U6643 ( .I(n6755), .Z(n6754) );
  BUFFD0 U6644 ( .I(n128), .Z(n6755) );
  IOA22D0 U6645 ( .B1(n9127), .B2(n59), .A1(n1), .A2(Decoder[4]), .ZN(n128) );
  BUFFD0 U6646 ( .I(n6757), .Z(n6756) );
  BUFFD0 U6647 ( .I(n6758), .Z(n6757) );
  BUFFD0 U6648 ( .I(n6759), .Z(n6758) );
  BUFFD0 U6649 ( .I(n127), .Z(n6759) );
  IOA22D0 U6650 ( .B1(n9127), .B2(n58), .A1(n1), .A2(Decoder[5]), .ZN(n127) );
  CKBD0 U6651 ( .CLK(n126), .C(n6763) );
  MOAI22D1 U6652 ( .A1(n9127), .A2(n57), .B1(n9129), .B2(Decoder[6]), .ZN(n126) );
  BUFFD0 U6653 ( .I(n6761), .Z(n6760) );
  BUFFD0 U6654 ( .I(n6762), .Z(n6761) );
  BUFFD0 U6655 ( .I(n6763), .Z(n6762) );
  IOA22D4 U6656 ( .B1(n9127), .B2(n56), .A1(n1), .A2(Decoder[7]), .ZN(n125) );
  BUFFD0 U6657 ( .I(n6765), .Z(n6764) );
  BUFFD0 U6658 ( .I(n6766), .Z(n6765) );
  BUFFD0 U6659 ( .I(n6767), .Z(n6766) );
  BUFFD0 U6660 ( .I(n125), .Z(n6767) );
  CKBD0 U6661 ( .CLK(n124), .C(n6771) );
  BUFFD0 U6662 ( .I(n6769), .Z(n6768) );
  BUFFD0 U6663 ( .I(n6770), .Z(n6769) );
  BUFFD0 U6664 ( .I(n6771), .Z(n6770) );
  CKBD0 U6665 ( .CLK(n123), .C(n6775) );
  BUFFD0 U6666 ( .I(n6773), .Z(n6772) );
  BUFFD0 U6667 ( .I(n6774), .Z(n6773) );
  BUFFD0 U6668 ( .I(n6775), .Z(n6774) );
  IOA22D4 U6669 ( .B1(n9127), .B2(n53), .A1(n9129), .A2(Decoder[10]), .ZN(n122) );
  BUFFD0 U6670 ( .I(n6777), .Z(n6776) );
  BUFFD0 U6671 ( .I(n6778), .Z(n6777) );
  BUFFD0 U6672 ( .I(n6779), .Z(n6778) );
  BUFFD0 U6673 ( .I(n122), .Z(n6779) );
  IOA22D4 U6674 ( .B1(n9127), .B2(n52), .A1(n9129), .A2(Decoder[11]), .ZN(n121) );
  BUFFD0 U6675 ( .I(n6781), .Z(n6780) );
  BUFFD0 U6676 ( .I(n6782), .Z(n6781) );
  BUFFD0 U6677 ( .I(n6783), .Z(n6782) );
  BUFFD0 U6678 ( .I(n121), .Z(n6783) );
  IOA22D4 U6679 ( .B1(n9127), .B2(n51), .A1(n9129), .A2(Decoder[12]), .ZN(n120) );
  BUFFD0 U6680 ( .I(n6785), .Z(n6784) );
  BUFFD0 U6681 ( .I(n6786), .Z(n6785) );
  BUFFD0 U6682 ( .I(n6787), .Z(n6786) );
  BUFFD0 U6683 ( .I(n120), .Z(n6787) );
  IOA22D4 U6684 ( .B1(n9127), .B2(n50), .A1(n9129), .A2(Decoder[13]), .ZN(n119) );
  BUFFD0 U6685 ( .I(n6789), .Z(n6788) );
  BUFFD0 U6686 ( .I(n6790), .Z(n6789) );
  BUFFD0 U6687 ( .I(n6791), .Z(n6790) );
  BUFFD0 U6688 ( .I(n119), .Z(n6791) );
  IOA22D4 U6689 ( .B1(n9128), .B2(n49), .A1(n9129), .A2(Decoder[14]), .ZN(n118) );
  BUFFD0 U6690 ( .I(n6793), .Z(n6792) );
  BUFFD0 U6691 ( .I(n6794), .Z(n6793) );
  BUFFD0 U6692 ( .I(n6795), .Z(n6794) );
  BUFFD0 U6693 ( .I(n118), .Z(n6795) );
  IOA22D4 U6694 ( .B1(n9128), .B2(n48), .A1(n9129), .A2(Decoder[15]), .ZN(n117) );
  BUFFD0 U6695 ( .I(n6797), .Z(n6796) );
  BUFFD0 U6696 ( .I(n6798), .Z(n6797) );
  BUFFD0 U6697 ( .I(n6799), .Z(n6798) );
  BUFFD0 U6698 ( .I(n117), .Z(n6799) );
  IOA22D4 U6699 ( .B1(n9128), .B2(n47), .A1(n9129), .A2(Decoder[16]), .ZN(n116) );
  BUFFD0 U6700 ( .I(n6801), .Z(n6800) );
  BUFFD0 U6701 ( .I(n6802), .Z(n6801) );
  BUFFD0 U6702 ( .I(n6803), .Z(n6802) );
  BUFFD0 U6703 ( .I(n116), .Z(n6803) );
  IOA22D4 U6704 ( .B1(n9128), .B2(n46), .A1(n9129), .A2(Decoder[17]), .ZN(n115) );
  BUFFD0 U6705 ( .I(n6805), .Z(n6804) );
  BUFFD0 U6706 ( .I(n6806), .Z(n6805) );
  BUFFD0 U6707 ( .I(n6807), .Z(n6806) );
  BUFFD0 U6708 ( .I(n115), .Z(n6807) );
  IOA22D4 U6709 ( .B1(n9128), .B2(n45), .A1(n9129), .A2(Decoder[18]), .ZN(n114) );
  BUFFD0 U6710 ( .I(n6809), .Z(n6808) );
  BUFFD0 U6711 ( .I(n6810), .Z(n6809) );
  BUFFD0 U6712 ( .I(n6811), .Z(n6810) );
  BUFFD0 U6713 ( .I(n114), .Z(n6811) );
  IOA22D4 U6714 ( .B1(n9128), .B2(n44), .A1(n9129), .A2(Decoder[19]), .ZN(n113) );
  BUFFD0 U6715 ( .I(n6813), .Z(n6812) );
  BUFFD0 U6716 ( .I(n6814), .Z(n6813) );
  BUFFD0 U6717 ( .I(n6815), .Z(n6814) );
  BUFFD0 U6718 ( .I(n113), .Z(n6815) );
  IOA22D4 U6719 ( .B1(n9128), .B2(n43), .A1(n9128), .A2(Decoder[20]), .ZN(n112) );
  BUFFD0 U6720 ( .I(n6817), .Z(n6816) );
  BUFFD0 U6721 ( .I(n6818), .Z(n6817) );
  BUFFD0 U6722 ( .I(n6819), .Z(n6818) );
  BUFFD0 U6723 ( .I(n112), .Z(n6819) );
  IOA22D4 U6724 ( .B1(n9128), .B2(n42), .A1(n9129), .A2(Decoder[21]), .ZN(n111) );
  BUFFD0 U6725 ( .I(n6821), .Z(n6820) );
  BUFFD0 U6726 ( .I(n6822), .Z(n6821) );
  BUFFD0 U6727 ( .I(n6823), .Z(n6822) );
  BUFFD0 U6728 ( .I(n111), .Z(n6823) );
  IOA22D4 U6729 ( .B1(n9128), .B2(n41), .A1(n9129), .A2(Decoder[22]), .ZN(n110) );
  BUFFD0 U6730 ( .I(n6825), .Z(n6824) );
  BUFFD0 U6731 ( .I(n6826), .Z(n6825) );
  BUFFD0 U6732 ( .I(n6827), .Z(n6826) );
  BUFFD0 U6733 ( .I(n110), .Z(n6827) );
  IOA22D4 U6734 ( .B1(n9128), .B2(n40), .A1(n9129), .A2(Decoder[23]), .ZN(n109) );
  BUFFD0 U6735 ( .I(n6829), .Z(n6828) );
  BUFFD0 U6736 ( .I(n6830), .Z(n6829) );
  BUFFD0 U6737 ( .I(n6831), .Z(n6830) );
  BUFFD0 U6738 ( .I(n109), .Z(n6831) );
  IOA22D4 U6739 ( .B1(n9128), .B2(n39), .A1(n9129), .A2(Decoder[24]), .ZN(n108) );
  BUFFD0 U6740 ( .I(n6833), .Z(n6832) );
  BUFFD0 U6741 ( .I(n6834), .Z(n6833) );
  BUFFD0 U6742 ( .I(n6835), .Z(n6834) );
  BUFFD0 U6743 ( .I(n108), .Z(n6835) );
  IOA22D4 U6744 ( .B1(n9128), .B2(n38), .A1(n9129), .A2(Decoder[25]), .ZN(n107) );
  BUFFD0 U6745 ( .I(n6837), .Z(n6836) );
  BUFFD0 U6746 ( .I(n6838), .Z(n6837) );
  BUFFD0 U6747 ( .I(n6839), .Z(n6838) );
  BUFFD0 U6748 ( .I(n107), .Z(n6839) );
  IOA22D4 U6749 ( .B1(n9128), .B2(n37), .A1(n9129), .A2(Decoder[26]), .ZN(n106) );
  BUFFD0 U6750 ( .I(n6841), .Z(n6840) );
  BUFFD0 U6751 ( .I(n6842), .Z(n6841) );
  BUFFD0 U6752 ( .I(n6843), .Z(n6842) );
  BUFFD0 U6753 ( .I(n106), .Z(n6843) );
  IOA22D4 U6754 ( .B1(n9128), .B2(n36), .A1(n9129), .A2(Decoder[27]), .ZN(n105) );
  BUFFD0 U6755 ( .I(n6845), .Z(n6844) );
  BUFFD0 U6756 ( .I(n6846), .Z(n6845) );
  BUFFD0 U6757 ( .I(n6847), .Z(n6846) );
  BUFFD0 U6758 ( .I(n105), .Z(n6847) );
  IOA22D4 U6759 ( .B1(n9128), .B2(n35), .A1(n1), .A2(Decoder[28]), .ZN(n104)
         );
  BUFFD0 U6760 ( .I(n6849), .Z(n6848) );
  BUFFD0 U6761 ( .I(n6850), .Z(n6849) );
  BUFFD0 U6762 ( .I(n6851), .Z(n6850) );
  BUFFD0 U6763 ( .I(n104), .Z(n6851) );
  IOA22D4 U6764 ( .B1(n9128), .B2(n34), .A1(n1), .A2(Decoder[29]), .ZN(n103)
         );
  BUFFD0 U6765 ( .I(n6853), .Z(n6852) );
  BUFFD0 U6766 ( .I(n6854), .Z(n6853) );
  BUFFD0 U6767 ( .I(n6855), .Z(n6854) );
  BUFFD0 U6768 ( .I(n103), .Z(n6855) );
  IOA22D4 U6769 ( .B1(n9128), .B2(n33), .A1(n1), .A2(Decoder[30]), .ZN(n102)
         );
  BUFFD0 U6770 ( .I(n6857), .Z(n6856) );
  BUFFD0 U6771 ( .I(n6858), .Z(n6857) );
  BUFFD0 U6772 ( .I(n6859), .Z(n6858) );
  BUFFD0 U6773 ( .I(n102), .Z(n6859) );
  BUFFD0 U6774 ( .I(n6861), .Z(n6860) );
  BUFFD0 U6775 ( .I(n6862), .Z(n6861) );
  BUFFD0 U6776 ( .I(n6863), .Z(n6862) );
  BUFFD0 U6777 ( .I(n101), .Z(n6863) );
  BUFFD0 U6778 ( .I(n6865), .Z(n6864) );
  BUFFD0 U6779 ( .I(N37), .Z(n6865) );
  BUFFD0 U6780 ( .I(n6867), .Z(n6866) );
  BUFFD0 U6781 ( .I(N43), .Z(n6867) );
  OAI21D0 U6782 ( .A1(n3), .A2(n29), .B(n231), .ZN(n96) );
  BUFFD0 U6783 ( .I(n6869), .Z(n6868) );
  BUFFD0 U6784 ( .I(n6870), .Z(n6869) );
  BUFFD0 U6785 ( .I(n6871), .Z(n6870) );
  BUFFD0 U6786 ( .I(n96), .Z(n6871) );
  NR2D0 U6787 ( .A1(n15), .A2(n14), .ZN(N47) );
  BUFFD0 U6788 ( .I(n1735), .Z(n6872) );
  CKBD0 U6789 ( .CLK(n1729), .C(n6873) );
  CKBD0 U6790 ( .CLK(n2272), .C(n6874) );
  CKBD0 U6791 ( .CLK(n1541), .C(n6875) );
  CKBD0 U6792 ( .CLK(n1360), .C(n6876) );
  CKBD0 U6793 ( .CLK(n1545), .C(n6877) );
  CKBD0 U6794 ( .CLK(n1732), .C(n6878) );
  CKBD0 U6795 ( .CLK(n1739), .C(n6879) );
  CKBD0 U6796 ( .CLK(n2006), .C(n6880) );
  CKBD0 U6797 ( .CLK(n1272), .C(n6881) );
  CKBD0 U6798 ( .CLK(n1917), .C(n6882) );
  CKBD0 U6799 ( .CLK(n2095), .C(n6883) );
  CKBD0 U6800 ( .CLK(n1257), .C(n6884) );
  CKBD0 U6801 ( .CLK(n1828), .C(n6885) );
  CKBD0 U6802 ( .CLK(n2184), .C(n6886) );
  CKBD0 U6803 ( .CLK(n856), .C(n6887) );
  CKBD0 U6804 ( .CLK(n1538), .C(n6888) );
  CKBD0 U6805 ( .CLK(n1153), .C(n6889) );
  CKBD0 U6806 ( .CLK(n219), .C(n6890) );
  BUFFD0 U6807 ( .I(n852), .Z(n6891) );
  CKBD0 U6808 ( .CLK(n1449), .C(n6892) );
  CKBD0 U6809 ( .CLK(n1724), .C(n6893) );
  CKBD0 U6810 ( .CLK(n762), .C(n6894) );
  CKBD0 U6811 ( .CLK(n959), .C(n6895) );
  CKBD0 U6812 ( .CLK(n670), .C(n6896) );
  CKBD0 U6813 ( .CLK(n1049), .C(n6897) );
  CKBD0 U6814 ( .CLK(n1634), .C(n6898) );
  CKBD0 U6815 ( .CLK(n2361), .C(n6899) );
  CKBD0 U6816 ( .CLK(n491), .C(n6900) );
  CKBD0 U6817 ( .CLK(n312), .C(n6901) );
  CKBD0 U6818 ( .CLK(n580), .C(n6902) );
  CKBD0 U6819 ( .CLK(n401), .C(n6903) );
  CKBD0 U6820 ( .CLK(n6873), .C(n6904) );
  CKBD0 U6821 ( .CLK(n6872), .C(n6905) );
  CKBD0 U6822 ( .CLK(n6874), .C(n6906) );
  CKBD0 U6823 ( .CLK(n6875), .C(n6907) );
  CKBD0 U6824 ( .CLK(n6876), .C(n6908) );
  CKBD0 U6825 ( .CLK(n6877), .C(n6909) );
  CKBD0 U6826 ( .CLK(n6878), .C(n6910) );
  CKBD0 U6827 ( .CLK(n6879), .C(n6911) );
  CKBD0 U6828 ( .CLK(n6880), .C(n6912) );
  CKBD0 U6829 ( .CLK(n6882), .C(n6913) );
  CKBD0 U6830 ( .CLK(n6881), .C(n6914) );
  CKBD0 U6831 ( .CLK(n6883), .C(n6915) );
  CKBD0 U6832 ( .CLK(n6884), .C(n6916) );
  CKBD0 U6833 ( .CLK(n6885), .C(n6917) );
  CKBD0 U6834 ( .CLK(n6886), .C(n6918) );
  CKBD0 U6835 ( .CLK(n6887), .C(n6919) );
  CKBD0 U6836 ( .CLK(n6888), .C(n6920) );
  CKBD0 U6837 ( .CLK(n6889), .C(n6921) );
  CKBD0 U6838 ( .CLK(n6891), .C(n6922) );
  BUFFD0 U6839 ( .I(n6890), .Z(n6923) );
  CKBD0 U6840 ( .CLK(n6892), .C(n6924) );
  CKBD0 U6841 ( .CLK(n6893), .C(n6925) );
  CKBD0 U6842 ( .CLK(n6894), .C(n6926) );
  CKBD0 U6843 ( .CLK(n6895), .C(n6927) );
  CKBD0 U6844 ( .CLK(n6896), .C(n6928) );
  CKBD0 U6845 ( .CLK(n6897), .C(n6929) );
  BUFFD0 U6846 ( .I(n6898), .Z(n6930) );
  CKBD0 U6847 ( .CLK(n6899), .C(n6931) );
  CKBD0 U6848 ( .CLK(n6900), .C(n6932) );
  CKBD0 U6849 ( .CLK(n6901), .C(n6933) );
  BUFFD0 U6850 ( .I(n6904), .Z(n6934) );
  CKBD0 U6851 ( .CLK(n6902), .C(n6935) );
  CKBD0 U6852 ( .CLK(n6903), .C(n6936) );
  CKBD0 U6853 ( .CLK(n6905), .C(n6937) );
  CKBD0 U6854 ( .CLK(n6906), .C(n6938) );
  CKBD0 U6855 ( .CLK(n6907), .C(n6939) );
  CKBD0 U6856 ( .CLK(n6908), .C(n6940) );
  CKBD0 U6857 ( .CLK(n6909), .C(n6941) );
  CKBD0 U6858 ( .CLK(n6910), .C(n6942) );
  CKBD0 U6859 ( .CLK(n6911), .C(n6943) );
  CKBD0 U6860 ( .CLK(n6912), .C(n6944) );
  CKBD0 U6861 ( .CLK(n6913), .C(n6945) );
  CKBD0 U6862 ( .CLK(n6914), .C(n6946) );
  CKBD0 U6863 ( .CLK(n6915), .C(n6947) );
  CKBD0 U6864 ( .CLK(n6916), .C(n6948) );
  CKBD0 U6865 ( .CLK(n6917), .C(n6949) );
  CKBD0 U6866 ( .CLK(n6918), .C(n6950) );
  CKBD0 U6867 ( .CLK(n6920), .C(n6951) );
  CKBD0 U6868 ( .CLK(n6919), .C(n6952) );
  CKBD0 U6869 ( .CLK(n6921), .C(n6953) );
  CKBD0 U6870 ( .CLK(n6922), .C(n6954) );
  CKBD0 U6871 ( .CLK(n6923), .C(n6955) );
  CKBD0 U6872 ( .CLK(n6924), .C(n6956) );
  CKBD0 U6873 ( .CLK(n6925), .C(n6957) );
  CKBD0 U6874 ( .CLK(n6926), .C(n6958) );
  CKBD0 U6875 ( .CLK(n6927), .C(n6959) );
  CKBD0 U6876 ( .CLK(n6929), .C(n6960) );
  CKBD0 U6877 ( .CLK(n6928), .C(n6961) );
  CKBD0 U6878 ( .CLK(n6930), .C(n6962) );
  CKBD0 U6879 ( .CLK(n6931), .C(n6963) );
  CKBD0 U6880 ( .CLK(n6932), .C(n6964) );
  CKBD0 U6881 ( .CLK(n6933), .C(n6965) );
  CKBD0 U6882 ( .CLK(n6934), .C(n6966) );
  CKBD0 U6883 ( .CLK(n6935), .C(n6967) );
  CKBD0 U6884 ( .CLK(n6936), .C(n6968) );
  CKBD0 U6885 ( .CLK(n6937), .C(n6969) );
  CKBD0 U6886 ( .CLK(n6938), .C(n6970) );
  CKBD0 U6887 ( .CLK(n6939), .C(n6971) );
  CKBD0 U6888 ( .CLK(n6940), .C(n6972) );
  CKBD0 U6889 ( .CLK(n6941), .C(n6973) );
  CKBD0 U6890 ( .CLK(n6942), .C(n6974) );
  CKBD0 U6891 ( .CLK(n6943), .C(n6975) );
  CKBD0 U6892 ( .CLK(n6944), .C(n6976) );
  CKBD0 U6893 ( .CLK(n6945), .C(n6977) );
  CKBD0 U6894 ( .CLK(n6947), .C(n6978) );
  CKBD0 U6895 ( .CLK(n6946), .C(n6979) );
  CKBD0 U6896 ( .CLK(n6948), .C(n6980) );
  CKBD0 U6897 ( .CLK(n6949), .C(n6981) );
  CKBD0 U6898 ( .CLK(n6950), .C(n6982) );
  CKBD0 U6899 ( .CLK(n6951), .C(n6983) );
  CKBD0 U6900 ( .CLK(n6952), .C(n6984) );
  CKBD0 U6901 ( .CLK(n6953), .C(n6985) );
  CKBD0 U6902 ( .CLK(n6954), .C(n6986) );
  CKBD0 U6903 ( .CLK(n6955), .C(n6987) );
  CKBD0 U6904 ( .CLK(n6956), .C(n6988) );
  CKBD0 U6905 ( .CLK(n6957), .C(n6989) );
  CKBD0 U6906 ( .CLK(n6958), .C(n6990) );
  CKBD0 U6907 ( .CLK(n6959), .C(n6991) );
  BUFFD0 U6908 ( .I(n6960), .Z(n6992) );
  CKBD0 U6909 ( .CLK(n6961), .C(n6993) );
  CKBD0 U6910 ( .CLK(n6962), .C(n6994) );
  BUFFD0 U6911 ( .I(n6963), .Z(n6995) );
  CKBD0 U6912 ( .CLK(n6964), .C(n6996) );
  BUFFD0 U6913 ( .I(n6967), .Z(n6997) );
  CKBD0 U6914 ( .CLK(n6965), .C(n6998) );
  CKBD0 U6915 ( .CLK(n6966), .C(n6999) );
  CKBD0 U6916 ( .CLK(n6968), .C(n7000) );
  CKBD0 U6917 ( .CLK(n6969), .C(n7001) );
  CKBD0 U6918 ( .CLK(n6970), .C(n7002) );
  CKBD0 U6919 ( .CLK(n6971), .C(n7003) );
  CKBD0 U6920 ( .CLK(n6972), .C(n7004) );
  CKBD0 U6921 ( .CLK(n6973), .C(n7005) );
  CKBD0 U6922 ( .CLK(n6974), .C(n7006) );
  CKBD0 U6923 ( .CLK(n6975), .C(n7007) );
  CKBD0 U6924 ( .CLK(n6976), .C(n7008) );
  CKBD0 U6925 ( .CLK(n6977), .C(n7009) );
  CKBD0 U6926 ( .CLK(n6979), .C(n7010) );
  CKBD0 U6927 ( .CLK(n6978), .C(n7011) );
  CKBD0 U6928 ( .CLK(n6980), .C(n7012) );
  CKBD0 U6929 ( .CLK(n6981), .C(n7013) );
  CKBD0 U6930 ( .CLK(n6982), .C(n7014) );
  CKBD0 U6931 ( .CLK(n6983), .C(n7015) );
  CKBD0 U6932 ( .CLK(n6985), .C(n7016) );
  CKBD0 U6933 ( .CLK(n6984), .C(n7017) );
  CKBD0 U6934 ( .CLK(n6986), .C(n7018) );
  CKBD0 U6935 ( .CLK(n6987), .C(n7019) );
  CKBD0 U6936 ( .CLK(n6988), .C(n7020) );
  CKBD0 U6937 ( .CLK(n6989), .C(n7021) );
  CKBD0 U6938 ( .CLK(n6990), .C(n7022) );
  CKBD0 U6939 ( .CLK(n6991), .C(n7023) );
  CKBD0 U6940 ( .CLK(n6992), .C(n7024) );
  CKBD0 U6941 ( .CLK(n6993), .C(n7025) );
  CKBD0 U6942 ( .CLK(n6994), .C(n7026) );
  CKBD0 U6943 ( .CLK(n6995), .C(n7027) );
  CKBD0 U6944 ( .CLK(n6996), .C(n7028) );
  CKBD0 U6945 ( .CLK(n6997), .C(n7029) );
  CKBD0 U6946 ( .CLK(n6998), .C(n7030) );
  CKBD0 U6947 ( .CLK(n6999), .C(n7031) );
  CKBD0 U6948 ( .CLK(n7000), .C(n7032) );
  CKBD0 U6949 ( .CLK(n7001), .C(n7033) );
  BUFFD0 U6950 ( .I(n7004), .Z(n7034) );
  CKBD0 U6951 ( .CLK(n7002), .C(n7035) );
  CKBD0 U6952 ( .CLK(n7003), .C(n7036) );
  CKBD0 U6953 ( .CLK(n7005), .C(n7037) );
  BUFFD0 U6954 ( .I(n7006), .Z(n7038) );
  CKBD0 U6955 ( .CLK(n7007), .C(n7039) );
  BUFFD0 U6956 ( .I(n7010), .Z(n7040) );
  CKBD0 U6957 ( .CLK(n7008), .C(n7041) );
  CKBD0 U6958 ( .CLK(n7009), .C(n7042) );
  CKBD0 U6959 ( .CLK(n7011), .C(n7043) );
  BUFFD0 U6960 ( .I(n7012), .Z(n7044) );
  CKBD0 U6961 ( .CLK(n7014), .C(n7045) );
  CKBD0 U6962 ( .CLK(n7013), .C(n7046) );
  CKBD0 U6963 ( .CLK(n7015), .C(n7047) );
  CKBD0 U6964 ( .CLK(n7016), .C(n7048) );
  CKBD0 U6965 ( .CLK(n7017), .C(n7049) );
  CKBD0 U6966 ( .CLK(n7018), .C(n7050) );
  CKBD0 U6967 ( .CLK(n7019), .C(n7051) );
  CKBD0 U6968 ( .CLK(n7020), .C(n7052) );
  CKBD0 U6969 ( .CLK(n7021), .C(n7053) );
  CKBD0 U6970 ( .CLK(n7022), .C(n7054) );
  CKBD0 U6971 ( .CLK(n7025), .C(n7055) );
  CKBD0 U6972 ( .CLK(n7023), .C(n7056) );
  CKBD0 U6973 ( .CLK(n7024), .C(n7057) );
  CKBD0 U6974 ( .CLK(n7026), .C(n7058) );
  CKBD0 U6975 ( .CLK(n7027), .C(n7059) );
  CKBD0 U6976 ( .CLK(n7028), .C(n7060) );
  CKBD0 U6977 ( .CLK(n7030), .C(n7061) );
  CKBD0 U6978 ( .CLK(n7029), .C(n7062) );
  CKBD0 U6979 ( .CLK(n7031), .C(n7063) );
  CKBD0 U6980 ( .CLK(n7032), .C(n7064) );
  BUFFD0 U6981 ( .I(n7036), .Z(n7065) );
  CKBD0 U6982 ( .CLK(n7033), .C(n7066) );
  CKBD0 U6983 ( .CLK(n7034), .C(n7067) );
  CKBD0 U6984 ( .CLK(n7035), .C(n7068) );
  BUFFD0 U6985 ( .I(n7037), .Z(n7069) );
  CKBD0 U6986 ( .CLK(n7038), .C(n7070) );
  CKBD0 U6987 ( .CLK(n7039), .C(n7071) );
  CKBD0 U6988 ( .CLK(n7040), .C(n7072) );
  CKBD0 U6989 ( .CLK(n7041), .C(n7073) );
  CKBD0 U6990 ( .CLK(n7042), .C(n7074) );
  CKBD0 U6991 ( .CLK(n7043), .C(n7075) );
  CKBD0 U6992 ( .CLK(n7044), .C(n7076) );
  BUFFD0 U6993 ( .I(n7045), .Z(n7077) );
  CKBD0 U6994 ( .CLK(n7046), .C(n7078) );
  CKBD0 U6995 ( .CLK(n7047), .C(n7079) );
  BUFFD0 U6996 ( .I(n7048), .Z(n7080) );
  CKBD0 U6997 ( .CLK(n7049), .C(n7081) );
  CKBD0 U6998 ( .CLK(n7050), .C(n7082) );
  CKBD0 U6999 ( .CLK(n7051), .C(n7083) );
  CKBD0 U7000 ( .CLK(n7052), .C(n7084) );
  CKBD0 U7001 ( .CLK(n7054), .C(n7085) );
  CKBD0 U7002 ( .CLK(n7053), .C(n7086) );
  CKBD0 U7003 ( .CLK(n7056), .C(n7087) );
  BUFFD0 U7004 ( .I(n7055), .Z(n7088) );
  CKBD0 U7005 ( .CLK(n7057), .C(n7089) );
  CKBD0 U7006 ( .CLK(n7058), .C(n7090) );
  CKBD0 U7007 ( .CLK(n7060), .C(n7091) );
  CKBD0 U7008 ( .CLK(n7059), .C(n7092) );
  BUFFD0 U7009 ( .I(n7061), .Z(n7093) );
  CKBD0 U7010 ( .CLK(n7062), .C(n7094) );
  CKBD0 U7011 ( .CLK(n7063), .C(n7095) );
  CKBD0 U7012 ( .CLK(n7064), .C(n7096) );
  CKBD0 U7013 ( .CLK(n7065), .C(n7097) );
  CKBD0 U7014 ( .CLK(n7066), .C(n7098) );
  CKBD0 U7015 ( .CLK(n7068), .C(n7099) );
  CKBD0 U7016 ( .CLK(n7067), .C(n7100) );
  CKBD0 U7017 ( .CLK(n7069), .C(n7101) );
  CKBD0 U7018 ( .CLK(n7070), .C(n7102) );
  BUFFD0 U7019 ( .I(n7071), .Z(n7103) );
  CKBD0 U7020 ( .CLK(n7072), .C(n7104) );
  CKBD0 U7021 ( .CLK(n7073), .C(n7105) );
  BUFFD0 U7022 ( .I(n7074), .Z(n7106) );
  CKBD0 U7023 ( .CLK(n7075), .C(n7107) );
  CKBD0 U7024 ( .CLK(n7076), .C(n7108) );
  CKBD0 U7025 ( .CLK(n7078), .C(n7109) );
  CKBD0 U7026 ( .CLK(n7077), .C(n7110) );
  BUFFD0 U7027 ( .I(n7079), .Z(n7111) );
  CKBD0 U7028 ( .CLK(n7080), .C(n7112) );
  CKBD0 U7029 ( .CLK(n7081), .C(n7113) );
  CKBD0 U7030 ( .CLK(n7082), .C(n7114) );
  CKBD0 U7031 ( .CLK(n7083), .C(n7115) );
  CKBD0 U7032 ( .CLK(n7086), .C(n7116) );
  CKBD0 U7033 ( .CLK(n7084), .C(n7117) );
  BUFFD0 U7034 ( .I(n7085), .Z(n7118) );
  BUFFD0 U7035 ( .I(n7087), .Z(n7119) );
  CKBD0 U7036 ( .CLK(n7088), .C(n7120) );
  CKBD0 U7037 ( .CLK(n7089), .C(n7121) );
  CKBD0 U7038 ( .CLK(n7090), .C(n7122) );
  CKBD0 U7039 ( .CLK(n7092), .C(n7123) );
  BUFFD0 U7040 ( .I(n7091), .Z(n7124) );
  CKBD0 U7041 ( .CLK(n7093), .C(n7125) );
  CKBD0 U7042 ( .CLK(n7094), .C(n7126) );
  CKBD0 U7043 ( .CLK(n7095), .C(n7127) );
  BUFFD0 U7044 ( .I(n7099), .Z(n7128) );
  CKBD0 U7045 ( .CLK(n7096), .C(n7129) );
  CKBD0 U7046 ( .CLK(n7097), .C(n7130) );
  CKBD0 U7047 ( .CLK(n7098), .C(n7131) );
  CKBD0 U7048 ( .CLK(n7100), .C(n7132) );
  CKBD0 U7049 ( .CLK(n7101), .C(n7133) );
  CKBD0 U7050 ( .CLK(n7102), .C(n7134) );
  CKBD0 U7051 ( .CLK(n7103), .C(n7135) );
  CKBD0 U7052 ( .CLK(n7104), .C(n7136) );
  CKBD0 U7053 ( .CLK(n7105), .C(n7137) );
  CKBD0 U7054 ( .CLK(n7106), .C(n7138) );
  BUFFD0 U7055 ( .I(n7107), .Z(n7139) );
  CKBD0 U7056 ( .CLK(n7108), .C(n7140) );
  BUFFD0 U7057 ( .I(n7113), .Z(n7141) );
  BUFFD0 U7058 ( .I(n7109), .Z(n7142) );
  CKBD0 U7059 ( .CLK(n7110), .C(n7143) );
  CKBD0 U7060 ( .CLK(n7111), .C(n7144) );
  CKBD0 U7061 ( .CLK(n7112), .C(n7145) );
  CKBD0 U7062 ( .CLK(n7114), .C(n7146) );
  CKBD0 U7063 ( .CLK(n7115), .C(n7147) );
  CKBD0 U7064 ( .CLK(n7117), .C(n7148) );
  BUFFD0 U7065 ( .I(n7116), .Z(n7149) );
  CKBD0 U7066 ( .CLK(n7118), .C(n7150) );
  CKBD0 U7067 ( .CLK(n7119), .C(n7151) );
  CKBD0 U7068 ( .CLK(n7120), .C(n7152) );
  CKBD0 U7069 ( .CLK(n7121), .C(n7153) );
  CKBD0 U7070 ( .CLK(n7122), .C(n7154) );
  CKBD0 U7071 ( .CLK(n7123), .C(n7155) );
  CKBD0 U7072 ( .CLK(n7124), .C(n7156) );
  CKBD0 U7073 ( .CLK(n7125), .C(n7157) );
  CKBD0 U7074 ( .CLK(n7126), .C(n7158) );
  BUFFD0 U7075 ( .I(n7129), .Z(n7159) );
  CKBD0 U7076 ( .CLK(n7127), .C(n7160) );
  CKBD0 U7077 ( .CLK(n7128), .C(n7161) );
  CKBD0 U7078 ( .CLK(n7130), .C(n7162) );
  CKBD0 U7079 ( .CLK(n7131), .C(n7163) );
  CKBD0 U7080 ( .CLK(n7132), .C(n7164) );
  CKBD0 U7081 ( .CLK(n7133), .C(n7165) );
  CKBD0 U7082 ( .CLK(n7134), .C(n7166) );
  CKBD0 U7083 ( .CLK(n7135), .C(n7167) );
  CKBD0 U7084 ( .CLK(n7137), .C(n7168) );
  CKBD0 U7085 ( .CLK(n7136), .C(n7169) );
  CKBD0 U7086 ( .CLK(n7138), .C(n7170) );
  CKBD0 U7087 ( .CLK(n7139), .C(n7171) );
  CKBD0 U7088 ( .CLK(n7140), .C(n7172) );
  CKBD0 U7089 ( .CLK(n7142), .C(n7173) );
  CKBD0 U7090 ( .CLK(n7143), .C(n7174) );
  CKBD0 U7091 ( .CLK(n7141), .C(n7175) );
  CKBD0 U7092 ( .CLK(n7144), .C(n7176) );
  CKBD0 U7093 ( .CLK(n7145), .C(n7177) );
  CKBD0 U7094 ( .CLK(n7146), .C(n7178) );
  CKBD0 U7095 ( .CLK(n7147), .C(n7179) );
  CKBD0 U7096 ( .CLK(n7148), .C(n7180) );
  CKBD0 U7097 ( .CLK(n7149), .C(n7181) );
  CKBD0 U7098 ( .CLK(n7150), .C(n7182) );
  CKBD0 U7099 ( .CLK(n7151), .C(n7183) );
  CKBD0 U7100 ( .CLK(n7152), .C(n7184) );
  CKBD0 U7101 ( .CLK(n7153), .C(n7185) );
  CKBD0 U7102 ( .CLK(n7154), .C(n7186) );
  CKBD0 U7103 ( .CLK(n7155), .C(n7187) );
  CKBD0 U7104 ( .CLK(n7156), .C(n7188) );
  CKBD0 U7105 ( .CLK(n7157), .C(n7189) );
  CKBD0 U7106 ( .CLK(n7158), .C(n7190) );
  CKBD0 U7107 ( .CLK(n7159), .C(n7191) );
  CKBD0 U7108 ( .CLK(n7160), .C(n7192) );
  CKBD0 U7109 ( .CLK(n7161), .C(n7193) );
  CKBD0 U7110 ( .CLK(n7162), .C(n7194) );
  CKBD0 U7111 ( .CLK(n7163), .C(n7195) );
  CKBD0 U7112 ( .CLK(n7164), .C(n7196) );
  CKBD0 U7113 ( .CLK(n7165), .C(n7197) );
  CKBD0 U7114 ( .CLK(n7166), .C(n7198) );
  CKBD0 U7115 ( .CLK(n7167), .C(n7199) );
  BUFFD0 U7116 ( .I(n7168), .Z(n7200) );
  CKBD0 U7117 ( .CLK(n7169), .C(n7201) );
  CKBD0 U7118 ( .CLK(n7170), .C(n7202) );
  CKBD0 U7119 ( .CLK(n7171), .C(n7203) );
  CKBD0 U7120 ( .CLK(n7172), .C(n7204) );
  CKBD0 U7121 ( .CLK(n7173), .C(n7205) );
  CKBD0 U7122 ( .CLK(n7174), .C(n7206) );
  CKBD0 U7123 ( .CLK(n7175), .C(n7207) );
  CKBD0 U7124 ( .CLK(n7176), .C(n7208) );
  CKBD0 U7125 ( .CLK(n7177), .C(n7209) );
  CKBD0 U7126 ( .CLK(n7178), .C(n7210) );
  CKBD0 U7127 ( .CLK(n7180), .C(n7211) );
  CKBD0 U7128 ( .CLK(n7179), .C(n7212) );
  CKBD0 U7129 ( .CLK(n7181), .C(n7213) );
  CKBD0 U7130 ( .CLK(n7182), .C(n7214) );
  CKBD0 U7131 ( .CLK(n7183), .C(n7215) );
  CKBD0 U7132 ( .CLK(n7184), .C(n7216) );
  CKBD0 U7133 ( .CLK(n7185), .C(n7217) );
  CKBD0 U7134 ( .CLK(n7186), .C(n7218) );
  CKBD0 U7135 ( .CLK(n7187), .C(n7219) );
  CKBD0 U7136 ( .CLK(n7188), .C(n7220) );
  CKBD0 U7137 ( .CLK(n7189), .C(n7221) );
  CKBD0 U7138 ( .CLK(n7190), .C(n7222) );
  CKBD0 U7139 ( .CLK(n7191), .C(n7223) );
  CKBD0 U7140 ( .CLK(n7192), .C(n7224) );
  CKBD0 U7141 ( .CLK(n7193), .C(n7225) );
  CKBD0 U7142 ( .CLK(n7195), .C(n7226) );
  CKBD0 U7143 ( .CLK(n7194), .C(n7227) );
  CKBD0 U7144 ( .CLK(n7196), .C(n7228) );
  CKBD0 U7145 ( .CLK(n7197), .C(n7229) );
  CKBD0 U7146 ( .CLK(n7198), .C(n7230) );
  CKBD0 U7147 ( .CLK(n7199), .C(n7231) );
  CKBD0 U7148 ( .CLK(n7200), .C(n7232) );
  CKBD0 U7149 ( .CLK(n7201), .C(n7233) );
  CKBD0 U7150 ( .CLK(n7202), .C(n7234) );
  CKBD0 U7151 ( .CLK(n7203), .C(n7235) );
  CKBD0 U7152 ( .CLK(n7204), .C(n7236) );
  CKBD0 U7153 ( .CLK(n7205), .C(n7237) );
  CKBD0 U7154 ( .CLK(n7206), .C(n7238) );
  CKBD0 U7155 ( .CLK(n7207), .C(n7239) );
  CKBD0 U7156 ( .CLK(n7208), .C(n7240) );
  CKBD0 U7157 ( .CLK(n7209), .C(n7241) );
  CKBD0 U7158 ( .CLK(n7212), .C(n7242) );
  BUFFD0 U7159 ( .I(n7210), .Z(n7243) );
  BUFFD0 U7160 ( .I(n7211), .Z(n7244) );
  CKBD0 U7161 ( .CLK(n7213), .C(n7245) );
  CKBD0 U7162 ( .CLK(n7214), .C(n7246) );
  CKBD0 U7163 ( .CLK(n7215), .C(n7247) );
  CKBD0 U7164 ( .CLK(n7216), .C(n7248) );
  CKBD0 U7165 ( .CLK(n7217), .C(n7249) );
  CKBD0 U7166 ( .CLK(n7218), .C(n7250) );
  CKBD0 U7167 ( .CLK(n7219), .C(n7251) );
  CKBD0 U7168 ( .CLK(n7220), .C(n7252) );
  CKBD0 U7169 ( .CLK(n7221), .C(n7253) );
  CKBD0 U7170 ( .CLK(n7222), .C(n7254) );
  CKBD0 U7171 ( .CLK(n7223), .C(n7255) );
  BUFFD0 U7172 ( .I(n7226), .Z(n7256) );
  CKBD0 U7173 ( .CLK(n7224), .C(n7257) );
  CKBD0 U7174 ( .CLK(n7225), .C(n7258) );
  CKBD0 U7175 ( .CLK(n7227), .C(n7259) );
  CKBD0 U7176 ( .CLK(n7228), .C(n7260) );
  CKBD0 U7177 ( .CLK(n7229), .C(n7261) );
  CKBD0 U7178 ( .CLK(n7230), .C(n7262) );
  CKBD0 U7179 ( .CLK(n7231), .C(n7263) );
  CKBD0 U7180 ( .CLK(n7232), .C(n7264) );
  CKBD0 U7181 ( .CLK(n7234), .C(n7265) );
  CKBD0 U7182 ( .CLK(n7233), .C(n7266) );
  CKBD0 U7183 ( .CLK(n7235), .C(n7267) );
  CKBD0 U7184 ( .CLK(n7236), .C(n7268) );
  CKBD0 U7185 ( .CLK(n7237), .C(n7269) );
  CKBD0 U7186 ( .CLK(n7238), .C(n7270) );
  CKBD0 U7187 ( .CLK(n7240), .C(n7271) );
  CKBD0 U7188 ( .CLK(n7239), .C(n7272) );
  CKBD0 U7189 ( .CLK(n7241), .C(n7273) );
  CKBD0 U7190 ( .CLK(n7243), .C(n7274) );
  BUFFD0 U7191 ( .I(n7242), .Z(n7275) );
  CKBD0 U7192 ( .CLK(n7244), .C(n7276) );
  CKBD0 U7193 ( .CLK(n7245), .C(n7277) );
  CKBD0 U7194 ( .CLK(n7246), .C(n7278) );
  CKBD0 U7195 ( .CLK(n7247), .C(n7279) );
  CKBD0 U7196 ( .CLK(n7248), .C(n7280) );
  CKBD0 U7197 ( .CLK(n7249), .C(n7281) );
  BUFFD0 U7198 ( .I(n7250), .Z(n7282) );
  CKBD0 U7199 ( .CLK(n7251), .C(n7283) );
  CKBD0 U7200 ( .CLK(n7252), .C(n7284) );
  CKBD0 U7201 ( .CLK(n7253), .C(n7285) );
  CKBD0 U7202 ( .CLK(n7254), .C(n7286) );
  CKBD0 U7203 ( .CLK(n7255), .C(n7287) );
  CKBD0 U7204 ( .CLK(n7257), .C(n7288) );
  CKBD0 U7205 ( .CLK(n7256), .C(n7289) );
  CKBD0 U7206 ( .CLK(n7258), .C(n7290) );
  CKBD0 U7207 ( .CLK(n7259), .C(n7291) );
  CKBD0 U7208 ( .CLK(n7260), .C(n7292) );
  CKBD0 U7209 ( .CLK(n7261), .C(n7293) );
  CKBD0 U7210 ( .CLK(n7262), .C(n7294) );
  CKBD0 U7211 ( .CLK(n7263), .C(n7295) );
  CKBD0 U7212 ( .CLK(n7264), .C(n7296) );
  CKBD0 U7213 ( .CLK(n7265), .C(n7297) );
  CKBD0 U7214 ( .CLK(n7266), .C(n7298) );
  CKBD0 U7215 ( .CLK(n7267), .C(n7299) );
  CKBD0 U7216 ( .CLK(n7268), .C(n7300) );
  CKBD0 U7217 ( .CLK(n7269), .C(n7301) );
  CKBD0 U7218 ( .CLK(n7270), .C(n7302) );
  CKBD0 U7219 ( .CLK(n7271), .C(n7303) );
  CKBD0 U7220 ( .CLK(n7272), .C(n7304) );
  CKBD0 U7221 ( .CLK(n7273), .C(n7305) );
  CKBD0 U7222 ( .CLK(n7274), .C(n7306) );
  CKBD0 U7223 ( .CLK(n7275), .C(n7307) );
  CKBD0 U7224 ( .CLK(n7276), .C(n7308) );
  CKBD0 U7225 ( .CLK(n7277), .C(n7309) );
  CKBD0 U7226 ( .CLK(n7278), .C(n7310) );
  CKBD0 U7227 ( .CLK(n7279), .C(n7311) );
  CKBD0 U7228 ( .CLK(n7281), .C(n7312) );
  CKBD0 U7229 ( .CLK(n7280), .C(n7313) );
  CKBD0 U7230 ( .CLK(n7282), .C(n7314) );
  BUFFD0 U7231 ( .I(n7283), .Z(n7315) );
  CKBD0 U7232 ( .CLK(n7284), .C(n7316) );
  CKBD0 U7233 ( .CLK(n7285), .C(n7317) );
  BUFFD0 U7234 ( .I(n7288), .Z(n7318) );
  CKBD0 U7235 ( .CLK(n7286), .C(n7319) );
  CKBD0 U7236 ( .CLK(n7287), .C(n7320) );
  CKBD0 U7237 ( .CLK(n7289), .C(n7321) );
  CKBD0 U7238 ( .CLK(n7290), .C(n7322) );
  CKBD0 U7239 ( .CLK(n7291), .C(n7323) );
  CKBD0 U7240 ( .CLK(n7292), .C(n7324) );
  CKBD0 U7241 ( .CLK(n7293), .C(n7325) );
  CKBD0 U7242 ( .CLK(n7294), .C(n7326) );
  CKBD0 U7243 ( .CLK(n7295), .C(n7327) );
  CKBD0 U7244 ( .CLK(n7296), .C(n7328) );
  CKBD0 U7245 ( .CLK(n7297), .C(n7329) );
  CKBD0 U7246 ( .CLK(n7299), .C(n7330) );
  CKBD0 U7247 ( .CLK(n7298), .C(n7331) );
  CKBD0 U7248 ( .CLK(n7300), .C(n7332) );
  CKBD0 U7249 ( .CLK(n7301), .C(n7333) );
  CKBD0 U7250 ( .CLK(n7302), .C(n7334) );
  CKBD0 U7251 ( .CLK(n7303), .C(n7335) );
  CKBD0 U7252 ( .CLK(n7304), .C(n7336) );
  CKBD0 U7253 ( .CLK(n7305), .C(n7337) );
  CKBD0 U7254 ( .CLK(n7306), .C(n7338) );
  CKBD0 U7255 ( .CLK(n7307), .C(n7339) );
  CKBD0 U7256 ( .CLK(n7308), .C(n7340) );
  CKBD0 U7257 ( .CLK(n7309), .C(n7341) );
  CKBD0 U7258 ( .CLK(n7310), .C(n7342) );
  CKBD0 U7259 ( .CLK(n7311), .C(n7343) );
  BUFFD0 U7260 ( .I(n7312), .Z(n7344) );
  CKBD0 U7261 ( .CLK(n7313), .C(n7345) );
  CKBD0 U7262 ( .CLK(n7314), .C(n7346) );
  CKBD0 U7263 ( .CLK(n7315), .C(n7347) );
  CKBD0 U7264 ( .CLK(n7316), .C(n7348) );
  CKBD0 U7265 ( .CLK(n7317), .C(n7349) );
  CKBD0 U7266 ( .CLK(n7318), .C(n7350) );
  CKBD0 U7267 ( .CLK(n7319), .C(n7351) );
  CKBD0 U7268 ( .CLK(n7320), .C(n7352) );
  CKBD0 U7269 ( .CLK(n7321), .C(n7353) );
  CKBD0 U7270 ( .CLK(n7322), .C(n7354) );
  CKBD0 U7271 ( .CLK(n7323), .C(n7355) );
  CKBD0 U7272 ( .CLK(n7324), .C(n7356) );
  CKBD0 U7273 ( .CLK(n7325), .C(n7357) );
  BUFFD0 U7274 ( .I(n7326), .Z(n7358) );
  CKBD0 U7275 ( .CLK(n7327), .C(n7359) );
  CKBD0 U7276 ( .CLK(n7328), .C(n7360) );
  CKBD0 U7277 ( .CLK(n7329), .C(n7361) );
  CKBD0 U7278 ( .CLK(n7331), .C(n7362) );
  CKBD0 U7279 ( .CLK(n7330), .C(n7363) );
  CKBD0 U7280 ( .CLK(n7332), .C(n7364) );
  CKBD0 U7281 ( .CLK(n7333), .C(n7365) );
  CKBD0 U7282 ( .CLK(n7334), .C(n7366) );
  CKBD0 U7283 ( .CLK(n7335), .C(n7367) );
  CKBD0 U7284 ( .CLK(n7337), .C(n7368) );
  CKBD0 U7285 ( .CLK(n7336), .C(n7369) );
  CKBD0 U7286 ( .CLK(n7338), .C(n7370) );
  CKBD0 U7287 ( .CLK(n7339), .C(n7371) );
  CKBD0 U7288 ( .CLK(n7340), .C(n7372) );
  CKBD0 U7289 ( .CLK(n7341), .C(n7373) );
  CKBD0 U7290 ( .CLK(n7342), .C(n7374) );
  CKBD0 U7291 ( .CLK(n7343), .C(n7375) );
  CKBD0 U7292 ( .CLK(n7344), .C(n7376) );
  CKBD0 U7293 ( .CLK(n7345), .C(n7377) );
  CKBD0 U7294 ( .CLK(n7346), .C(n7378) );
  CKBD0 U7295 ( .CLK(n7347), .C(n7379) );
  CKBD0 U7296 ( .CLK(n7348), .C(n7380) );
  CKBD0 U7297 ( .CLK(n7349), .C(n7381) );
  CKBD0 U7298 ( .CLK(n7350), .C(n7382) );
  CKBD0 U7299 ( .CLK(n7351), .C(n7383) );
  CKBD0 U7300 ( .CLK(n7352), .C(n7384) );
  CKBD0 U7301 ( .CLK(n7353), .C(n7385) );
  BUFFD0 U7302 ( .I(n7356), .Z(n7386) );
  CKBD0 U7303 ( .CLK(n7354), .C(n7387) );
  CKBD0 U7304 ( .CLK(n7355), .C(n7388) );
  CKBD0 U7305 ( .CLK(n7357), .C(n7389) );
  CKBD0 U7306 ( .CLK(n7358), .C(n7390) );
  CKBD0 U7307 ( .CLK(n7359), .C(n7391) );
  BUFFD0 U7308 ( .I(n7362), .Z(n7392) );
  CKBD0 U7309 ( .CLK(n7360), .C(n7393) );
  CKBD0 U7310 ( .CLK(n7361), .C(n7394) );
  CKBD0 U7311 ( .CLK(n7363), .C(n7395) );
  BUFFD0 U7312 ( .I(n7364), .Z(n7396) );
  CKBD0 U7313 ( .CLK(n7366), .C(n7397) );
  CKBD0 U7314 ( .CLK(n7365), .C(n7398) );
  CKBD0 U7315 ( .CLK(n7367), .C(n7399) );
  BUFFD0 U7316 ( .I(n7368), .Z(n7400) );
  CKBD0 U7317 ( .CLK(n7369), .C(n7401) );
  CKBD0 U7318 ( .CLK(n7370), .C(n7402) );
  CKBD0 U7319 ( .CLK(n7371), .C(n7403) );
  CKBD0 U7320 ( .CLK(n7372), .C(n7404) );
  CKBD0 U7321 ( .CLK(n7373), .C(n7405) );
  CKBD0 U7322 ( .CLK(n7374), .C(n7406) );
  CKBD0 U7323 ( .CLK(n7377), .C(n7407) );
  CKBD0 U7324 ( .CLK(n7375), .C(n7408) );
  CKBD0 U7325 ( .CLK(n7376), .C(n7409) );
  CKBD0 U7326 ( .CLK(n7378), .C(n7410) );
  CKBD0 U7327 ( .CLK(n7379), .C(n7411) );
  CKBD0 U7328 ( .CLK(n7380), .C(n7412) );
  CKBD0 U7329 ( .CLK(n7381), .C(n7413) );
  CKBD0 U7330 ( .CLK(n7382), .C(n7414) );
  CKBD0 U7331 ( .CLK(n7383), .C(n7415) );
  CKBD0 U7332 ( .CLK(n7384), .C(n7416) );
  BUFFD0 U7333 ( .I(n7388), .Z(n7417) );
  CKBD0 U7334 ( .CLK(n7385), .C(n7418) );
  CKBD0 U7335 ( .CLK(n7386), .C(n7419) );
  CKBD0 U7336 ( .CLK(n7387), .C(n7420) );
  CKBD0 U7337 ( .CLK(n7389), .C(n7421) );
  CKBD0 U7338 ( .CLK(n7390), .C(n7422) );
  CKBD0 U7339 ( .CLK(n7391), .C(n7423) );
  CKBD0 U7340 ( .CLK(n7392), .C(n7424) );
  CKBD0 U7341 ( .CLK(n7393), .C(n7425) );
  CKBD0 U7342 ( .CLK(n7394), .C(n7426) );
  CKBD0 U7343 ( .CLK(n7395), .C(n7427) );
  CKBD0 U7344 ( .CLK(n7396), .C(n7428) );
  BUFFD0 U7345 ( .I(n7397), .Z(n7429) );
  CKBD0 U7346 ( .CLK(n7398), .C(n7430) );
  CKBD0 U7347 ( .CLK(n7399), .C(n7431) );
  CKBD0 U7348 ( .CLK(n7400), .C(n7432) );
  CKBD0 U7349 ( .CLK(n7401), .C(n7433) );
  CKBD0 U7350 ( .CLK(n7402), .C(n7434) );
  CKBD0 U7351 ( .CLK(n7403), .C(n7435) );
  CKBD0 U7352 ( .CLK(n7404), .C(n7436) );
  CKBD0 U7353 ( .CLK(n7406), .C(n7437) );
  CKBD0 U7354 ( .CLK(n7405), .C(n7438) );
  CKBD0 U7355 ( .CLK(n7408), .C(n7439) );
  BUFFD0 U7356 ( .I(n7407), .Z(n7440) );
  CKBD0 U7357 ( .CLK(n7409), .C(n7441) );
  CKBD0 U7358 ( .CLK(n7410), .C(n7442) );
  CKBD0 U7359 ( .CLK(n7412), .C(n7443) );
  CKBD0 U7360 ( .CLK(n7411), .C(n7444) );
  BUFFD0 U7361 ( .I(n7413), .Z(n7445) );
  BUFFD0 U7362 ( .I(n7415), .Z(n7446) );
  CKBD0 U7363 ( .CLK(n7414), .C(n7447) );
  CKBD0 U7364 ( .CLK(n7416), .C(n7448) );
  CKBD0 U7365 ( .CLK(n7417), .C(n7449) );
  CKBD0 U7366 ( .CLK(n7418), .C(n7450) );
  CKBD0 U7367 ( .CLK(n7419), .C(n7451) );
  CKBD0 U7368 ( .CLK(n7420), .C(n7452) );
  BUFFD0 U7369 ( .I(n7421), .Z(n7453) );
  CKBD0 U7370 ( .CLK(n7422), .C(n7454) );
  BUFFD0 U7371 ( .I(n7423), .Z(n7455) );
  CKBD0 U7372 ( .CLK(n7424), .C(n7456) );
  CKBD0 U7373 ( .CLK(n7425), .C(n7457) );
  BUFFD0 U7374 ( .I(n7426), .Z(n7458) );
  CKBD0 U7375 ( .CLK(n7427), .C(n7459) );
  CKBD0 U7376 ( .CLK(n7428), .C(n7460) );
  CKBD0 U7377 ( .CLK(n7430), .C(n7461) );
  CKBD0 U7378 ( .CLK(n7429), .C(n7462) );
  BUFFD0 U7379 ( .I(n7431), .Z(n7463) );
  CKBD0 U7380 ( .CLK(n7432), .C(n7464) );
  CKBD0 U7381 ( .CLK(n7433), .C(n7465) );
  CKBD0 U7382 ( .CLK(n7434), .C(n7466) );
  CKBD0 U7383 ( .CLK(n7435), .C(n7467) );
  CKBD0 U7384 ( .CLK(n7438), .C(n7468) );
  CKBD0 U7385 ( .CLK(n7436), .C(n7469) );
  BUFFD0 U7386 ( .I(n7437), .Z(n7470) );
  CKBD0 U7387 ( .CLK(n7439), .C(n7471) );
  CKBD0 U7388 ( .CLK(n7440), .C(n7472) );
  CKBD0 U7389 ( .CLK(n7441), .C(n7473) );
  CKBD0 U7390 ( .CLK(n7442), .C(n7474) );
  CKBD0 U7391 ( .CLK(n7444), .C(n7475) );
  BUFFD0 U7392 ( .I(n7443), .Z(n7476) );
  CKBD0 U7393 ( .CLK(n7445), .C(n7477) );
  CKBD0 U7394 ( .CLK(n7446), .C(n7478) );
  CKBD0 U7395 ( .CLK(n7447), .C(n7479) );
  CKBD0 U7396 ( .CLK(n7448), .C(n7480) );
  CKBD0 U7397 ( .CLK(n7449), .C(n7481) );
  CKBD0 U7398 ( .CLK(n7450), .C(n7482) );
  CKBD0 U7399 ( .CLK(n7452), .C(n7483) );
  CKBD0 U7400 ( .CLK(n7451), .C(n7484) );
  CKBD0 U7401 ( .CLK(n7453), .C(n7485) );
  CKBD0 U7402 ( .CLK(n7454), .C(n7486) );
  CKBD0 U7403 ( .CLK(n7457), .C(n7487) );
  CKBD0 U7404 ( .CLK(n7458), .C(n7488) );
  BUFFD0 U7405 ( .I(n7459), .Z(n7489) );
  CKBD0 U7406 ( .CLK(n7460), .C(n7490) );
  BUFFD0 U7407 ( .I(n7461), .Z(n7491) );
  CKBD0 U7408 ( .CLK(n7462), .C(n7492) );
  CKBD0 U7409 ( .CLK(n7463), .C(n7493) );
  CKBD0 U7410 ( .CLK(n7464), .C(n7494) );
  CKBD0 U7411 ( .CLK(n7455), .C(n7495) );
  CKBD0 U7412 ( .CLK(n7456), .C(n7496) );
  CKBD0 U7413 ( .CLK(n7466), .C(n7497) );
  CKBD0 U7414 ( .CLK(n7467), .C(n7498) );
  CKBD0 U7415 ( .CLK(n7469), .C(n7499) );
  BUFFD0 U7416 ( .I(n7468), .Z(n7500) );
  CKBD0 U7417 ( .CLK(n7470), .C(n7501) );
  CKBD0 U7418 ( .CLK(n7471), .C(n7502) );
  CKBD0 U7419 ( .CLK(n7472), .C(n7503) );
  CKBD0 U7420 ( .CLK(n7473), .C(n7504) );
  BUFFD0 U7421 ( .I(n7465), .Z(n7505) );
  CKBD0 U7422 ( .CLK(n7474), .C(n7506) );
  CKBD0 U7423 ( .CLK(n7475), .C(n7507) );
  CKBD0 U7424 ( .CLK(n7476), .C(n7508) );
  CKBD0 U7425 ( .CLK(n7477), .C(n7509) );
  CKBD0 U7426 ( .CLK(n7478), .C(n7510) );
  CKBD0 U7427 ( .CLK(n7479), .C(n7511) );
  CKBD0 U7428 ( .CLK(n7481), .C(n7512) );
  CKBD0 U7429 ( .CLK(n7482), .C(n7513) );
  CKBD0 U7430 ( .CLK(n7485), .C(n7514) );
  CKBD0 U7431 ( .CLK(n7486), .C(n7515) );
  CKBD0 U7432 ( .CLK(n7495), .C(n7516) );
  CKBD0 U7433 ( .CLK(n7496), .C(n7517) );
  BUFFD0 U7434 ( .I(n7480), .Z(n7518) );
  BUFFD0 U7435 ( .I(n7483), .Z(n7519) );
  CKBD0 U7436 ( .CLK(n7505), .C(n7520) );
  CKBD0 U7437 ( .CLK(n7484), .C(n7521) );
  CKBD0 U7438 ( .CLK(n7511), .C(n7522) );
  CKBD0 U7439 ( .CLK(n7513), .C(n7523) );
  CKBD0 U7440 ( .CLK(n7512), .C(n7524) );
  BUFFD0 U7441 ( .I(n7487), .Z(n7525) );
  CKBD0 U7442 ( .CLK(n7514), .C(n7526) );
  CKBD0 U7443 ( .CLK(n7488), .C(n7527) );
  CKBD0 U7444 ( .CLK(n7489), .C(n7528) );
  CKBD0 U7445 ( .CLK(n7490), .C(n7529) );
  CKBD0 U7446 ( .CLK(n7491), .C(n7530) );
  CKBD0 U7447 ( .CLK(n7492), .C(n7531) );
  CKBD0 U7448 ( .CLK(n7493), .C(n7532) );
  CKBD0 U7449 ( .CLK(n7515), .C(n7533) );
  CKBD0 U7450 ( .CLK(n7494), .C(n7534) );
  CKBD0 U7451 ( .CLK(n7497), .C(n7535) );
  CKBD0 U7452 ( .CLK(n7498), .C(n7536) );
  CKBD0 U7453 ( .CLK(n7499), .C(n7537) );
  CKBD0 U7454 ( .CLK(n7500), .C(n7538) );
  CKBD0 U7455 ( .CLK(n7501), .C(n7539) );
  CKBD0 U7456 ( .CLK(n7516), .C(n7540) );
  BUFFD0 U7457 ( .I(n7502), .Z(n7541) );
  CKBD0 U7458 ( .CLK(n7517), .C(n7542) );
  CKBD0 U7459 ( .CLK(n7520), .C(n7543) );
  CKBD0 U7460 ( .CLK(n7522), .C(n7544) );
  BUFFD0 U7461 ( .I(n7523), .Z(n7545) );
  CKBD0 U7462 ( .CLK(n7524), .C(n7546) );
  CKBD0 U7463 ( .CLK(n7526), .C(n7547) );
  CKBD0 U7464 ( .CLK(n7533), .C(n7548) );
  CKBD0 U7465 ( .CLK(n7503), .C(n7549) );
  CKBD0 U7466 ( .CLK(n7504), .C(n7550) );
  CKBD0 U7467 ( .CLK(n7506), .C(n7551) );
  CKBD0 U7468 ( .CLK(n7507), .C(n7552) );
  CKBD0 U7469 ( .CLK(n7508), .C(n7553) );
  CKBD0 U7470 ( .CLK(n7540), .C(n7554) );
  CKBD0 U7471 ( .CLK(n7542), .C(n7555) );
  CKBD0 U7472 ( .CLK(n7543), .C(n7556) );
  BUFFD0 U7473 ( .I(n7544), .Z(n7557) );
  CKBD0 U7474 ( .CLK(n7545), .C(n7558) );
  CKBD0 U7475 ( .CLK(n7546), .C(n7559) );
  CKBD0 U7476 ( .CLK(n7547), .C(n7560) );
  CKBD0 U7477 ( .CLK(n7548), .C(n7561) );
  CKBD0 U7478 ( .CLK(n7509), .C(n7562) );
  CKBD0 U7479 ( .CLK(n7510), .C(n7563) );
  CKBD0 U7480 ( .CLK(n7554), .C(n7564) );
  CKBD0 U7481 ( .CLK(n7518), .C(n7565) );
  CKBD0 U7482 ( .CLK(n7519), .C(n7566) );
  CKBD0 U7483 ( .CLK(n7521), .C(n7567) );
  CKBD0 U7484 ( .CLK(n7555), .C(n7568) );
  CKBD0 U7485 ( .CLK(n7556), .C(n7569) );
  CKBD0 U7486 ( .CLK(n7557), .C(n7570) );
  CKBD0 U7487 ( .CLK(n7525), .C(n7571) );
  CKBD0 U7488 ( .CLK(n7527), .C(n7572) );
  CKBD0 U7489 ( .CLK(n7528), .C(n7573) );
  CKBD0 U7490 ( .CLK(n7558), .C(n7574) );
  CKBD0 U7491 ( .CLK(n7529), .C(n7575) );
  CKBD0 U7492 ( .CLK(n7530), .C(n7576) );
  CKBD0 U7493 ( .CLK(n7531), .C(n7577) );
  CKBD0 U7494 ( .CLK(n7532), .C(n7578) );
  CKBD0 U7495 ( .CLK(n7559), .C(n7579) );
  CKBD0 U7496 ( .CLK(n7534), .C(n7580) );
  CKBD0 U7497 ( .CLK(n7535), .C(n7581) );
  CKBD0 U7498 ( .CLK(n7537), .C(n7582) );
  CKBD0 U7499 ( .CLK(n7536), .C(n7583) );
  CKBD0 U7500 ( .CLK(n7538), .C(n7584) );
  CKBD0 U7501 ( .CLK(n7539), .C(n7585) );
  CKBD0 U7502 ( .CLK(n7560), .C(n7586) );
  CKBD0 U7503 ( .CLK(n7541), .C(n7587) );
  CKBD0 U7504 ( .CLK(n7549), .C(n7588) );
  CKBD0 U7505 ( .CLK(n7550), .C(n7589) );
  CKBD0 U7506 ( .CLK(n7551), .C(n7590) );
  CKBD0 U7507 ( .CLK(n7552), .C(n7591) );
  CKBD0 U7508 ( .CLK(n7553), .C(n7592) );
  CKBD0 U7509 ( .CLK(n7561), .C(n7593) );
  CKBD0 U7510 ( .CLK(n7562), .C(n7594) );
  CKBD0 U7511 ( .CLK(n7563), .C(n7595) );
  CKBD0 U7512 ( .CLK(n7564), .C(n7596) );
  CKBD0 U7513 ( .CLK(n7565), .C(n7597) );
  CKBD0 U7514 ( .CLK(n7566), .C(n7598) );
  CKBD0 U7515 ( .CLK(n7567), .C(n7599) );
  CKBD0 U7516 ( .CLK(n7568), .C(n7600) );
  CKBD0 U7517 ( .CLK(n7569), .C(n7601) );
  CKBD0 U7518 ( .CLK(n7570), .C(n7602) );
  CKBD0 U7519 ( .CLK(n7571), .C(n7603) );
  CKBD0 U7520 ( .CLK(n7572), .C(n7604) );
  CKBD0 U7521 ( .CLK(n7573), .C(n7605) );
  CKBD0 U7522 ( .CLK(n7574), .C(n7606) );
  CKBD0 U7523 ( .CLK(n7575), .C(n7607) );
  CKBD0 U7524 ( .CLK(n7576), .C(n7608) );
  CKBD0 U7525 ( .CLK(n7577), .C(n7609) );
  CKBD0 U7526 ( .CLK(n7578), .C(n7610) );
  CKBD0 U7527 ( .CLK(n7580), .C(n7611) );
  CKBD0 U7528 ( .CLK(n7579), .C(n7612) );
  BUFFD0 U7529 ( .I(n7581), .Z(n7613) );
  BUFFD0 U7530 ( .I(n7582), .Z(n7614) );
  CKBD0 U7531 ( .CLK(n7583), .C(n7615) );
  CKBD0 U7532 ( .CLK(n7584), .C(n7616) );
  CKBD0 U7533 ( .CLK(n7585), .C(n7617) );
  CKBD0 U7534 ( .CLK(n7587), .C(n7618) );
  CKBD0 U7535 ( .CLK(n7586), .C(n7619) );
  CKBD0 U7536 ( .CLK(n7588), .C(n7620) );
  BUFFD0 U7537 ( .I(n7593), .Z(n7621) );
  CKBD0 U7538 ( .CLK(n7589), .C(n7622) );
  BUFFD0 U7539 ( .I(n7590), .Z(n7623) );
  CKBD0 U7540 ( .CLK(n7591), .C(n7624) );
  CKBD0 U7541 ( .CLK(n7592), .C(n7625) );
  CKBD0 U7542 ( .CLK(n7594), .C(n7626) );
  CKBD0 U7543 ( .CLK(n7595), .C(n7627) );
  CKBD0 U7544 ( .CLK(n7596), .C(n7628) );
  CKBD0 U7545 ( .CLK(n7597), .C(n7629) );
  CKBD0 U7546 ( .CLK(n7598), .C(n7630) );
  CKBD0 U7547 ( .CLK(n7599), .C(n7631) );
  CKBD0 U7548 ( .CLK(n7600), .C(n7632) );
  CKBD0 U7549 ( .CLK(n7601), .C(n7633) );
  CKBD0 U7550 ( .CLK(n7602), .C(n7634) );
  CKBD0 U7551 ( .CLK(n7603), .C(n7635) );
  CKBD0 U7552 ( .CLK(n7604), .C(n7636) );
  CKBD0 U7553 ( .CLK(n7605), .C(n7637) );
  CKBD0 U7554 ( .CLK(n7606), .C(n7638) );
  CKBD0 U7555 ( .CLK(n7612), .C(n7639) );
  CKBD0 U7556 ( .CLK(n7619), .C(n7640) );
  CKBD0 U7557 ( .CLK(n7621), .C(n7641) );
  CKBD0 U7558 ( .CLK(n7628), .C(n7642) );
  CKBD0 U7559 ( .CLK(n7632), .C(n7643) );
  CKBD0 U7560 ( .CLK(n7633), .C(n7644) );
  CKBD0 U7561 ( .CLK(n7634), .C(n7645) );
  CKBD0 U7562 ( .CLK(n7607), .C(n7646) );
  CKBD0 U7563 ( .CLK(n7608), .C(n7647) );
  CKBD0 U7564 ( .CLK(n7609), .C(n7648) );
  CKBD0 U7565 ( .CLK(n7610), .C(n7649) );
  CKBD0 U7566 ( .CLK(n7611), .C(n7650) );
  CKBD0 U7567 ( .CLK(n7638), .C(n7651) );
  CKBD0 U7568 ( .CLK(n7639), .C(n7652) );
  CKBD0 U7569 ( .CLK(n7640), .C(n7653) );
  CKBD0 U7570 ( .CLK(n7641), .C(n7654) );
  BUFFD0 U7571 ( .I(n7642), .Z(n7655) );
  BUFFD0 U7572 ( .I(n7643), .Z(n7656) );
  CKBD0 U7573 ( .CLK(n7644), .C(n7657) );
  CKBD0 U7574 ( .CLK(n7645), .C(n7658) );
  CKBD0 U7575 ( .CLK(n7615), .C(n7659) );
  CKBD0 U7576 ( .CLK(n7613), .C(n7660) );
  CKBD0 U7577 ( .CLK(n7651), .C(n7661) );
  CKBD0 U7578 ( .CLK(n7652), .C(n7662) );
  BUFFD0 U7579 ( .I(n7653), .Z(n7663) );
  CKBD0 U7580 ( .CLK(n7654), .C(n7664) );
  CKBD0 U7581 ( .CLK(n7655), .C(n7665) );
  CKBD0 U7582 ( .CLK(n7656), .C(n7666) );
  CKBD0 U7583 ( .CLK(n7657), .C(n7667) );
  CKBD0 U7584 ( .CLK(n7658), .C(n7668) );
  BUFFD0 U7585 ( .I(n7662), .Z(n7669) );
  CKBD0 U7586 ( .CLK(n7661), .C(n7670) );
  CKBD0 U7587 ( .CLK(n7663), .C(n7671) );
  CKBD0 U7588 ( .CLK(n7664), .C(n7672) );
  CKBD0 U7589 ( .CLK(n7665), .C(n7673) );
  CKBD0 U7590 ( .CLK(n7666), .C(n7674) );
  BUFFD0 U7591 ( .I(n7667), .Z(n7675) );
  CKBD0 U7592 ( .CLK(n7668), .C(n7676) );
  CKBD0 U7593 ( .CLK(n7669), .C(n7677) );
  CKBD0 U7594 ( .CLK(n7670), .C(n7678) );
  CKBD0 U7595 ( .CLK(n7671), .C(n7679) );
  CKBD0 U7596 ( .CLK(n7672), .C(n7680) );
  CKBD0 U7597 ( .CLK(n7673), .C(n7681) );
  CKBD0 U7598 ( .CLK(n7674), .C(n7682) );
  CKBD0 U7599 ( .CLK(n7675), .C(n7683) );
  CKBD0 U7600 ( .CLK(n7676), .C(n7684) );
  CKBD0 U7601 ( .CLK(n7677), .C(n7685) );
  CKBD0 U7602 ( .CLK(n7678), .C(n7686) );
  CKBD0 U7603 ( .CLK(n7679), .C(n7687) );
  CKBD0 U7604 ( .CLK(n7680), .C(n7688) );
  CKBD0 U7605 ( .CLK(n7681), .C(n7689) );
  CKBD0 U7606 ( .CLK(n7682), .C(n7690) );
  CKBD0 U7607 ( .CLK(n7683), .C(n7691) );
  CKBD0 U7608 ( .CLK(n7614), .C(n7692) );
  CKBD0 U7609 ( .CLK(n7684), .C(n7693) );
  CKBD0 U7610 ( .CLK(n7686), .C(n7694) );
  CKBD0 U7611 ( .CLK(n7685), .C(n7695) );
  CKBD0 U7612 ( .CLK(n7687), .C(n7696) );
  CKBD0 U7613 ( .CLK(n7688), .C(n7697) );
  CKBD0 U7614 ( .CLK(n7689), .C(n7698) );
  CKBD0 U7615 ( .CLK(n7690), .C(n7699) );
  CKBD0 U7616 ( .CLK(n7616), .C(n7700) );
  CKBD0 U7617 ( .CLK(n7617), .C(n7701) );
  CKBD0 U7618 ( .CLK(n7618), .C(n7702) );
  CKBD0 U7619 ( .CLK(n7620), .C(n7703) );
  CKBD0 U7620 ( .CLK(n7622), .C(n7704) );
  CKBD0 U7621 ( .CLK(n7623), .C(n7705) );
  CKBD0 U7622 ( .CLK(n7691), .C(n7706) );
  CKBD0 U7623 ( .CLK(n7624), .C(n7707) );
  BUFFD0 U7624 ( .I(n7694), .Z(n7708) );
  CKBD0 U7625 ( .CLK(n7693), .C(n7709) );
  CKBD0 U7626 ( .CLK(n7695), .C(n7710) );
  CKBD0 U7627 ( .CLK(n7696), .C(n7711) );
  CKBD0 U7628 ( .CLK(n7697), .C(n7712) );
  CKBD0 U7629 ( .CLK(n7698), .C(n7713) );
  CKBD0 U7630 ( .CLK(n7699), .C(n7714) );
  CKBD0 U7631 ( .CLK(n7625), .C(n7715) );
  CKBD0 U7632 ( .CLK(n7626), .C(n7716) );
  CKBD0 U7633 ( .CLK(n7706), .C(n7717) );
  CKBD0 U7634 ( .CLK(n7627), .C(n7718) );
  CKBD0 U7635 ( .CLK(n7629), .C(n7719) );
  CKBD0 U7636 ( .CLK(n7630), .C(n7720) );
  CKBD0 U7637 ( .CLK(n7631), .C(n7721) );
  CKBD0 U7638 ( .CLK(n7709), .C(n7722) );
  CKBD0 U7639 ( .CLK(n7708), .C(n7723) );
  CKBD0 U7640 ( .CLK(n7710), .C(n7724) );
  CKBD0 U7641 ( .CLK(n7711), .C(n7725) );
  CKBD0 U7642 ( .CLK(n7635), .C(n7726) );
  CKBD0 U7643 ( .CLK(n7636), .C(n7727) );
  CKBD0 U7644 ( .CLK(n7712), .C(n7728) );
  CKBD0 U7645 ( .CLK(n7637), .C(n7729) );
  CKBD0 U7646 ( .CLK(n7646), .C(n7730) );
  CKBD0 U7647 ( .CLK(n7647), .C(n7731) );
  CKBD0 U7648 ( .CLK(n7648), .C(n7732) );
  CKBD0 U7649 ( .CLK(n7713), .C(n7733) );
  CKBD0 U7650 ( .CLK(n7714), .C(n7734) );
  CKBD0 U7651 ( .CLK(n7717), .C(n7735) );
  BUFFD0 U7652 ( .I(n7722), .Z(n7736) );
  CKBD0 U7653 ( .CLK(n7723), .C(n7737) );
  CKBD0 U7654 ( .CLK(n7724), .C(n7738) );
  CKBD0 U7655 ( .CLK(n7725), .C(n7739) );
  CKBD0 U7656 ( .CLK(n7649), .C(n7740) );
  CKBD0 U7657 ( .CLK(n7728), .C(n7741) );
  CKBD0 U7658 ( .CLK(n7650), .C(n7742) );
  CKBD0 U7659 ( .CLK(n7660), .C(n7743) );
  BUFFD0 U7660 ( .I(n7659), .Z(n7744) );
  CKBD0 U7661 ( .CLK(n7692), .C(n7745) );
  CKBD0 U7662 ( .CLK(n7700), .C(n7746) );
  CKBD0 U7663 ( .CLK(n7733), .C(n7747) );
  CKBD0 U7664 ( .CLK(n7701), .C(n7748) );
  CKBD0 U7665 ( .CLK(n7702), .C(n7749) );
  CKBD0 U7666 ( .CLK(n7704), .C(n7750) );
  CKBD0 U7667 ( .CLK(n7703), .C(n7751) );
  CKBD0 U7668 ( .CLK(n7705), .C(n7752) );
  BUFFD0 U7669 ( .I(n7707), .Z(n7753) );
  CKBD0 U7670 ( .CLK(n7715), .C(n7754) );
  CKBD0 U7671 ( .CLK(n7716), .C(n7755) );
  CKBD0 U7672 ( .CLK(n7734), .C(n7756) );
  CKBD0 U7673 ( .CLK(n7718), .C(n7757) );
  CKBD0 U7674 ( .CLK(n7719), .C(n7758) );
  CKBD0 U7675 ( .CLK(n7735), .C(n7759) );
  CKBD0 U7676 ( .CLK(n7720), .C(n7760) );
  CKBD0 U7677 ( .CLK(n7721), .C(n7761) );
  CKBD0 U7678 ( .CLK(n7736), .C(n7762) );
  CKBD0 U7679 ( .CLK(n7737), .C(n7763) );
  CKBD0 U7680 ( .CLK(n7738), .C(n7764) );
  CKBD0 U7681 ( .CLK(n7726), .C(n7765) );
  CKBD0 U7682 ( .CLK(n7739), .C(n7766) );
  CKBD0 U7683 ( .CLK(n7727), .C(n7767) );
  CKBD0 U7684 ( .CLK(n7729), .C(n7768) );
  CKBD0 U7685 ( .CLK(n7730), .C(n7769) );
  CKBD0 U7686 ( .CLK(n7731), .C(n7770) );
  CKBD0 U7687 ( .CLK(n7732), .C(n7771) );
  CKBD0 U7688 ( .CLK(n7741), .C(n7772) );
  CKBD0 U7689 ( .CLK(n7740), .C(n7773) );
  CKBD0 U7690 ( .CLK(n7742), .C(n7774) );
  CKBD0 U7691 ( .CLK(n7743), .C(n7775) );
  CKBD0 U7692 ( .CLK(n7744), .C(n7776) );
  CKBD0 U7693 ( .CLK(n7745), .C(n7777) );
  CKBD0 U7694 ( .CLK(n7746), .C(n7778) );
  CKBD0 U7695 ( .CLK(n7747), .C(n7779) );
  CKBD0 U7696 ( .CLK(n7748), .C(n7780) );
  CKBD0 U7697 ( .CLK(n7749), .C(n7781) );
  BUFFD0 U7698 ( .I(n7750), .Z(n7782) );
  CKBD0 U7699 ( .CLK(n7751), .C(n7783) );
  CKBD0 U7700 ( .CLK(n7752), .C(n7784) );
  CKBD0 U7701 ( .CLK(n7753), .C(n7785) );
  CKBD0 U7702 ( .CLK(n7756), .C(n7786) );
  CKBD0 U7703 ( .CLK(n7759), .C(n7787) );
  CKBD0 U7704 ( .CLK(n7762), .C(n7788) );
  CKBD0 U7705 ( .CLK(n7763), .C(n7789) );
  CKBD0 U7706 ( .CLK(n7764), .C(n7790) );
  CKBD0 U7707 ( .CLK(n7766), .C(n7791) );
  BUFFD0 U7708 ( .I(n7772), .Z(n7792) );
  CKBD0 U7709 ( .CLK(n7779), .C(n7793) );
  CKBD0 U7710 ( .CLK(n7754), .C(n7794) );
  CKBD0 U7711 ( .CLK(n7755), .C(n7795) );
  BUFFD0 U7712 ( .I(n7786), .Z(n7796) );
  CKBD0 U7713 ( .CLK(n7757), .C(n7797) );
  CKBD0 U7714 ( .CLK(n7758), .C(n7798) );
  CKBD0 U7715 ( .CLK(n7787), .C(n7799) );
  CKBD0 U7716 ( .CLK(n7788), .C(n7800) );
  CKBD0 U7717 ( .CLK(n7789), .C(n7801) );
  CKBD0 U7718 ( .CLK(n7790), .C(n7802) );
  CKBD0 U7719 ( .CLK(n7791), .C(n7803) );
  CKBD0 U7720 ( .CLK(n7792), .C(n7804) );
  BUFFD0 U7721 ( .I(n7793), .Z(n7805) );
  CKBD0 U7722 ( .CLK(n7796), .C(n7806) );
  CKBD0 U7723 ( .CLK(n7760), .C(n7807) );
  CKBD0 U7724 ( .CLK(n7761), .C(n7808) );
  CKBD0 U7725 ( .CLK(n7799), .C(n7809) );
  CKBD0 U7726 ( .CLK(n7800), .C(n7810) );
  CKBD0 U7727 ( .CLK(n7765), .C(n7811) );
  CKBD0 U7728 ( .CLK(n7767), .C(n7812) );
  BUFFD0 U7729 ( .I(n7802), .Z(n7813) );
  CKBD0 U7730 ( .CLK(n7801), .C(n7814) );
  CKBD0 U7731 ( .CLK(n7768), .C(n7815) );
  CKBD0 U7732 ( .CLK(n7771), .C(n7816) );
  CKBD0 U7733 ( .CLK(n7769), .C(n7817) );
  CKBD0 U7734 ( .CLK(n7770), .C(n7818) );
  BUFFD0 U7735 ( .I(n7803), .Z(n7819) );
  CKBD0 U7736 ( .CLK(n7773), .C(n7820) );
  CKBD0 U7737 ( .CLK(n7774), .C(n7821) );
  CKBD0 U7738 ( .CLK(n7775), .C(n7822) );
  CKBD0 U7739 ( .CLK(n7776), .C(n7823) );
  CKBD0 U7740 ( .CLK(n7777), .C(n7824) );
  CKBD0 U7741 ( .CLK(n7778), .C(n7825) );
  CKBD0 U7742 ( .CLK(n7780), .C(n7826) );
  CKBD0 U7743 ( .CLK(n7804), .C(n7827) );
  CKBD0 U7744 ( .CLK(n7781), .C(n7828) );
  CKBD0 U7745 ( .CLK(n7782), .C(n7829) );
  CKBD0 U7746 ( .CLK(n7783), .C(n7830) );
  CKBD0 U7747 ( .CLK(n7784), .C(n7831) );
  CKBD0 U7748 ( .CLK(n7794), .C(n7832) );
  CKBD0 U7749 ( .CLK(n7785), .C(n7833) );
  CKBD0 U7750 ( .CLK(n7805), .C(n7834) );
  CKBD0 U7751 ( .CLK(n7795), .C(n7835) );
  CKBD0 U7752 ( .CLK(n7797), .C(n7836) );
  CKBD0 U7753 ( .CLK(n7798), .C(n7837) );
  CKBD0 U7754 ( .CLK(n7806), .C(n7838) );
  CKBD0 U7755 ( .CLK(n7807), .C(n7839) );
  CKBD0 U7756 ( .CLK(n7808), .C(n7840) );
  CKBD0 U7757 ( .CLK(n7809), .C(n7841) );
  CKBD0 U7758 ( .CLK(n7810), .C(n7842) );
  CKBD0 U7759 ( .CLK(n7811), .C(n7843) );
  BUFFD0 U7760 ( .I(n7812), .Z(n7844) );
  CKBD0 U7761 ( .CLK(n7813), .C(n7845) );
  CKBD0 U7762 ( .CLK(n7815), .C(n7846) );
  CKBD0 U7763 ( .CLK(n7814), .C(n7847) );
  CKBD0 U7764 ( .CLK(n7819), .C(n7848) );
  CKBD0 U7765 ( .CLK(n7827), .C(n7849) );
  CKBD0 U7766 ( .CLK(n7834), .C(n7850) );
  CKBD0 U7767 ( .CLK(n7838), .C(n7851) );
  BUFFD0 U7768 ( .I(n7841), .Z(n7852) );
  CKBD0 U7769 ( .CLK(n7842), .C(n7853) );
  CKBD0 U7770 ( .CLK(n7817), .C(n7854) );
  BUFFD0 U7771 ( .I(n7816), .Z(n7855) );
  CKBD0 U7772 ( .CLK(n7818), .C(n7856) );
  CKBD0 U7773 ( .CLK(n7820), .C(n7857) );
  CKBD0 U7774 ( .CLK(n7821), .C(n7858) );
  CKBD0 U7775 ( .CLK(n7845), .C(n7859) );
  CKBD0 U7776 ( .CLK(n7847), .C(n7860) );
  CKBD0 U7777 ( .CLK(n7848), .C(n7861) );
  CKBD0 U7778 ( .CLK(n7849), .C(n7862) );
  CKBD0 U7779 ( .CLK(n7850), .C(n7863) );
  CKBD0 U7780 ( .CLK(n7851), .C(n7864) );
  CKBD0 U7781 ( .CLK(n7852), .C(n7865) );
  CKBD0 U7782 ( .CLK(n7853), .C(n7866) );
  CKBD0 U7783 ( .CLK(n7822), .C(n7867) );
  CKBD0 U7784 ( .CLK(n7823), .C(n7868) );
  CKBD0 U7785 ( .CLK(n7824), .C(n7869) );
  CKBD0 U7786 ( .CLK(n7826), .C(n7870) );
  CKBD0 U7787 ( .CLK(n7825), .C(n7871) );
  CKBD0 U7788 ( .CLK(n7860), .C(n7872) );
  CKBD0 U7789 ( .CLK(n7859), .C(n7873) );
  CKBD0 U7790 ( .CLK(n7828), .C(n7874) );
  CKBD0 U7791 ( .CLK(n7861), .C(n7875) );
  CKBD0 U7792 ( .CLK(n7862), .C(n7876) );
  CKBD0 U7793 ( .CLK(n7863), .C(n7877) );
  CKBD0 U7794 ( .CLK(n7864), .C(n7878) );
  CKBD0 U7795 ( .CLK(n7865), .C(n7879) );
  BUFFD0 U7796 ( .I(n7872), .Z(n7880) );
  CKBD0 U7797 ( .CLK(n7829), .C(n7881) );
  CKBD0 U7798 ( .CLK(n7830), .C(n7882) );
  CKBD0 U7799 ( .CLK(n7866), .C(n7883) );
  CKBD0 U7800 ( .CLK(n7831), .C(n7884) );
  CKBD0 U7801 ( .CLK(n7833), .C(n7885) );
  BUFFD0 U7802 ( .I(n7832), .Z(n7886) );
  CKBD0 U7803 ( .CLK(n7873), .C(n7887) );
  CKBD0 U7804 ( .CLK(n7875), .C(n7888) );
  CKBD0 U7805 ( .CLK(n7876), .C(n7889) );
  CKBD0 U7806 ( .CLK(n7877), .C(n7890) );
  CKBD0 U7807 ( .CLK(n7878), .C(n7891) );
  CKBD0 U7808 ( .CLK(n7879), .C(n7892) );
  CKBD0 U7809 ( .CLK(n7880), .C(n7893) );
  CKBD0 U7810 ( .CLK(n7883), .C(n7894) );
  BUFFD0 U7811 ( .I(n7836), .Z(n7895) );
  CKBD0 U7812 ( .CLK(n7835), .C(n7896) );
  CKBD0 U7813 ( .CLK(n7887), .C(n7897) );
  CKBD0 U7814 ( .CLK(n7888), .C(n7898) );
  CKBD0 U7815 ( .CLK(n7889), .C(n7899) );
  CKBD0 U7816 ( .CLK(n7890), .C(n7900) );
  CKBD0 U7817 ( .CLK(n7891), .C(n7901) );
  CKBD0 U7818 ( .CLK(n7892), .C(n7902) );
  CKBD0 U7819 ( .CLK(n7893), .C(n7903) );
  CKBD0 U7820 ( .CLK(n7894), .C(n7904) );
  CKBD0 U7821 ( .CLK(n7837), .C(n7905) );
  CKBD0 U7822 ( .CLK(n7839), .C(n7906) );
  CKBD0 U7823 ( .CLK(n7897), .C(n7907) );
  BUFFD0 U7824 ( .I(n7840), .Z(n7908) );
  CKBD0 U7825 ( .CLK(n7898), .C(n7909) );
  CKBD0 U7826 ( .CLK(n7899), .C(n7910) );
  CKBD0 U7827 ( .CLK(n7900), .C(n7911) );
  CKBD0 U7828 ( .CLK(n7843), .C(n7912) );
  CKBD0 U7829 ( .CLK(n7901), .C(n7913) );
  CKBD0 U7830 ( .CLK(n7844), .C(n7914) );
  CKBD0 U7831 ( .CLK(n7846), .C(n7915) );
  BUFFD0 U7832 ( .I(n7854), .Z(n7916) );
  CKBD0 U7833 ( .CLK(n7856), .C(n7917) );
  CKBD0 U7834 ( .CLK(n7855), .C(n7918) );
  CKBD0 U7835 ( .CLK(n7902), .C(n7919) );
  CKBD0 U7836 ( .CLK(n7904), .C(n7920) );
  CKBD0 U7837 ( .CLK(n7903), .C(n7921) );
  CKBD0 U7838 ( .CLK(n7907), .C(n7922) );
  CKBD0 U7839 ( .CLK(n7909), .C(n7923) );
  CKBD0 U7840 ( .CLK(n7910), .C(n7924) );
  CKBD0 U7841 ( .CLK(n7911), .C(n7925) );
  CKBD0 U7842 ( .CLK(n7913), .C(n7926) );
  CKBD0 U7843 ( .CLK(n7857), .C(n7927) );
  BUFFD0 U7844 ( .I(n7858), .Z(n7928) );
  CKBD0 U7845 ( .CLK(n7919), .C(n7929) );
  BUFFD0 U7846 ( .I(n7920), .Z(n7930) );
  CKBD0 U7847 ( .CLK(n7921), .C(n7931) );
  CKBD0 U7848 ( .CLK(n7922), .C(n7932) );
  CKBD0 U7849 ( .CLK(n7923), .C(n7933) );
  BUFFD0 U7850 ( .I(n7924), .Z(n7934) );
  CKBD0 U7851 ( .CLK(n7925), .C(n7935) );
  CKBD0 U7852 ( .CLK(n7926), .C(n7936) );
  CKBD0 U7853 ( .CLK(n7867), .C(n7937) );
  CKBD0 U7854 ( .CLK(n7868), .C(n7938) );
  CKBD0 U7855 ( .CLK(n7871), .C(n7939) );
  CKBD0 U7856 ( .CLK(n7869), .C(n7940) );
  BUFFD0 U7857 ( .I(n7870), .Z(n7941) );
  CKBD0 U7858 ( .CLK(n7874), .C(n7942) );
  CKBD0 U7859 ( .CLK(n7882), .C(n7943) );
  CKBD0 U7860 ( .CLK(n7881), .C(n7944) );
  CKBD0 U7861 ( .CLK(n7929), .C(n7945) );
  CKBD0 U7862 ( .CLK(n7884), .C(n7946) );
  CKBD0 U7863 ( .CLK(n7885), .C(n7947) );
  CKBD0 U7864 ( .CLK(n7886), .C(n7948) );
  CKBD0 U7865 ( .CLK(n7896), .C(n7949) );
  CKBD0 U7866 ( .CLK(n7895), .C(n7950) );
  CKBD0 U7867 ( .CLK(n7930), .C(n7951) );
  CKBD0 U7868 ( .CLK(n7931), .C(n7952) );
  CKBD0 U7869 ( .CLK(n7932), .C(n7953) );
  CKBD0 U7870 ( .CLK(n7933), .C(n7954) );
  CKBD0 U7871 ( .CLK(n7934), .C(n7955) );
  CKBD0 U7872 ( .CLK(n7935), .C(n7956) );
  BUFFD0 U7873 ( .I(n7936), .Z(n7957) );
  CKBD0 U7874 ( .CLK(n7945), .C(n7958) );
  BUFFD0 U7875 ( .I(n7906), .Z(n7959) );
  CKBD0 U7876 ( .CLK(n7905), .C(n7960) );
  CKBD0 U7877 ( .CLK(n7951), .C(n7961) );
  BUFFD0 U7878 ( .I(n7953), .Z(n7962) );
  CKBD0 U7879 ( .CLK(n7952), .C(n7963) );
  CKBD0 U7880 ( .CLK(n7954), .C(n7964) );
  CKBD0 U7881 ( .CLK(n7955), .C(n7965) );
  CKBD0 U7882 ( .CLK(n7956), .C(n7966) );
  CKBD0 U7883 ( .CLK(n7957), .C(n7967) );
  CKBD0 U7884 ( .CLK(n7958), .C(n7968) );
  CKBD0 U7885 ( .CLK(n7908), .C(n7969) );
  CKBD0 U7886 ( .CLK(n7961), .C(n7970) );
  CKBD0 U7887 ( .CLK(n7962), .C(n7971) );
  CKBD0 U7888 ( .CLK(n7963), .C(n7972) );
  BUFFD0 U7889 ( .I(n7964), .Z(n7973) );
  CKBD0 U7890 ( .CLK(n7912), .C(n7974) );
  CKBD0 U7891 ( .CLK(n7914), .C(n7975) );
  CKBD0 U7892 ( .CLK(n7965), .C(n7976) );
  BUFFD0 U7893 ( .I(n7915), .Z(n7977) );
  CKBD0 U7894 ( .CLK(n7916), .C(n7978) );
  BUFFD0 U7895 ( .I(n7917), .Z(n7979) );
  CKBD0 U7896 ( .CLK(n7918), .C(n7980) );
  BUFFD0 U7897 ( .I(n7927), .Z(n7981) );
  CKBD0 U7898 ( .CLK(n7928), .C(n7982) );
  CKBD0 U7899 ( .CLK(n7966), .C(n7983) );
  CKBD0 U7900 ( .CLK(n7937), .C(n7984) );
  CKBD0 U7901 ( .CLK(n7938), .C(n7985) );
  CKBD0 U7902 ( .CLK(n7940), .C(n7986) );
  BUFFD0 U7903 ( .I(n7939), .Z(n7987) );
  CKBD0 U7904 ( .CLK(n7967), .C(n7988) );
  CKBD0 U7905 ( .CLK(n7968), .C(n7989) );
  CKBD0 U7906 ( .CLK(n7970), .C(n7990) );
  CKBD0 U7907 ( .CLK(n7971), .C(n7991) );
  CKBD0 U7908 ( .CLK(n7972), .C(n7992) );
  CKBD0 U7909 ( .CLK(n7973), .C(n7993) );
  CKBD0 U7910 ( .CLK(n7976), .C(n7994) );
  BUFFD0 U7911 ( .I(n7983), .Z(n7995) );
  CKBD0 U7912 ( .CLK(n7941), .C(n7996) );
  CKBD0 U7913 ( .CLK(n7988), .C(n7997) );
  BUFFD0 U7914 ( .I(n7989), .Z(n7998) );
  CKBD0 U7915 ( .CLK(n7990), .C(n7999) );
  CKBD0 U7916 ( .CLK(n7992), .C(n8000) );
  CKBD0 U7917 ( .CLK(n7991), .C(n8001) );
  CKBD0 U7918 ( .CLK(n7993), .C(n8002) );
  CKBD0 U7919 ( .CLK(n7994), .C(n8003) );
  BUFFD0 U7920 ( .I(n7942), .Z(n8004) );
  BUFFD0 U7921 ( .I(n7943), .Z(n8005) );
  CKBD0 U7922 ( .CLK(n7944), .C(n8006) );
  CKBD0 U7923 ( .CLK(n7946), .C(n8007) );
  CKBD0 U7924 ( .CLK(n7947), .C(n8008) );
  CKBD0 U7925 ( .CLK(n7995), .C(n8009) );
  CKBD0 U7926 ( .CLK(n7948), .C(n8010) );
  BUFFD0 U7927 ( .I(n7949), .Z(n8011) );
  CKBD0 U7928 ( .CLK(n7950), .C(n8012) );
  BUFFD0 U7929 ( .I(n7960), .Z(n8013) );
  CKBD0 U7930 ( .CLK(n7959), .C(n8014) );
  CKBD0 U7931 ( .CLK(n7997), .C(n8015) );
  CKBD0 U7932 ( .CLK(n7969), .C(n8016) );
  CKBD0 U7933 ( .CLK(n7998), .C(n8017) );
  BUFFD0 U7934 ( .I(n8000), .Z(n8018) );
  CKBD0 U7935 ( .CLK(n7999), .C(n8019) );
  CKBD0 U7936 ( .CLK(n7974), .C(n8020) );
  CKBD0 U7937 ( .CLK(n8001), .C(n8021) );
  CKBD0 U7938 ( .CLK(n7975), .C(n8022) );
  CKBD0 U7939 ( .CLK(n8002), .C(n8023) );
  CKBD0 U7940 ( .CLK(n8003), .C(n8024) );
  CKBD0 U7941 ( .CLK(n8009), .C(n8025) );
  CKBD0 U7942 ( .CLK(n8015), .C(n8026) );
  CKBD0 U7943 ( .CLK(n8017), .C(n8027) );
  CKBD0 U7944 ( .CLK(n8018), .C(n8028) );
  CKBD0 U7945 ( .CLK(n7977), .C(n8029) );
  CKBD0 U7946 ( .CLK(n8019), .C(n8030) );
  CKBD0 U7947 ( .CLK(n7978), .C(n8031) );
  CKBD0 U7948 ( .CLK(n7979), .C(n8032) );
  CKBD0 U7949 ( .CLK(n7980), .C(n8033) );
  CKBD0 U7950 ( .CLK(n7981), .C(n8034) );
  CKBD0 U7951 ( .CLK(n8021), .C(n8035) );
  CKBD0 U7952 ( .CLK(n8023), .C(n8036) );
  CKBD0 U7953 ( .CLK(n8024), .C(n8037) );
  CKBD0 U7954 ( .CLK(n8025), .C(n8038) );
  CKBD0 U7955 ( .CLK(n8026), .C(n8039) );
  CKBD0 U7956 ( .CLK(n8027), .C(n8040) );
  CKBD0 U7957 ( .CLK(n8030), .C(n8041) );
  CKBD0 U7958 ( .CLK(n8028), .C(n8042) );
  CKBD0 U7959 ( .CLK(n8035), .C(n8043) );
  CKBD0 U7960 ( .CLK(n8036), .C(n8044) );
  CKBD0 U7961 ( .CLK(n8037), .C(n8045) );
  CKBD0 U7962 ( .CLK(n8038), .C(n8046) );
  CKBD0 U7963 ( .CLK(n8039), .C(n8047) );
  CKBD0 U7964 ( .CLK(n8040), .C(n8048) );
  BUFFD0 U7965 ( .I(n8041), .Z(n8049) );
  CKBD0 U7966 ( .CLK(n7982), .C(n8050) );
  CKBD0 U7967 ( .CLK(n7986), .C(n8051) );
  CKBD0 U7968 ( .CLK(n7984), .C(n8052) );
  CKBD0 U7969 ( .CLK(n7985), .C(n8053) );
  CKBD0 U7970 ( .CLK(n7987), .C(n8054) );
  CKBD0 U7971 ( .CLK(n7996), .C(n8055) );
  CKBD0 U7972 ( .CLK(n8042), .C(n8056) );
  CKBD0 U7973 ( .CLK(n8004), .C(n8057) );
  CKBD0 U7974 ( .CLK(n8043), .C(n8058) );
  CKBD0 U7975 ( .CLK(n8044), .C(n8059) );
  CKBD0 U7976 ( .CLK(n8045), .C(n8060) );
  CKBD0 U7977 ( .CLK(n8046), .C(n8061) );
  CKBD0 U7978 ( .CLK(n8047), .C(n8062) );
  CKBD0 U7979 ( .CLK(n8048), .C(n8063) );
  CKBD0 U7980 ( .CLK(n8049), .C(n8064) );
  CKBD0 U7981 ( .CLK(n8005), .C(n8065) );
  CKBD0 U7982 ( .CLK(n8006), .C(n8066) );
  CKBD0 U7983 ( .CLK(n8007), .C(n8067) );
  CKBD0 U7984 ( .CLK(n8008), .C(n8068) );
  CKBD0 U7985 ( .CLK(n8010), .C(n8069) );
  CKBD0 U7986 ( .CLK(n8056), .C(n8070) );
  CKBD0 U7987 ( .CLK(n8058), .C(n8071) );
  CKBD0 U7988 ( .CLK(n8059), .C(n8072) );
  CKBD0 U7989 ( .CLK(n8060), .C(n8073) );
  CKBD0 U7990 ( .CLK(n8061), .C(n8074) );
  CKBD0 U7991 ( .CLK(n8062), .C(n8075) );
  CKBD0 U7992 ( .CLK(n8063), .C(n8076) );
  CKBD0 U7993 ( .CLK(n8064), .C(n8077) );
  CKBD0 U7994 ( .CLK(n8011), .C(n8078) );
  CKBD0 U7995 ( .CLK(n8012), .C(n8079) );
  CKBD0 U7996 ( .CLK(n8013), .C(n8080) );
  CKBD0 U7997 ( .CLK(n8070), .C(n8081) );
  CKBD0 U7998 ( .CLK(n8014), .C(n8082) );
  CKBD0 U7999 ( .CLK(n8071), .C(n8083) );
  CKBD0 U8000 ( .CLK(n8016), .C(n8084) );
  CKBD0 U8001 ( .CLK(n8072), .C(n8085) );
  BUFFD0 U8002 ( .I(n8073), .Z(n8086) );
  CKBD0 U8003 ( .CLK(n8074), .C(n8087) );
  CKBD0 U8004 ( .CLK(n8075), .C(n8088) );
  CKBD0 U8005 ( .CLK(n8020), .C(n8089) );
  CKBD0 U8006 ( .CLK(n8022), .C(n8090) );
  CKBD0 U8007 ( .CLK(n8029), .C(n8091) );
  CKBD0 U8008 ( .CLK(n8076), .C(n8092) );
  CKBD0 U8009 ( .CLK(n8077), .C(n8093) );
  CKBD0 U8010 ( .CLK(n8081), .C(n8094) );
  CKBD0 U8011 ( .CLK(n8083), .C(n8095) );
  CKBD0 U8012 ( .CLK(n8085), .C(n8096) );
  CKBD0 U8013 ( .CLK(n8086), .C(n8097) );
  CKBD0 U8014 ( .CLK(n8087), .C(n8098) );
  CKBD0 U8015 ( .CLK(n8088), .C(n8099) );
  CKBD0 U8016 ( .CLK(n8031), .C(n8100) );
  CKBD0 U8017 ( .CLK(n8032), .C(n8101) );
  CKBD0 U8018 ( .CLK(n8033), .C(n8102) );
  CKBD0 U8019 ( .CLK(n8034), .C(n8103) );
  CKBD0 U8020 ( .CLK(n8050), .C(n8104) );
  CKBD0 U8021 ( .CLK(n8092), .C(n8105) );
  CKBD0 U8022 ( .CLK(n8052), .C(n8106) );
  BUFFD0 U8023 ( .I(n8051), .Z(n8107) );
  CKBD0 U8024 ( .CLK(n8053), .C(n8108) );
  CKBD0 U8025 ( .CLK(n8054), .C(n8109) );
  CKBD0 U8026 ( .CLK(n8055), .C(n8110) );
  CKBD0 U8027 ( .CLK(n8057), .C(n8111) );
  CKBD0 U8028 ( .CLK(n8066), .C(n8112) );
  CKBD0 U8029 ( .CLK(n8065), .C(n8113) );
  CKBD0 U8030 ( .CLK(n8093), .C(n8114) );
  CKBD0 U8031 ( .CLK(n8094), .C(n8115) );
  CKBD0 U8032 ( .CLK(n8095), .C(n8116) );
  CKBD0 U8033 ( .CLK(n8096), .C(n8117) );
  CKBD0 U8034 ( .CLK(n8097), .C(n8118) );
  BUFFD0 U8035 ( .I(n8098), .Z(n8119) );
  BUFFD0 U8036 ( .I(n8099), .Z(n8120) );
  CKBD0 U8037 ( .CLK(n8105), .C(n8121) );
  CKBD0 U8038 ( .CLK(n8068), .C(n8122) );
  CKBD0 U8039 ( .CLK(n8067), .C(n8123) );
  CKBD0 U8040 ( .CLK(n8069), .C(n8124) );
  CKBD0 U8041 ( .CLK(n8114), .C(n8125) );
  BUFFD0 U8042 ( .I(n8116), .Z(n8126) );
  CKBD0 U8043 ( .CLK(n8115), .C(n8127) );
  BUFFD0 U8044 ( .I(n8117), .Z(n8128) );
  CKBD0 U8045 ( .CLK(n8118), .C(n8129) );
  CKBD0 U8046 ( .CLK(n8119), .C(n8130) );
  CKBD0 U8047 ( .CLK(n8120), .C(n8131) );
  CKBD0 U8048 ( .CLK(n8121), .C(n8132) );
  CKBD0 U8049 ( .CLK(n8078), .C(n8133) );
  CKBD0 U8050 ( .CLK(n8079), .C(n8134) );
  CKBD0 U8051 ( .CLK(n8080), .C(n8135) );
  CKBD0 U8052 ( .CLK(n8125), .C(n8136) );
  CKBD0 U8053 ( .CLK(n8126), .C(n8137) );
  CKBD0 U8054 ( .CLK(n8127), .C(n8138) );
  CKBD0 U8055 ( .CLK(n8128), .C(n8139) );
  CKBD0 U8056 ( .CLK(n8129), .C(n8140) );
  CKBD0 U8057 ( .CLK(n8130), .C(n8141) );
  CKBD0 U8058 ( .CLK(n8131), .C(n8142) );
  CKBD0 U8059 ( .CLK(n8132), .C(n8143) );
  CKBD0 U8060 ( .CLK(n8082), .C(n8144) );
  CKBD0 U8061 ( .CLK(n8084), .C(n8145) );
  CKBD0 U8062 ( .CLK(n8136), .C(n8146) );
  CKBD0 U8063 ( .CLK(n8138), .C(n8147) );
  CKBD0 U8064 ( .CLK(n8137), .C(n8148) );
  CKBD0 U8065 ( .CLK(n8139), .C(n8149) );
  CKBD0 U8066 ( .CLK(n8089), .C(n8150) );
  CKBD0 U8067 ( .CLK(n8140), .C(n8151) );
  CKBD0 U8068 ( .CLK(n8090), .C(n8152) );
  CKBD0 U8069 ( .CLK(n8091), .C(n8153) );
  CKBD0 U8070 ( .CLK(n8100), .C(n8154) );
  CKBD0 U8071 ( .CLK(n8102), .C(n8155) );
  CKBD0 U8072 ( .CLK(n8141), .C(n8156) );
  CKBD0 U8073 ( .CLK(n8142), .C(n8157) );
  BUFFD0 U8074 ( .I(n8143), .Z(n8158) );
  BUFFD0 U8075 ( .I(n8147), .Z(n8159) );
  CKBD0 U8076 ( .CLK(n8146), .C(n8160) );
  CKBD0 U8077 ( .CLK(n8148), .C(n8161) );
  CKBD0 U8078 ( .CLK(n8149), .C(n8162) );
  CKBD0 U8079 ( .CLK(n8101), .C(n8163) );
  CKBD0 U8080 ( .CLK(n8151), .C(n8164) );
  CKBD0 U8081 ( .CLK(n8103), .C(n8165) );
  CKBD0 U8082 ( .CLK(n8104), .C(n8166) );
  BUFFD0 U8083 ( .I(n8106), .Z(n8167) );
  CKBD0 U8084 ( .CLK(n8156), .C(n8168) );
  CKBD0 U8085 ( .CLK(n8109), .C(n8169) );
  CKBD0 U8086 ( .CLK(n8107), .C(n8170) );
  CKBD0 U8087 ( .CLK(n8157), .C(n8171) );
  CKBD0 U8088 ( .CLK(n8158), .C(n8172) );
  CKBD0 U8089 ( .CLK(n8159), .C(n8173) );
  CKBD0 U8090 ( .CLK(n8160), .C(n8174) );
  CKBD0 U8091 ( .CLK(n8161), .C(n8175) );
  CKBD0 U8092 ( .CLK(n8162), .C(n8176) );
  CKBD0 U8093 ( .CLK(n8164), .C(n8177) );
  CKBD0 U8094 ( .CLK(n8108), .C(n8178) );
  CKBD0 U8095 ( .CLK(n8110), .C(n8179) );
  BUFFD0 U8096 ( .I(n8355), .Z(n8180) );
  CKBD0 U8097 ( .CLK(n8113), .C(n8181) );
  CKBD0 U8098 ( .CLK(n8111), .C(n8182) );
  CKBD0 U8099 ( .CLK(n8168), .C(n8183) );
  CKBD0 U8100 ( .CLK(n8124), .C(n8184) );
  CKBD0 U8101 ( .CLK(n8123), .C(n8185) );
  BUFFD0 U8102 ( .I(n8122), .Z(n8186) );
  CKBD0 U8103 ( .CLK(n8171), .C(n8187) );
  CKBD0 U8104 ( .CLK(n8172), .C(n8188) );
  CKBD0 U8105 ( .CLK(n8174), .C(n8189) );
  CKBD0 U8106 ( .CLK(n8173), .C(n8190) );
  CKBD0 U8107 ( .CLK(n8175), .C(n8191) );
  CKBD0 U8108 ( .CLK(n8176), .C(n8192) );
  CKBD0 U8109 ( .CLK(n8177), .C(n8193) );
  CKBD0 U8110 ( .CLK(n8133), .C(n8194) );
  CKBD0 U8111 ( .CLK(n8183), .C(n8195) );
  CKBD0 U8112 ( .CLK(n8134), .C(n8196) );
  CKBD0 U8113 ( .CLK(n8135), .C(n8197) );
  CKBD0 U8114 ( .CLK(n8144), .C(n8198) );
  CKBD0 U8115 ( .CLK(n8187), .C(n8199) );
  CKBD0 U8116 ( .CLK(n8145), .C(n8200) );
  CKBD0 U8117 ( .CLK(n8188), .C(n8201) );
  BUFFD0 U8118 ( .I(n8189), .Z(n8202) );
  BUFFD0 U8119 ( .I(n8150), .Z(n8203) );
  CKBD0 U8120 ( .CLK(n8190), .C(n8204) );
  BUFFD0 U8121 ( .I(n8152), .Z(n8205) );
  CKBD0 U8122 ( .CLK(n8191), .C(n8206) );
  CKBD0 U8123 ( .CLK(n8192), .C(n8207) );
  CKBD0 U8124 ( .CLK(n8193), .C(n8208) );
  CKBD0 U8125 ( .CLK(n8195), .C(n8209) );
  CKBD0 U8126 ( .CLK(n8199), .C(n8210) );
  CKBD0 U8127 ( .CLK(n8201), .C(n8211) );
  CKBD0 U8128 ( .CLK(n8202), .C(n8212) );
  CKBD0 U8129 ( .CLK(n8153), .C(n8213) );
  BUFFD0 U8130 ( .I(n8276), .Z(n8214) );
  BUFFD0 U8131 ( .I(n8277), .Z(n8215) );
  CKBD0 U8132 ( .CLK(n8163), .C(n8216) );
  CKBD0 U8133 ( .CLK(n8165), .C(n8217) );
  CKBD0 U8134 ( .CLK(n8204), .C(n8218) );
  BUFFD0 U8135 ( .I(n8166), .Z(n8219) );
  CKBD0 U8136 ( .CLK(n8178), .C(n8220) );
  CKBD0 U8137 ( .CLK(n8167), .C(n8221) );
  CKBD0 U8138 ( .CLK(n8170), .C(n8222) );
  CKBD0 U8139 ( .CLK(n8206), .C(n8223) );
  BUFFD0 U8140 ( .I(n8169), .Z(n8224) );
  CKBD0 U8141 ( .CLK(n8207), .C(n8225) );
  CKBD0 U8142 ( .CLK(n8208), .C(n8226) );
  CKBD0 U8143 ( .CLK(n8209), .C(n8227) );
  CKBD0 U8144 ( .CLK(n8210), .C(n8228) );
  CKBD0 U8145 ( .CLK(n8211), .C(n8229) );
  CKBD0 U8146 ( .CLK(n8212), .C(n8230) );
  CKBD0 U8147 ( .CLK(n8218), .C(n8231) );
  BUFFD0 U8148 ( .I(n8179), .Z(n8232) );
  CKBD0 U8149 ( .CLK(n8223), .C(n8233) );
  CKBD0 U8150 ( .CLK(n8225), .C(n8234) );
  BUFFD0 U8151 ( .I(n8226), .Z(n8235) );
  CKBD0 U8152 ( .CLK(n8227), .C(n8236) );
  CKBD0 U8153 ( .CLK(n8228), .C(n8237) );
  CKBD0 U8154 ( .CLK(n8229), .C(n8238) );
  CKBD0 U8155 ( .CLK(n8230), .C(n8239) );
  CKBD0 U8156 ( .CLK(n8182), .C(n8240) );
  BUFFD0 U8157 ( .I(n8112), .Z(n8241) );
  BUFFD0 U8158 ( .I(n8181), .Z(n8242) );
  CKBD0 U8159 ( .CLK(n8185), .C(n8243) );
  CKBD0 U8160 ( .CLK(n8186), .C(n8244) );
  BUFFD0 U8161 ( .I(n8184), .Z(n8245) );
  CKBD0 U8162 ( .CLK(n8231), .C(n8246) );
  CKBD0 U8163 ( .CLK(n8233), .C(n8247) );
  BUFFD0 U8164 ( .I(n8234), .Z(n8248) );
  CKBD0 U8165 ( .CLK(n8235), .C(n8249) );
  BUFFD0 U8166 ( .I(n8236), .Z(n8250) );
  BUFFD0 U8167 ( .I(n8237), .Z(n8251) );
  CKBD0 U8168 ( .CLK(n8238), .C(n8252) );
  CKBD0 U8169 ( .CLK(n8239), .C(n8253) );
  BUFFD0 U8170 ( .I(n8316), .Z(n8254) );
  BUFFD0 U8171 ( .I(n8247), .Z(n8255) );
  CKBD0 U8172 ( .CLK(n8246), .C(n8256) );
  CKBD0 U8173 ( .CLK(n8196), .C(n8257) );
  CKBD0 U8174 ( .CLK(n8248), .C(n8258) );
  CKBD0 U8175 ( .CLK(n8249), .C(n8259) );
  CKBD0 U8176 ( .CLK(n8250), .C(n8260) );
  CKBD0 U8177 ( .CLK(n8251), .C(n8261) );
  CKBD0 U8178 ( .CLK(n8252), .C(n8262) );
  CKBD0 U8179 ( .CLK(n8253), .C(n8263) );
  CKBD0 U8180 ( .CLK(n8197), .C(n8264) );
  CKBD0 U8181 ( .CLK(n8198), .C(n8265) );
  CKBD0 U8182 ( .CLK(n8255), .C(n8266) );
  CKBD0 U8183 ( .CLK(n8256), .C(n8267) );
  CKBD0 U8184 ( .CLK(n8258), .C(n8268) );
  CKBD0 U8185 ( .CLK(n8200), .C(n8269) );
  CKBD0 U8186 ( .CLK(n8259), .C(n8270) );
  CKBD0 U8187 ( .CLK(n8260), .C(n8271) );
  CKBD0 U8188 ( .CLK(n8261), .C(n8272) );
  CKBD0 U8189 ( .CLK(n8203), .C(n8273) );
  CKBD0 U8190 ( .CLK(n8205), .C(n8274) );
  BUFFD0 U8191 ( .I(n8421), .Z(n8275) );
  BUFFD0 U8192 ( .I(n8335), .Z(n8276) );
  BUFFD0 U8193 ( .I(n8993), .Z(n8277) );
  CKBD0 U8194 ( .CLK(n8262), .C(n8278) );
  CKBD0 U8195 ( .CLK(n8263), .C(n8279) );
  CKBD0 U8196 ( .CLK(n8266), .C(n8280) );
  CKBD0 U8197 ( .CLK(n8267), .C(n8281) );
  CKBD0 U8198 ( .CLK(n8268), .C(n8282) );
  CKBD0 U8199 ( .CLK(n8270), .C(n8283) );
  CKBD0 U8200 ( .CLK(n8271), .C(n8284) );
  CKBD0 U8201 ( .CLK(n8272), .C(n8285) );
  BUFFD0 U8202 ( .I(n8432), .Z(n8286) );
  BUFFD0 U8203 ( .I(n8216), .Z(n8287) );
  CKBD0 U8204 ( .CLK(n8219), .C(n8288) );
  BUFFD0 U8205 ( .I(n8278), .Z(n8289) );
  CKBD0 U8206 ( .CLK(n8279), .C(n8290) );
  CKBD0 U8207 ( .CLK(n8281), .C(n8291) );
  CKBD0 U8208 ( .CLK(n8280), .C(n8292) );
  CKBD0 U8209 ( .CLK(n8282), .C(n8293) );
  CKBD0 U8210 ( .CLK(n8283), .C(n8294) );
  CKBD0 U8211 ( .CLK(n8284), .C(n8295) );
  CKBD0 U8212 ( .CLK(n8285), .C(n8296) );
  CKBD0 U8213 ( .CLK(n8221), .C(n8297) );
  CKBD0 U8214 ( .CLK(n8222), .C(n8298) );
  CKBD0 U8215 ( .CLK(n8224), .C(n8299) );
  BUFFD0 U8216 ( .I(n8220), .Z(n8300) );
  CKBD0 U8217 ( .CLK(n8232), .C(n8301) );
  CKBD0 U8218 ( .CLK(n8241), .C(n8302) );
  CKBD0 U8219 ( .CLK(n8242), .C(n8303) );
  BUFFD0 U8220 ( .I(n8240), .Z(n8304) );
  CKBD0 U8221 ( .CLK(n8289), .C(n8305) );
  BUFFD0 U8222 ( .I(n8291), .Z(n8306) );
  CKBD0 U8223 ( .CLK(n8290), .C(n8307) );
  CKBD0 U8224 ( .CLK(n8292), .C(n8308) );
  CKBD0 U8225 ( .CLK(n8293), .C(n8309) );
  CKBD0 U8226 ( .CLK(n8294), .C(n8310) );
  CKBD0 U8227 ( .CLK(n8295), .C(n8311) );
  CKBD0 U8228 ( .CLK(n8296), .C(n8312) );
  CKBD0 U8229 ( .CLK(n8245), .C(n8313) );
  BUFFD0 U8230 ( .I(n8243), .Z(n8314) );
  BUFFD0 U8231 ( .I(n8244), .Z(n8315) );
  BUFFD0 U8232 ( .I(n8495), .Z(n8316) );
  BUFFD0 U8233 ( .I(n8257), .Z(n8317) );
  CKBD0 U8234 ( .CLK(n8305), .C(n8318) );
  CKBD0 U8235 ( .CLK(n8307), .C(n8319) );
  CKBD0 U8236 ( .CLK(n8306), .C(n8320) );
  CKBD0 U8237 ( .CLK(n8308), .C(n8321) );
  CKBD0 U8238 ( .CLK(n8309), .C(n8322) );
  CKBD0 U8239 ( .CLK(n8310), .C(n8323) );
  CKBD0 U8240 ( .CLK(n8311), .C(n8324) );
  CKBD0 U8241 ( .CLK(n8312), .C(n8325) );
  BUFFD0 U8242 ( .I(n8265), .Z(n8326) );
  CKBD0 U8243 ( .CLK(n8264), .C(n8327) );
  CKBD0 U8244 ( .CLK(n8318), .C(n8328) );
  CKBD0 U8245 ( .CLK(n8269), .C(n8329) );
  BUFFD0 U8246 ( .I(n8319), .Z(n8330) );
  CKBD0 U8247 ( .CLK(n8320), .C(n8331) );
  CKBD0 U8248 ( .CLK(n8321), .C(n8332) );
  BUFFD0 U8249 ( .I(n8524), .Z(n8333) );
  CKBD0 U8250 ( .CLK(n8322), .C(n8334) );
  BUFFD0 U8251 ( .I(n8954), .Z(n8335) );
  BUFFD0 U8252 ( .I(n8274), .Z(n8336) );
  BUFFD0 U8253 ( .I(n8213), .Z(n8337) );
  BUFFD0 U8254 ( .I(n8155), .Z(n8338) );
  CKBD0 U8255 ( .CLK(n8287), .C(n8339) );
  CKBD0 U8256 ( .CLK(n8323), .C(n8340) );
  BUFFD0 U8257 ( .I(n8217), .Z(n8341) );
  BUFFD0 U8258 ( .I(n8678), .Z(n8342) );
  BUFFD0 U8259 ( .I(n8682), .Z(n8343) );
  CKBD0 U8260 ( .CLK(n8324), .C(n8344) );
  BUFFD0 U8261 ( .I(n8536), .Z(n8345) );
  CKBD0 U8262 ( .CLK(n8300), .C(n8346) );
  BUFFD0 U8263 ( .I(n8297), .Z(n8347) );
  CKBD0 U8264 ( .CLK(n8325), .C(n8348) );
  CKBD0 U8265 ( .CLK(n8328), .C(n8349) );
  CKBD0 U8266 ( .CLK(n8330), .C(n8350) );
  CKBD0 U8267 ( .CLK(n8331), .C(n8351) );
  CKBD0 U8268 ( .CLK(n8332), .C(n8352) );
  CKBD0 U8269 ( .CLK(n8334), .C(n8353) );
  CKBD0 U8270 ( .CLK(n8340), .C(n8354) );
  BUFFD0 U8271 ( .I(n8971), .Z(n8355) );
  BUFFD0 U8272 ( .I(n8299), .Z(n8356) );
  BUFFD0 U8273 ( .I(n8401), .Z(n8357) );
  CKBD0 U8274 ( .CLK(n8304), .C(n8358) );
  BUFFD0 U8275 ( .I(n8708), .Z(n8359) );
  CKBD0 U8276 ( .CLK(n8344), .C(n8360) );
  CKBD0 U8277 ( .CLK(n8314), .C(n8361) );
  CKBD0 U8278 ( .CLK(n8315), .C(n8362) );
  CKBD0 U8279 ( .CLK(n8348), .C(n8363) );
  CKBD0 U8280 ( .CLK(n8349), .C(n8364) );
  CKBD0 U8281 ( .CLK(n8350), .C(n8365) );
  CKBD0 U8282 ( .CLK(n8351), .C(n8366) );
  CKBD0 U8283 ( .CLK(n8352), .C(n8367) );
  CKBD0 U8284 ( .CLK(n8353), .C(n8368) );
  CKBD0 U8285 ( .CLK(n8354), .C(n8369) );
  CKBD0 U8286 ( .CLK(n8360), .C(n8370) );
  BUFFD0 U8287 ( .I(n8194), .Z(n8371) );
  CKBD0 U8288 ( .CLK(n8317), .C(n8372) );
  BUFFD0 U8289 ( .I(n8408), .Z(n8373) );
  CKBD0 U8290 ( .CLK(n8363), .C(n8374) );
  CKBD0 U8291 ( .CLK(n8364), .C(n8375) );
  CKBD0 U8292 ( .CLK(n8365), .C(n8376) );
  CKBD0 U8293 ( .CLK(n8366), .C(n8377) );
  CKBD0 U8294 ( .CLK(n8367), .C(n8378) );
  CKBD0 U8295 ( .CLK(n8368), .C(n8379) );
  BUFFD0 U8296 ( .I(n8369), .Z(n8380) );
  CKBD0 U8297 ( .CLK(n8370), .C(n8381) );
  CKBD0 U8298 ( .CLK(n8326), .C(n8382) );
  BUFFD0 U8299 ( .I(n8558), .Z(n8383) );
  CKBD0 U8300 ( .CLK(n8374), .C(n8384) );
  CKBD0 U8301 ( .CLK(n8375), .C(n8385) );
  CKBD0 U8302 ( .CLK(n8376), .C(n8386) );
  BUFFD0 U8303 ( .I(n8273), .Z(n8387) );
  CKBD0 U8304 ( .CLK(n8336), .C(n8388) );
  BUFFD0 U8305 ( .I(n8154), .Z(n8389) );
  CKBD0 U8306 ( .CLK(n8337), .C(n8390) );
  CKBD0 U8307 ( .CLK(n8338), .C(n8391) );
  CKBD0 U8308 ( .CLK(n8377), .C(n8392) );
  CKBD0 U8309 ( .CLK(n8341), .C(n8393) );
  BUFFD0 U8310 ( .I(n8339), .Z(n8394) );
  CKBD0 U8311 ( .CLK(n8378), .C(n8395) );
  BUFFD0 U8312 ( .I(n8288), .Z(n8396) );
  BUFFD0 U8313 ( .I(n8379), .Z(n8397) );
  BUFFD0 U8314 ( .I(n8588), .Z(n8398) );
  BUFFD0 U8315 ( .I(n8298), .Z(n8399) );
  CKBD0 U8316 ( .CLK(n8347), .C(n8400) );
  BUFFD0 U8317 ( .I(n8880), .Z(n8401) );
  BUFFD0 U8318 ( .I(n8301), .Z(n8402) );
  BUFFD0 U8319 ( .I(n8302), .Z(n8403) );
  CKBD0 U8320 ( .CLK(n8356), .C(n8404) );
  BUFFD0 U8321 ( .I(n8358), .Z(n8405) );
  CKBD0 U8322 ( .CLK(n8380), .C(n8406) );
  BUFFD0 U8323 ( .I(n8372), .Z(n8407) );
  BUFFD0 U8324 ( .I(n8447), .Z(n8408) );
  BUFFD0 U8325 ( .I(n8313), .Z(n8409) );
  BUFFD0 U8326 ( .I(n8361), .Z(n8410) );
  BUFFD0 U8327 ( .I(n8362), .Z(n8411) );
  CKBD0 U8328 ( .CLK(n8371), .C(n8412) );
  CKBD0 U8329 ( .CLK(n8381), .C(n8413) );
  CKBD0 U8330 ( .CLK(n8382), .C(n8414) );
  BUFFD0 U8331 ( .I(n8329), .Z(n8415) );
  BUFFD0 U8332 ( .I(n8384), .Z(n8416) );
  CKBD0 U8333 ( .CLK(n8385), .C(n8417) );
  CKBD0 U8334 ( .CLK(n8387), .C(n8418) );
  CKBD0 U8335 ( .CLK(n8386), .C(n8419) );
  BUFFD0 U8336 ( .I(n8808), .Z(n8420) );
  BUFFD0 U8337 ( .I(n8824), .Z(n8421) );
  CKBD0 U8338 ( .CLK(n8389), .C(n8422) );
  BUFFD0 U8339 ( .I(n8391), .Z(n8423) );
  BUFFD0 U8340 ( .I(n8395), .Z(n8424) );
  CKBD0 U8341 ( .CLK(n8392), .C(n8425) );
  CKBD0 U8342 ( .CLK(n8397), .C(n8426) );
  CKBD0 U8343 ( .CLK(n8406), .C(n8427) );
  CKBD0 U8344 ( .CLK(n8413), .C(n8428) );
  CKBD0 U8345 ( .CLK(n8416), .C(n8429) );
  CKBD0 U8346 ( .CLK(n8417), .C(n8430) );
  CKBD0 U8347 ( .CLK(n8419), .C(n8431) );
  BUFFD0 U8348 ( .I(n8675), .Z(n8432) );
  CKBD0 U8349 ( .CLK(n8394), .C(n8433) );
  CKBD0 U8350 ( .CLK(n8396), .C(n8434) );
  CKBD0 U8351 ( .CLK(n8424), .C(n8435) );
  CKBD0 U8352 ( .CLK(n8425), .C(n8436) );
  BUFFD0 U8353 ( .I(n8681), .Z(n8437) );
  CKBD0 U8354 ( .CLK(n8426), .C(n8438) );
  CKBD0 U8355 ( .CLK(n8427), .C(n8439) );
  BUFFD0 U8356 ( .I(n8428), .Z(n8440) );
  CKBD0 U8357 ( .CLK(n8429), .C(n8441) );
  BUFFD0 U8358 ( .I(n8430), .Z(n8442) );
  CKBD0 U8359 ( .CLK(n8431), .C(n8443) );
  CKBD0 U8360 ( .CLK(n8399), .C(n8444) );
  BUFFD0 U8361 ( .I(n8346), .Z(n8445) );
  CKBD0 U8362 ( .CLK(n8402), .C(n8446) );
  BUFFD0 U8363 ( .I(n8809), .Z(n8447) );
  CKBD0 U8364 ( .CLK(n8403), .C(n8448) );
  CKBD0 U8365 ( .CLK(n8404), .C(n8449) );
  BUFFD0 U8366 ( .I(n8303), .Z(n8450) );
  CKBD0 U8367 ( .CLK(n8405), .C(n8451) );
  CKBD0 U8368 ( .CLK(n8435), .C(n8452) );
  CKBD0 U8369 ( .CLK(n8436), .C(n8453) );
  CKBD0 U8370 ( .CLK(n8438), .C(n8454) );
  CKBD0 U8371 ( .CLK(n8439), .C(n8455) );
  CKBD0 U8372 ( .CLK(n8440), .C(n8456) );
  CKBD0 U8373 ( .CLK(n8441), .C(n8457) );
  CKBD0 U8374 ( .CLK(n8442), .C(n8458) );
  CKBD0 U8375 ( .CLK(n8443), .C(n8459) );
  CKBD0 U8376 ( .CLK(n8407), .C(n8460) );
  CKBD0 U8377 ( .CLK(n8409), .C(n8461) );
  CKBD0 U8378 ( .CLK(n8453), .C(n8462) );
  CKBD0 U8379 ( .CLK(n8452), .C(n8463) );
  CKBD0 U8380 ( .CLK(n8454), .C(n8464) );
  CKBD0 U8381 ( .CLK(n8455), .C(n8465) );
  CKBD0 U8382 ( .CLK(n8456), .C(n8466) );
  CKBD0 U8383 ( .CLK(n8457), .C(n8467) );
  CKBD0 U8384 ( .CLK(n8458), .C(n8468) );
  BUFFD0 U8385 ( .I(n8462), .Z(n8469) );
  CKBD0 U8386 ( .CLK(n8459), .C(n8470) );
  CKBD0 U8387 ( .CLK(n8463), .C(n8471) );
  CKBD0 U8388 ( .CLK(n8464), .C(n8472) );
  CKBD0 U8389 ( .CLK(n8465), .C(n8473) );
  CKBD0 U8390 ( .CLK(n8466), .C(n8474) );
  CKBD0 U8391 ( .CLK(n8467), .C(n8475) );
  CKBD0 U8392 ( .CLK(n8468), .C(n8476) );
  CKBD0 U8393 ( .CLK(n8469), .C(n8477) );
  CKBD0 U8394 ( .CLK(n8470), .C(n8478) );
  CKBD0 U8395 ( .CLK(n8471), .C(n8479) );
  CKBD0 U8396 ( .CLK(n8472), .C(n8480) );
  CKBD0 U8397 ( .CLK(n8473), .C(n8481) );
  CKBD0 U8398 ( .CLK(n8474), .C(n8482) );
  CKBD0 U8399 ( .CLK(n8475), .C(n8483) );
  CKBD0 U8400 ( .CLK(n8476), .C(n8484) );
  CKBD0 U8401 ( .CLK(n8478), .C(n8485) );
  CKBD0 U8402 ( .CLK(n8477), .C(n8486) );
  CKBD0 U8403 ( .CLK(n8479), .C(n8487) );
  CKBD0 U8404 ( .CLK(n8480), .C(n8488) );
  CKBD0 U8405 ( .CLK(n8481), .C(n8489) );
  CKBD0 U8406 ( .CLK(n8482), .C(n8490) );
  CKBD0 U8407 ( .CLK(n8483), .C(n8491) );
  CKBD0 U8408 ( .CLK(n8484), .C(n8492) );
  CKBD0 U8409 ( .CLK(n8410), .C(n8493) );
  CKBD0 U8410 ( .CLK(n8411), .C(n8494) );
  BUFFD0 U8411 ( .I(n8973), .Z(n8495) );
  BUFFD0 U8412 ( .I(n8485), .Z(n8496) );
  CKBD0 U8413 ( .CLK(n8486), .C(n8497) );
  CKBD0 U8414 ( .CLK(n8487), .C(n8498) );
  CKBD0 U8415 ( .CLK(n8488), .C(n8499) );
  CKBD0 U8416 ( .CLK(n8489), .C(n8500) );
  CKBD0 U8417 ( .CLK(n8490), .C(n8501) );
  CKBD0 U8418 ( .CLK(n8491), .C(n8502) );
  CKBD0 U8419 ( .CLK(n8492), .C(n8503) );
  CKBD0 U8420 ( .CLK(n8496), .C(n8504) );
  CKBD0 U8421 ( .CLK(n8497), .C(n8505) );
  CKBD0 U8422 ( .CLK(n8498), .C(n8506) );
  CKBD0 U8423 ( .CLK(n8499), .C(n8507) );
  CKBD0 U8424 ( .CLK(n8500), .C(n8508) );
  CKBD0 U8425 ( .CLK(n8501), .C(n8509) );
  CKBD0 U8426 ( .CLK(n8502), .C(n8510) );
  CKBD0 U8427 ( .CLK(n8503), .C(n8511) );
  CKBD0 U8428 ( .CLK(n8504), .C(n8512) );
  CKBD0 U8429 ( .CLK(n8505), .C(n8513) );
  CKBD0 U8430 ( .CLK(n8506), .C(n8514) );
  CKBD0 U8431 ( .CLK(n8507), .C(n8515) );
  BUFFD0 U8432 ( .I(n8508), .Z(n8516) );
  CKBD0 U8433 ( .CLK(n8509), .C(n8517) );
  BUFFD0 U8434 ( .I(n8554), .Z(n8518) );
  CKBD0 U8435 ( .CLK(n8415), .C(n8519) );
  CKBD0 U8436 ( .CLK(n8510), .C(n8520) );
  CKBD0 U8437 ( .CLK(n8511), .C(n8521) );
  CKBD0 U8438 ( .CLK(n8512), .C(n8522) );
  CKBD0 U8439 ( .CLK(n8513), .C(n8523) );
  BUFFD0 U8440 ( .I(n8562), .Z(n8524) );
  CKBD0 U8441 ( .CLK(n8514), .C(n8525) );
  BUFFD0 U8442 ( .I(n8388), .Z(n8526) );
  BUFFD0 U8443 ( .I(n8390), .Z(n8527) );
  BUFFD0 U8444 ( .I(n8422), .Z(n8528) );
  CKBD0 U8445 ( .CLK(n8423), .C(n8529) );
  BUFFD0 U8446 ( .I(n8720), .Z(n8530) );
  BUFFD0 U8447 ( .I(n8393), .Z(n8531) );
  CKBD0 U8448 ( .CLK(n8515), .C(n8532) );
  BUFFD0 U8449 ( .I(n8434), .Z(n8533) );
  CKBD0 U8450 ( .CLK(n8516), .C(n8534) );
  BUFFD0 U8451 ( .I(n8327), .Z(n8535) );
  BUFFD0 U8452 ( .I(n8879), .Z(n8536) );
  CKBD0 U8453 ( .CLK(n8445), .C(n8537) );
  BUFFD0 U8454 ( .I(n8400), .Z(n8538) );
  BUFFD0 U8455 ( .I(n8775), .Z(n8539) );
  BUFFD0 U8456 ( .I(n8444), .Z(n8540) );
  CKBD0 U8457 ( .CLK(n8517), .C(n8541) );
  CKBD0 U8458 ( .CLK(n8520), .C(n8542) );
  CKBD0 U8459 ( .CLK(n8521), .C(n8543) );
  CKBD0 U8460 ( .CLK(n8522), .C(n8544) );
  BUFFD0 U8461 ( .I(n8525), .Z(n8545) );
  CKBD0 U8462 ( .CLK(n8523), .C(n8546) );
  CKBD0 U8463 ( .CLK(n8532), .C(n8547) );
  CKBD0 U8464 ( .CLK(n8450), .C(n8548) );
  BUFFD0 U8465 ( .I(n8460), .Z(n8549) );
  BUFFD0 U8466 ( .I(n8645), .Z(n8550) );
  BUFFD0 U8467 ( .I(n8448), .Z(n8551) );
  CKBD0 U8468 ( .CLK(n8534), .C(n8552) );
  BUFFD0 U8469 ( .I(n8651), .Z(n8553) );
  BUFFD0 U8470 ( .I(n8862), .Z(n8554) );
  BUFFD0 U8471 ( .I(n8461), .Z(n8555) );
  BUFFD0 U8472 ( .I(n8494), .Z(n8556) );
  BUFFD0 U8473 ( .I(n8412), .Z(n8557) );
  BUFFD0 U8474 ( .I(n8661), .Z(n8558) );
  CKBD0 U8475 ( .CLK(n8541), .C(n8559) );
  BUFFD0 U8476 ( .I(n8542), .Z(n8560) );
  BUFFD0 U8477 ( .I(n8543), .Z(n8561) );
  BUFFD0 U8478 ( .I(n8667), .Z(n8562) );
  CKBD0 U8479 ( .CLK(n8544), .C(n8563) );
  CKBD0 U8480 ( .CLK(n8526), .C(n8564) );
  CKBD0 U8481 ( .CLK(n8527), .C(n8565) );
  CKBD0 U8482 ( .CLK(n8528), .C(n8566) );
  CKBD0 U8483 ( .CLK(n8545), .C(n8567) );
  CKBD0 U8484 ( .CLK(n8546), .C(n8568) );
  BUFFD0 U8485 ( .I(n8529), .Z(n8569) );
  BUFFD0 U8486 ( .I(n8547), .Z(n8570) );
  CKBD0 U8487 ( .CLK(n8552), .C(n8571) );
  BUFFD0 U8488 ( .I(n8559), .Z(n8572) );
  CKBD0 U8489 ( .CLK(n8560), .C(n8573) );
  CKBD0 U8490 ( .CLK(n8561), .C(n8574) );
  CKBD0 U8491 ( .CLK(n8563), .C(n8575) );
  CKBD0 U8492 ( .CLK(n8531), .C(n8576) );
  BUFFD0 U8493 ( .I(n8433), .Z(n8577) );
  CKBD0 U8494 ( .CLK(n8533), .C(n8578) );
  CKBD0 U8495 ( .CLK(n8535), .C(n8579) );
  CKBD0 U8496 ( .CLK(n8567), .C(n8580) );
  CKBD0 U8497 ( .CLK(n8568), .C(n8581) );
  CKBD0 U8498 ( .CLK(n8570), .C(n8582) );
  CKBD0 U8499 ( .CLK(n8571), .C(n8583) );
  CKBD0 U8500 ( .CLK(n8572), .C(n8584) );
  CKBD0 U8501 ( .CLK(n8573), .C(n8585) );
  CKBD0 U8502 ( .CLK(n8574), .C(n8586) );
  CKBD0 U8503 ( .CLK(n8575), .C(n8587) );
  BUFFD0 U8504 ( .I(n8836), .Z(n8588) );
  CKBD0 U8505 ( .CLK(n8538), .C(n8589) );
  CKBD0 U8506 ( .CLK(n8581), .C(n8590) );
  CKBD0 U8507 ( .CLK(n8580), .C(n8591) );
  CKBD0 U8508 ( .CLK(n8582), .C(n8592) );
  CKBD0 U8509 ( .CLK(n8583), .C(n8593) );
  CKBD0 U8510 ( .CLK(n8584), .C(n8594) );
  CKBD0 U8511 ( .CLK(n8585), .C(n8595) );
  CKBD0 U8512 ( .CLK(n8586), .C(n8596) );
  BUFFD0 U8513 ( .I(n8590), .Z(n8597) );
  CKBD0 U8514 ( .CLK(n8587), .C(n8598) );
  CKBD0 U8515 ( .CLK(n8591), .C(n8599) );
  CKBD0 U8516 ( .CLK(n8592), .C(n8600) );
  CKBD0 U8517 ( .CLK(n8593), .C(n8601) );
  CKBD0 U8518 ( .CLK(n8594), .C(n8602) );
  CKBD0 U8519 ( .CLK(n8595), .C(n8603) );
  CKBD0 U8520 ( .CLK(n8596), .C(n8604) );
  CKBD0 U8521 ( .CLK(n8597), .C(n8605) );
  CKBD0 U8522 ( .CLK(n8598), .C(n8606) );
  CKBD0 U8523 ( .CLK(n8599), .C(n8607) );
  CKBD0 U8524 ( .CLK(n8600), .C(n8608) );
  CKBD0 U8525 ( .CLK(n8601), .C(n8609) );
  CKBD0 U8526 ( .CLK(n8602), .C(n8610) );
  CKBD0 U8527 ( .CLK(n8603), .C(n8611) );
  CKBD0 U8528 ( .CLK(n8604), .C(n8612) );
  CKBD0 U8529 ( .CLK(n8606), .C(n8613) );
  CKBD0 U8530 ( .CLK(n8605), .C(n8614) );
  CKBD0 U8531 ( .CLK(n8607), .C(n8615) );
  CKBD0 U8532 ( .CLK(n8608), .C(n8616) );
  CKBD0 U8533 ( .CLK(n8609), .C(n8617) );
  CKBD0 U8534 ( .CLK(n8610), .C(n8618) );
  CKBD0 U8535 ( .CLK(n8611), .C(n8619) );
  CKBD0 U8536 ( .CLK(n8612), .C(n8620) );
  CKBD0 U8537 ( .CLK(n8540), .C(n8621) );
  BUFFD0 U8538 ( .I(n8613), .Z(n8622) );
  CKBD0 U8539 ( .CLK(n8614), .C(n8623) );
  CKBD0 U8540 ( .CLK(n8615), .C(n8624) );
  CKBD0 U8541 ( .CLK(n8616), .C(n8625) );
  CKBD0 U8542 ( .CLK(n8617), .C(n8626) );
  CKBD0 U8543 ( .CLK(n8618), .C(n8627) );
  CKBD0 U8544 ( .CLK(n8619), .C(n8628) );
  CKBD0 U8545 ( .CLK(n8620), .C(n8629) );
  CKBD0 U8546 ( .CLK(n8622), .C(n8630) );
  CKBD0 U8547 ( .CLK(n8623), .C(n8631) );
  CKBD0 U8548 ( .CLK(n8624), .C(n8632) );
  CKBD0 U8549 ( .CLK(n8625), .C(n8633) );
  CKBD0 U8550 ( .CLK(n8626), .C(n8634) );
  CKBD0 U8551 ( .CLK(n8627), .C(n8635) );
  BUFFD0 U8552 ( .I(n8446), .Z(n8636) );
  CKBD0 U8553 ( .CLK(n8628), .C(n8637) );
  CKBD0 U8554 ( .CLK(n8629), .C(n8638) );
  CKBD0 U8555 ( .CLK(n8630), .C(n8639) );
  CKBD0 U8556 ( .CLK(n8631), .C(n8640) );
  CKBD0 U8557 ( .CLK(n8632), .C(n8641) );
  CKBD0 U8558 ( .CLK(n8633), .C(n8642) );
  CKBD0 U8559 ( .CLK(n8634), .C(n8643) );
  CKBD0 U8560 ( .CLK(n8635), .C(n8644) );
  BUFFD0 U8561 ( .I(n8967), .Z(n8645) );
  BUFFD0 U8562 ( .I(n8449), .Z(n8646) );
  CKBD0 U8563 ( .CLK(n8549), .C(n8647) );
  BUFFD0 U8564 ( .I(n8414), .Z(n8648) );
  CKBD0 U8565 ( .CLK(n8551), .C(n8649) );
  BUFFD0 U8566 ( .I(n8548), .Z(n8650) );
  BUFFD0 U8567 ( .I(n8700), .Z(n8651) );
  CKBD0 U8568 ( .CLK(n8637), .C(n8652) );
  CKBD0 U8569 ( .CLK(n8638), .C(n8653) );
  CKBD0 U8570 ( .CLK(n8639), .C(n8654) );
  CKBD0 U8571 ( .CLK(n8640), .C(n8655) );
  BUFFD0 U8572 ( .I(n8642), .Z(n8656) );
  CKBD0 U8573 ( .CLK(n8641), .C(n8657) );
  BUFFD0 U8574 ( .I(n8643), .Z(n8658) );
  CKBD0 U8575 ( .CLK(n8644), .C(n8659) );
  CKBD0 U8576 ( .CLK(n8555), .C(n8660) );
  BUFFD0 U8577 ( .I(n8690), .Z(n8661) );
  CKBD0 U8578 ( .CLK(n8556), .C(n8662) );
  CKBD0 U8579 ( .CLK(n8557), .C(n8663) );
  CKBD0 U8580 ( .CLK(n8652), .C(n8664) );
  CKBD0 U8581 ( .CLK(n8653), .C(n8665) );
  CKBD0 U8582 ( .CLK(n8654), .C(n8666) );
  BUFFD0 U8583 ( .I(n8988), .Z(n8667) );
  CKBD0 U8584 ( .CLK(n8655), .C(n8668) );
  CKBD0 U8585 ( .CLK(n8657), .C(n8669) );
  CKBD0 U8586 ( .CLK(n8656), .C(n8670) );
  BUFFD0 U8587 ( .I(n8564), .Z(n8671) );
  BUFFD0 U8588 ( .I(n8565), .Z(n8672) );
  BUFFD0 U8589 ( .I(n8566), .Z(n8673) );
  CKBD0 U8590 ( .CLK(n8569), .C(n8674) );
  BUFFD0 U8591 ( .I(n8996), .Z(n8675) );
  BUFFD0 U8592 ( .I(n8579), .Z(n8676) );
  CKBD0 U8593 ( .CLK(n8577), .C(n8677) );
  BUFFD0 U8594 ( .I(n8732), .Z(n8678) );
  CKBD0 U8595 ( .CLK(n8658), .C(n8679) );
  BUFFD0 U8596 ( .I(n8855), .Z(n8680) );
  BUFFD0 U8597 ( .I(n8772), .Z(n8681) );
  BUFFD0 U8598 ( .I(n8878), .Z(n8682) );
  BUFFD0 U8599 ( .I(n8537), .Z(n8683) );
  CKBD0 U8600 ( .CLK(n8636), .C(n8684) );
  CKBD0 U8601 ( .CLK(n8646), .C(n8685) );
  BUFFD0 U8602 ( .I(n8659), .Z(n8686) );
  CKBD0 U8603 ( .CLK(n8650), .C(n8687) );
  CKBD0 U8604 ( .CLK(n8648), .C(n8688) );
  BUFFD0 U8605 ( .I(n8451), .Z(n8689) );
  BUFFD0 U8606 ( .I(n8771), .Z(n8690) );
  BUFFD0 U8607 ( .I(n8664), .Z(n8691) );
  CKBD0 U8608 ( .CLK(n8665), .C(n8692) );
  CKBD0 U8609 ( .CLK(n8666), .C(n8693) );
  BUFFD0 U8610 ( .I(n8669), .Z(n8694) );
  CKBD0 U8611 ( .CLK(n8668), .C(n8695) );
  CKBD0 U8612 ( .CLK(n8670), .C(n8696) );
  CKBD0 U8613 ( .CLK(n8679), .C(n8697) );
  BUFFD0 U8614 ( .I(n8649), .Z(n8698) );
  CKBD0 U8615 ( .CLK(n8686), .C(n8699) );
  BUFFD0 U8616 ( .I(n8789), .Z(n8700) );
  CKBD0 U8617 ( .CLK(n8691), .C(n8701) );
  CKBD0 U8618 ( .CLK(n8692), .C(n8702) );
  CKBD0 U8619 ( .CLK(n8693), .C(n8703) );
  CKBD0 U8620 ( .CLK(n8694), .C(n8704) );
  CKBD0 U8621 ( .CLK(n8695), .C(n8705) );
  CKBD0 U8622 ( .CLK(n8696), .C(n8706) );
  CKBD0 U8623 ( .CLK(n8697), .C(n8707) );
  BUFFD0 U8624 ( .I(n8790), .Z(n8708) );
  BUFFD0 U8625 ( .I(n8662), .Z(n8709) );
  BUFFD0 U8626 ( .I(n8663), .Z(n8710) );
  CKBD0 U8627 ( .CLK(n8699), .C(n8711) );
  CKBD0 U8628 ( .CLK(n8701), .C(n8712) );
  BUFFD0 U8629 ( .I(n8702), .Z(n8713) );
  BUFFD0 U8630 ( .I(n8418), .Z(n8714) );
  CKBD0 U8631 ( .CLK(n8703), .C(n8715) );
  CKBD0 U8632 ( .CLK(n8671), .C(n8716) );
  CKBD0 U8633 ( .CLK(n8672), .C(n8717) );
  CKBD0 U8634 ( .CLK(n8673), .C(n8718) );
  CKBD0 U8635 ( .CLK(n8704), .C(n8719) );
  BUFFD0 U8636 ( .I(n8827), .Z(n8720) );
  BUFFD0 U8637 ( .I(n8647), .Z(n8721) );
  BUFFD0 U8638 ( .I(n8674), .Z(n8722) );
  CKBD0 U8639 ( .CLK(n8676), .C(n8723) );
  CKBD0 U8640 ( .CLK(n8705), .C(n8724) );
  BUFFD0 U8641 ( .I(n8576), .Z(n8725) );
  CKBD0 U8642 ( .CLK(n8706), .C(n8726) );
  CKBD0 U8643 ( .CLK(n8707), .C(n8727) );
  CKBD0 U8644 ( .CLK(n8711), .C(n8728) );
  CKBD0 U8645 ( .CLK(n8712), .C(n8729) );
  CKBD0 U8646 ( .CLK(n8713), .C(n8730) );
  CKBD0 U8647 ( .CLK(n8715), .C(n8731) );
  BUFFD0 U8648 ( .I(n8958), .Z(n8732) );
  CKBD0 U8649 ( .CLK(n8724), .C(n8733) );
  CKBD0 U8650 ( .CLK(n8719), .C(n8734) );
  CKBD0 U8651 ( .CLK(n8726), .C(n8735) );
  CKBD0 U8652 ( .CLK(n8727), .C(n8736) );
  CKBD0 U8653 ( .CLK(n8728), .C(n8737) );
  CKBD0 U8654 ( .CLK(n8729), .C(n8738) );
  CKBD0 U8655 ( .CLK(n8730), .C(n8739) );
  BUFFD0 U8656 ( .I(n8733), .Z(n8740) );
  CKBD0 U8657 ( .CLK(n8731), .C(n8741) );
  CKBD0 U8658 ( .CLK(n8734), .C(n8742) );
  CKBD0 U8659 ( .CLK(n8735), .C(n8743) );
  CKBD0 U8660 ( .CLK(n8736), .C(n8744) );
  CKBD0 U8661 ( .CLK(n8737), .C(n8745) );
  CKBD0 U8662 ( .CLK(n8738), .C(n8746) );
  CKBD0 U8663 ( .CLK(n8739), .C(n8747) );
  CKBD0 U8664 ( .CLK(n8741), .C(n8748) );
  CKBD0 U8665 ( .CLK(n8740), .C(n8749) );
  CKBD0 U8666 ( .CLK(n8742), .C(n8750) );
  CKBD0 U8667 ( .CLK(n8743), .C(n8751) );
  CKBD0 U8668 ( .CLK(n8744), .C(n8752) );
  CKBD0 U8669 ( .CLK(n8745), .C(n8753) );
  CKBD0 U8670 ( .CLK(n8746), .C(n8754) );
  CKBD0 U8671 ( .CLK(n8747), .C(n8755) );
  BUFFD0 U8672 ( .I(n8748), .Z(n8756) );
  CKBD0 U8673 ( .CLK(n8749), .C(n8757) );
  CKBD0 U8674 ( .CLK(n8750), .C(n8758) );
  CKBD0 U8675 ( .CLK(n8751), .C(n8759) );
  CKBD0 U8676 ( .CLK(n8752), .C(n8760) );
  CKBD0 U8677 ( .CLK(n8753), .C(n8761) );
  CKBD0 U8678 ( .CLK(n8754), .C(n8762) );
  CKBD0 U8679 ( .CLK(n8755), .C(n8763) );
  CKBD0 U8680 ( .CLK(n8756), .C(n8764) );
  CKBD0 U8681 ( .CLK(n8757), .C(n8765) );
  CKBD0 U8682 ( .CLK(n8758), .C(n8766) );
  CKBD0 U8683 ( .CLK(n8759), .C(n8767) );
  CKBD0 U8684 ( .CLK(n8760), .C(n8768) );
  CKBD0 U8685 ( .CLK(n8761), .C(n8769) );
  CKBD0 U8686 ( .CLK(n8762), .C(n8770) );
  BUFFD0 U8687 ( .I(n8828), .Z(n8771) );
  BUFFD0 U8688 ( .I(n8833), .Z(n8772) );
  BUFFD0 U8689 ( .I(n8688), .Z(n8773) );
  CKBD0 U8690 ( .CLK(n8683), .C(n8774) );
  BUFFD0 U8691 ( .I(n8837), .Z(n8775) );
  BUFFD0 U8692 ( .I(n8621), .Z(n8776) );
  CKBD0 U8693 ( .CLK(n8763), .C(n8777) );
  CKBD0 U8694 ( .CLK(n8764), .C(n8778) );
  CKBD0 U8695 ( .CLK(n8765), .C(n8779) );
  CKBD0 U8696 ( .CLK(n8766), .C(n8780) );
  CKBD0 U8697 ( .CLK(n8767), .C(n8781) );
  BUFFD0 U8698 ( .I(n8768), .Z(n8782) );
  CKBD0 U8699 ( .CLK(n8769), .C(n8783) );
  CKBD0 U8700 ( .CLK(n8770), .C(n8784) );
  BUFFD0 U8701 ( .I(n8684), .Z(n8785) );
  CKBD0 U8702 ( .CLK(n8689), .C(n8786) );
  CKBD0 U8703 ( .CLK(n8698), .C(n8787) );
  BUFFD0 U8704 ( .I(n8687), .Z(n8788) );
  BUFFD0 U8705 ( .I(n8956), .Z(n8789) );
  BUFFD0 U8706 ( .I(n8974), .Z(n8790) );
  CKBD0 U8707 ( .CLK(n8777), .C(n8791) );
  CKBD0 U8708 ( .CLK(n8709), .C(n8792) );
  CKBD0 U8709 ( .CLK(n8710), .C(n8793) );
  CKBD0 U8710 ( .CLK(n8778), .C(n8794) );
  BUFFD0 U8711 ( .I(n8780), .Z(n8795) );
  CKBD0 U8712 ( .CLK(n8779), .C(n8796) );
  CKBD0 U8713 ( .CLK(n8781), .C(n8797) );
  CKBD0 U8714 ( .CLK(n8782), .C(n8798) );
  CKBD0 U8715 ( .CLK(n8783), .C(n8799) );
  BUFFD0 U8716 ( .I(n8784), .Z(n8800) );
  CKBD0 U8717 ( .CLK(n8791), .C(n8801) );
  CKBD0 U8718 ( .CLK(n8794), .C(n8802) );
  CKBD0 U8719 ( .CLK(n8795), .C(n8803) );
  CKBD0 U8720 ( .CLK(n8796), .C(n8804) );
  BUFFD0 U8721 ( .I(n8797), .Z(n8805) );
  CKBD0 U8722 ( .CLK(n8714), .C(n8806) );
  CKBD0 U8723 ( .CLK(n8798), .C(n8807) );
  BUFFD0 U8724 ( .I(n8990), .Z(n8808) );
  BUFFD0 U8725 ( .I(n8979), .Z(n8809) );
  BUFFD0 U8726 ( .I(n8799), .Z(n8810) );
  CKBD0 U8727 ( .CLK(n8800), .C(n8811) );
  CKBD0 U8728 ( .CLK(n8801), .C(n8812) );
  CKBD0 U8729 ( .CLK(n8802), .C(n8813) );
  CKBD0 U8730 ( .CLK(n8804), .C(n8814) );
  CKBD0 U8731 ( .CLK(n8803), .C(n8815) );
  CKBD0 U8732 ( .CLK(n8805), .C(n8816) );
  CKBD0 U8733 ( .CLK(n8807), .C(n8817) );
  CKBD0 U8734 ( .CLK(n8810), .C(n8818) );
  CKBD0 U8735 ( .CLK(n8811), .C(n8819) );
  BUFFD0 U8736 ( .I(n8812), .Z(n8820) );
  CKBD0 U8737 ( .CLK(n8813), .C(n8821) );
  BUFFD0 U8738 ( .I(n8814), .Z(n8822) );
  CKBD0 U8739 ( .CLK(n8815), .C(n8823) );
  BUFFD0 U8740 ( .I(n8991), .Z(n8824) );
  CKBD0 U8741 ( .CLK(n8816), .C(n8825) );
  BUFFD0 U8742 ( .I(n8718), .Z(n8826) );
  BUFFD0 U8743 ( .I(n8989), .Z(n8827) );
  BUFFD0 U8744 ( .I(n8982), .Z(n8828) );
  CKBD0 U8745 ( .CLK(n8722), .C(n8829) );
  CKBD0 U8746 ( .CLK(n8721), .C(n8830) );
  CKBD0 U8747 ( .CLK(n8725), .C(n8831) );
  BUFFD0 U8748 ( .I(n8578), .Z(n8832) );
  BUFFD0 U8749 ( .I(n8866), .Z(n8833) );
  CKBD0 U8750 ( .CLK(n8817), .C(n8834) );
  CKBD0 U8751 ( .CLK(n8773), .C(n8835) );
  BUFFD0 U8752 ( .I(n8867), .Z(n8836) );
  BUFFD0 U8753 ( .I(n8869), .Z(n8837) );
  CKBD0 U8754 ( .CLK(n8776), .C(n8838) );
  CKBD0 U8755 ( .CLK(n8785), .C(n8839) );
  CKBD0 U8756 ( .CLK(n8788), .C(n8840) );
  BUFFD0 U8757 ( .I(n8786), .Z(n8841) );
  CKBD0 U8758 ( .CLK(n8818), .C(n8842) );
  BUFFD0 U8759 ( .I(n8787), .Z(n8843) );
  BUFFD0 U8760 ( .I(n8493), .Z(n8844) );
  BUFFD0 U8761 ( .I(n8660), .Z(n8845) );
  BUFFD0 U8762 ( .I(n9013), .Z(n8846) );
  BUFFD0 U8763 ( .I(n8793), .Z(n8847) );
  CKBD0 U8764 ( .CLK(n8819), .C(n8848) );
  CKBD0 U8765 ( .CLK(n8820), .C(n8849) );
  BUFFD0 U8766 ( .I(n8821), .Z(n8850) );
  CKBD0 U8767 ( .CLK(n8822), .C(n8851) );
  BUFFD0 U8768 ( .I(n8723), .Z(n8852) );
  BUFFD0 U8769 ( .I(n8806), .Z(n8853) );
  CKBD0 U8770 ( .CLK(n8823), .C(n8854) );
  BUFFD0 U8771 ( .I(n8900), .Z(n8855) );
  BUFFD0 U8772 ( .I(n8519), .Z(n8856) );
  BUFFD0 U8773 ( .I(n8716), .Z(n8857) );
  BUFFD0 U8774 ( .I(n8717), .Z(n8858) );
  CKBD0 U8775 ( .CLK(n8825), .C(n8859) );
  CKBD0 U8776 ( .CLK(n8826), .C(n8860) );
  BUFFD0 U8777 ( .I(n8677), .Z(n8861) );
  BUFFD0 U8778 ( .I(n8903), .Z(n8862) );
  BUFFD0 U8779 ( .I(n8829), .Z(n8863) );
  BUFFD0 U8780 ( .I(n8831), .Z(n8864) );
  CKBD0 U8781 ( .CLK(n8832), .C(n8865) );
  BUFFD0 U8782 ( .I(n8957), .Z(n8866) );
  BUFFD0 U8783 ( .I(n8950), .Z(n8867) );
  CKBD0 U8784 ( .CLK(n8834), .C(n8868) );
  BUFFD0 U8785 ( .I(n8968), .Z(n8869) );
  CKBD0 U8786 ( .CLK(n8842), .C(n8870) );
  CKBD0 U8787 ( .CLK(n8848), .C(n8871) );
  CKBD0 U8788 ( .CLK(n8849), .C(n8872) );
  CKBD0 U8789 ( .CLK(n8850), .C(n8873) );
  BUFFD0 U8790 ( .I(n8851), .Z(n8874) );
  BUFFD0 U8791 ( .I(n8889), .Z(n8875) );
  CKBD0 U8792 ( .CLK(n8854), .C(n8876) );
  BUFFD0 U8793 ( .I(n8868), .Z(n8877) );
  BUFFD0 U8794 ( .I(n8969), .Z(n8878) );
  BUFFD0 U8795 ( .I(n8970), .Z(n8879) );
  BUFFD0 U8796 ( .I(n8972), .Z(n8880) );
  CKBD0 U8797 ( .CLK(n8841), .C(n8881) );
  BUFFD0 U8798 ( .I(n8940), .Z(n8882) );
  CKBD0 U8799 ( .CLK(n8843), .C(n8883) );
  CKBD0 U8800 ( .CLK(n8844), .C(n8884) );
  CKBD0 U8801 ( .CLK(n8871), .C(n8885) );
  CKBD0 U8802 ( .CLK(n8872), .C(n8886) );
  BUFFD0 U8803 ( .I(n8873), .Z(n8887) );
  CKBD0 U8804 ( .CLK(n8874), .C(n8888) );
  BUFFD0 U8805 ( .I(n8938), .Z(n8889) );
  BUFFD0 U8806 ( .I(n8876), .Z(n8890) );
  CKBD0 U8807 ( .CLK(n8877), .C(n8891) );
  BUFFD0 U8808 ( .I(n8870), .Z(n8892) );
  CKBD0 U8809 ( .CLK(n8845), .C(n8893) );
  CKBD0 U8810 ( .CLK(n8847), .C(n8894) );
  BUFFD0 U8811 ( .I(n8792), .Z(n8895) );
  BUFFD0 U8812 ( .I(n8885), .Z(n8896) );
  BUFFD0 U8813 ( .I(n8908), .Z(n8897) );
  CKBD0 U8814 ( .CLK(n8887), .C(n8898) );
  BUFFD0 U8815 ( .I(n8888), .Z(n8899) );
  BUFFD0 U8816 ( .I(n8978), .Z(n8900) );
  CKBD0 U8817 ( .CLK(n8852), .C(n8901) );
  BUFFD0 U8818 ( .I(n8859), .Z(n8902) );
  BUFFD0 U8819 ( .I(n8980), .Z(n8903) );
  CKBD0 U8820 ( .CLK(n8856), .C(n8904) );
  CKBD0 U8821 ( .CLK(n8890), .C(n8905) );
  BUFFD0 U8822 ( .I(n8930), .Z(n8906) );
  CKBD0 U8823 ( .CLK(n8892), .C(n8907) );
  BUFFD0 U8824 ( .I(n8932), .Z(n8908) );
  CKBD0 U8825 ( .CLK(n8896), .C(n8909) );
  BUFFD0 U8826 ( .I(n8961), .Z(n8910) );
  CKBD0 U8827 ( .CLK(n8899), .C(n8911) );
  CKBD0 U8828 ( .CLK(n8902), .C(n8912) );
  BUFFD0 U8829 ( .I(n8920), .Z(n8913) );
  BUFFD0 U8830 ( .I(n8891), .Z(n8914) );
  BUFFD0 U8831 ( .I(n8907), .Z(n8915) );
  BUFFD0 U8832 ( .I(n8941), .Z(n8916) );
  BUFFD0 U8833 ( .I(n8886), .Z(n8917) );
  BUFFD0 U8834 ( .I(n8898), .Z(n8918) );
  BUFFD0 U8835 ( .I(n9011), .Z(n8919) );
  BUFFD0 U8836 ( .I(n8928), .Z(n8920) );
  BUFFD0 U8837 ( .I(n8912), .Z(n8921) );
  CKBD0 U8838 ( .CLK(n8914), .C(n8922) );
  CKBD0 U8839 ( .CLK(n8915), .C(n8923) );
  BUFFD0 U8840 ( .I(n8909), .Z(n8924) );
  CKBD0 U8841 ( .CLK(n8917), .C(n8925) );
  CKBD0 U8842 ( .CLK(n8918), .C(n8926) );
  BUFFD0 U8843 ( .I(n8911), .Z(n8927) );
  BUFFD0 U8844 ( .I(n8936), .Z(n8928) );
  CKBD0 U8845 ( .CLK(n8921), .C(n8929) );
  BUFFD0 U8846 ( .I(n8965), .Z(n8930) );
  BUFFD0 U8847 ( .I(n8923), .Z(n8931) );
  BUFFD0 U8848 ( .I(n8976), .Z(n8932) );
  CKBD0 U8849 ( .CLK(n8924), .C(n8933) );
  BUFFD0 U8850 ( .I(n8926), .Z(n8934) );
  CKBD0 U8851 ( .CLK(n8853), .C(n8935) );
  BUFFD0 U8852 ( .I(n9010), .Z(n8936) );
  CKBD0 U8853 ( .CLK(n8927), .C(n8937) );
  BUFFD0 U8854 ( .I(n9012), .Z(n8938) );
  BUFFD0 U8855 ( .I(n8922), .Z(n8939) );
  BUFFD0 U8856 ( .I(n9015), .Z(n8940) );
  BUFFD0 U8857 ( .I(n8959), .Z(n8941) );
  BUFFD0 U8858 ( .I(n8925), .Z(n8942) );
  CKBD0 U8859 ( .CLK(n8934), .C(n8943) );
  BUFFD0 U8860 ( .I(n8905), .Z(n8944) );
  BUFFD0 U8861 ( .I(n8937), .Z(n8945) );
  CKBD0 U8862 ( .CLK(n8861), .C(n8946) );
  CKBD0 U8863 ( .CLK(n8857), .C(n8947) );
  CKBD0 U8864 ( .CLK(n8858), .C(n8948) );
  BUFFD0 U8865 ( .I(n8929), .Z(n8949) );
  BUFFD0 U8866 ( .I(n8992), .Z(n8950) );
  CKBD0 U8867 ( .CLK(n8863), .C(n8951) );
  CKBD0 U8868 ( .CLK(n8864), .C(n8952) );
  CKBD0 U8869 ( .CLK(n8939), .C(n8953) );
  BUFFD0 U8870 ( .I(n8860), .Z(n8954) );
  BUFFD0 U8871 ( .I(n8931), .Z(n8955) );
  BUFFD0 U8872 ( .I(n9009), .Z(n8956) );
  BUFFD0 U8873 ( .I(n8589), .Z(n8957) );
  BUFFD0 U8874 ( .I(n8865), .Z(n8958) );
  BUFFD0 U8875 ( .I(n8975), .Z(n8959) );
  CKBD0 U8876 ( .CLK(n8942), .C(n8960) );
  BUFFD0 U8877 ( .I(n9007), .Z(n8961) );
  CKBD0 U8878 ( .CLK(n8944), .C(n8962) );
  CKBD0 U8879 ( .CLK(n8945), .C(n8963) );
  CKBD0 U8880 ( .CLK(n8949), .C(n8964) );
  BUFFD0 U8881 ( .I(n9014), .Z(n8965) );
  CKBD0 U8882 ( .CLK(n8955), .C(n8966) );
  BUFFD0 U8883 ( .I(n9008), .Z(n8967) );
  BUFFD0 U8884 ( .I(n8685), .Z(n8968) );
  BUFFD0 U8885 ( .I(n8997), .Z(n8969) );
  BUFFD0 U8886 ( .I(n8839), .Z(n8970) );
  BUFFD0 U8887 ( .I(n8883), .Z(n8971) );
  BUFFD0 U8888 ( .I(n8840), .Z(n8972) );
  BUFFD0 U8889 ( .I(n8894), .Z(n8973) );
  BUFFD0 U8890 ( .I(n8893), .Z(n8974) );
  BUFFD0 U8891 ( .I(n9016), .Z(n8975) );
  BUFFD0 U8892 ( .I(n9017), .Z(n8976) );
  CKBD0 U8893 ( .CLK(n8895), .C(n8977) );
  BUFFD0 U8894 ( .I(n8830), .Z(n8978) );
  BUFFD0 U8895 ( .I(n8901), .Z(n8979) );
  BUFFD0 U8896 ( .I(n8835), .Z(n8980) );
  BUFFD0 U8897 ( .I(n8943), .Z(n8981) );
  BUFFD0 U8898 ( .I(n8904), .Z(n8982) );
  BUFFD0 U8899 ( .I(n8962), .Z(n8983) );
  BUFFD0 U8900 ( .I(n8963), .Z(n8984) );
  BUFFD0 U8901 ( .I(n8964), .Z(n8985) );
  BUFFD0 U8902 ( .I(n8953), .Z(n8986) );
  BUFFD0 U8903 ( .I(n8966), .Z(n8987) );
  BUFFD0 U8904 ( .I(n8935), .Z(n8988) );
  BUFFD0 U8905 ( .I(n8946), .Z(n8989) );
  BUFFD0 U8906 ( .I(n8947), .Z(n8990) );
  BUFFD0 U8907 ( .I(n8948), .Z(n8991) );
  BUFFD0 U8908 ( .I(n8774), .Z(n8992) );
  BUFFD0 U8909 ( .I(n8951), .Z(n8993) );
  BUFFD0 U8910 ( .I(n8933), .Z(n8994) );
  BUFFD0 U8911 ( .I(n8960), .Z(n8995) );
  BUFFD0 U8912 ( .I(n8952), .Z(n8996) );
  BUFFD0 U8913 ( .I(n8838), .Z(n8997) );
  CKBD0 U8914 ( .CLK(n8981), .C(n8998) );
  CKBD0 U8915 ( .CLK(n8983), .C(n8999) );
  CKBD0 U8916 ( .CLK(n8984), .C(n9000) );
  BUFFD0 U8917 ( .I(n9125), .Z(n9001) );
  CKBD0 U8918 ( .CLK(n8985), .C(n9002) );
  CKBD0 U8919 ( .CLK(n8986), .C(n9003) );
  CKBD0 U8920 ( .CLK(n8987), .C(n9004) );
  CKBD0 U8921 ( .CLK(n8994), .C(n9005) );
  CKBD0 U8922 ( .CLK(n8995), .C(n9006) );
  BUFFD0 U8923 ( .I(n8998), .Z(n9007) );
  BUFFD0 U8924 ( .I(n8881), .Z(n9008) );
  BUFFD0 U8925 ( .I(n8884), .Z(n9009) );
  BUFFD0 U8926 ( .I(n8999), .Z(n9010) );
  BUFFD0 U8927 ( .I(n9000), .Z(n9011) );
  BUFFD0 U8928 ( .I(n9002), .Z(n9012) );
  BUFFD0 U8929 ( .I(n8977), .Z(n9013) );
  BUFFD0 U8930 ( .I(n9003), .Z(n9014) );
  BUFFD0 U8931 ( .I(n9004), .Z(n9015) );
  BUFFD0 U8932 ( .I(n9005), .Z(n9016) );
  BUFFD0 U8933 ( .I(n9006), .Z(n9017) );
  INR2XD0 U8934 ( .A1(n9026), .B1(n9127), .ZN(n97) );
  BUFFD0 U8935 ( .I(n9019), .Z(n9018) );
  BUFFD0 U8936 ( .I(n97), .Z(n9019) );
  CKBD0 U8937 ( .CLK(ParValidTimer[1]), .C(n9020) );
  BUFFD0 U8938 ( .I(n98), .Z(n9021) );
  BUFFD0 U8939 ( .I(n9023), .Z(n9022) );
  BUFFD0 U8940 ( .I(n8), .Z(n9023) );
  BUFFD1 U8941 ( .I(n9159), .Z(n9160) );
  BUFFD1 U8942 ( .I(n9161), .Z(n9159) );
  BUFFD1 U8943 ( .I(n9162), .Z(n9158) );
  BUFFD1 U8944 ( .I(n9162), .Z(n9157) );
  BUFFD1 U8945 ( .I(n9163), .Z(n9161) );
  BUFFD1 U8946 ( .I(n9163), .Z(n9162) );
  BUFFD1 U8947 ( .I(n9164), .Z(n9163) );
  INVD1 U8948 ( .I(Reset), .ZN(n9164) );
  INVD1 U8949 ( .I(n13), .ZN(n9125) );
  BUFFD1 U8950 ( .I(n9130), .Z(n9141) );
  BUFFD1 U8951 ( .I(n9130), .Z(n9142) );
  BUFFD1 U8952 ( .I(n9131), .Z(n9143) );
  BUFFD1 U8953 ( .I(n9131), .Z(n9144) );
  BUFFD1 U8954 ( .I(n9132), .Z(n9145) );
  BUFFD1 U8955 ( .I(n9132), .Z(n9146) );
  BUFFD1 U8956 ( .I(n9133), .Z(n9147) );
  BUFFD1 U8957 ( .I(n9133), .Z(n9148) );
  BUFFD1 U8958 ( .I(n9134), .Z(n9149) );
  BUFFD1 U8959 ( .I(n9134), .Z(n9150) );
  BUFFD1 U8960 ( .I(n9135), .Z(n9151) );
  BUFFD1 U8961 ( .I(n9135), .Z(n9152) );
  BUFFD1 U8962 ( .I(n9136), .Z(n9153) );
  BUFFD1 U8963 ( .I(n9136), .Z(n9154) );
  BUFFD1 U8964 ( .I(n9137), .Z(n9155) );
  BUFFD1 U8965 ( .I(n9137), .Z(n9156) );
  INVD1 U8966 ( .I(n231), .ZN(n9127) );
  INVD1 U8967 ( .I(n231), .ZN(n9128) );
  INVD1 U8968 ( .I(n231), .ZN(n9129) );
  BUFFD1 U8969 ( .I(n13), .Z(n9126) );
  BUFFD1 U8970 ( .I(n9139), .Z(n9132) );
  BUFFD1 U8971 ( .I(n9139), .Z(n9133) );
  BUFFD1 U8972 ( .I(n9139), .Z(n9134) );
  BUFFD1 U8973 ( .I(n9138), .Z(n9135) );
  BUFFD1 U8974 ( .I(n9138), .Z(n9136) );
  BUFFD1 U8975 ( .I(n9138), .Z(n9137) );
  BUFFD1 U8976 ( .I(n9140), .Z(n9130) );
  BUFFD1 U8977 ( .I(n9140), .Z(n9131) );
  IND2D1 U8978 ( .A1(n14), .B1(n15), .ZN(n13) );
  BUFFD1 U8979 ( .I(SerClock), .Z(n9139) );
  BUFFD1 U8980 ( .I(SerClock), .Z(n9138) );
  BUFFD1 U8981 ( .I(SerClock), .Z(n9140) );
  NR2D1 U8982 ( .A1(ParClk), .A2(n232), .ZN(n3) );
  NR2D1 U8983 ( .A1(ParClk), .A2(n27), .ZN(N37) );
  NR4D0 U8984 ( .A1(n28), .A2(Count32[2]), .A3(Count32[4]), .A4(Count32[3]), 
        .ZN(n26) );
  AN2D1 U8985 ( .A1(N34), .A2(n2), .Z(N42) );
  AN2D1 U8986 ( .A1(N33), .A2(n2), .Z(N41) );
  AN2D1 U8987 ( .A1(N32), .A2(n2), .Z(N40) );
  AN2D1 U8988 ( .A1(N31), .A2(n2), .Z(N39) );
  INVD1 U8989 ( .I(n9020), .ZN(n7) );
  AO22D0 U8990 ( .A1(n6723), .A2(n9001), .B1(n6588), .B2(n13), .Z(n133) );
  AO22D0 U8991 ( .A1(n6586), .A2(n9001), .B1(n6451), .B2(n13), .Z(n134) );
  AO22D0 U8992 ( .A1(n6449), .A2(n9001), .B1(n6314), .B2(n13), .Z(n135) );
  AO22D0 U8993 ( .A1(n6312), .A2(n9001), .B1(n6177), .B2(n13), .Z(n136) );
  AO22D0 U8994 ( .A1(n6175), .A2(n9001), .B1(n6040), .B2(n13), .Z(n137) );
  AO22D0 U8995 ( .A1(n6038), .A2(n9001), .B1(n5903), .B2(n13), .Z(n138) );
  AO22D0 U8996 ( .A1(n5901), .A2(n9001), .B1(Decoder[6]), .B2(n9126), .Z(n139)
         );
  AO22D0 U8997 ( .A1(n5764), .A2(n9001), .B1(Decoder[7]), .B2(n13), .Z(n140)
         );
  AO22D0 U8998 ( .A1(n5628), .A2(n9125), .B1(Decoder[8]), .B2(n9126), .Z(n141)
         );
  AO22D0 U8999 ( .A1(n5354), .A2(n9125), .B1(Decoder[10]), .B2(n9126), .Z(n143) );
  AO22D0 U9000 ( .A1(n5218), .A2(n9125), .B1(Decoder[11]), .B2(n9126), .Z(n144) );
  AO22D0 U9001 ( .A1(n5082), .A2(n9001), .B1(Decoder[12]), .B2(n9126), .Z(n145) );
  AO22D0 U9002 ( .A1(n4946), .A2(n9125), .B1(Decoder[13]), .B2(n9126), .Z(n146) );
  AO22D0 U9003 ( .A1(n4810), .A2(n9125), .B1(Decoder[14]), .B2(n9126), .Z(n147) );
  AO22D0 U9004 ( .A1(n4674), .A2(n9125), .B1(Decoder[15]), .B2(n9126), .Z(n148) );
  AO22D0 U9005 ( .A1(n4538), .A2(n9125), .B1(Decoder[16]), .B2(n9126), .Z(n149) );
  AO22D0 U9006 ( .A1(n4402), .A2(n9001), .B1(Decoder[17]), .B2(n9126), .Z(n150) );
  AO22D0 U9007 ( .A1(n4266), .A2(n9001), .B1(Decoder[18]), .B2(n9126), .Z(n151) );
  AO22D0 U9008 ( .A1(n4130), .A2(n9001), .B1(Decoder[19]), .B2(n9126), .Z(n152) );
  AO22D0 U9009 ( .A1(n3994), .A2(n9125), .B1(Decoder[20]), .B2(n9126), .Z(n153) );
  AO22D0 U9010 ( .A1(n3858), .A2(n9125), .B1(Decoder[21]), .B2(n9126), .Z(n154) );
  AO22D0 U9011 ( .A1(n3722), .A2(n9125), .B1(Decoder[22]), .B2(n9126), .Z(n155) );
  AO22D0 U9012 ( .A1(n3586), .A2(n9125), .B1(Decoder[23]), .B2(n9126), .Z(n156) );
  AO22D0 U9013 ( .A1(n3450), .A2(n9125), .B1(Decoder[24]), .B2(n13), .Z(n157)
         );
  AO22D0 U9014 ( .A1(n3314), .A2(n9125), .B1(Decoder[25]), .B2(n13), .Z(n158)
         );
  AO22D0 U9015 ( .A1(n3178), .A2(n9125), .B1(Decoder[26]), .B2(n13), .Z(n159)
         );
  AO22D0 U9016 ( .A1(n3042), .A2(n9125), .B1(Decoder[27]), .B2(n13), .Z(n160)
         );
  AO22D0 U9017 ( .A1(n2906), .A2(n9125), .B1(Decoder[28]), .B2(n13), .Z(n161)
         );
  AO22D0 U9018 ( .A1(n2770), .A2(n9001), .B1(Decoder[29]), .B2(n13), .Z(n162)
         );
  AO22D0 U9019 ( .A1(n2634), .A2(n9125), .B1(Decoder[30]), .B2(n13), .Z(n163)
         );
  AO22D0 U9020 ( .A1(n2495), .A2(n9125), .B1(Decoder[31]), .B2(n9126), .Z(n164) );
  OAI31D0 U9021 ( .A1(n6), .A2(n230), .A3(n7), .B(n232), .ZN(n9026) );
  NR2D1 U9022 ( .A1(n11), .A2(n9127), .ZN(n99) );
  NR2D1 U9023 ( .A1(n6729), .A2(n9127), .ZN(n100) );
  NR2D1 U9024 ( .A1(n9127), .A2(n9022), .ZN(n98) );
  XOR2D1 U9025 ( .A1(n230), .A2(n9), .Z(n8) );
  NR2D1 U9026 ( .A1(n7), .A2(n10), .ZN(n9) );
  NR4D0 U9027 ( .A1(n22), .A2(n8286), .A3(n8275), .A4(n8333), .ZN(n21) );
  ND2D1 U9028 ( .A1(n16), .A2(n17), .ZN(n14) );
  NR4D0 U9029 ( .A1(n8916), .A2(n8906), .A3(n8913), .A4(n8910), .ZN(n16) );
  NR4D0 U9030 ( .A1(n8897), .A2(n8882), .A3(n8875), .A4(n8919), .ZN(n17) );
  AN4D1 U9031 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .Z(n15) );
  INR4D0 U9032 ( .A1(n8383), .B1(n25), .B2(n8553), .B3(n8846), .ZN(n18) );
  NR4D0 U9033 ( .A1(n24), .A2(n8550), .A3(n8398), .A4(n8530), .ZN(n19) );
  NR4D0 U9034 ( .A1(n23), .A2(n8343), .A3(n8215), .A4(n8420), .ZN(n20) );
  ND3D1 U9035 ( .A1(n8518), .A2(n8373), .A3(n8680), .ZN(n25) );
  AN2D1 U9036 ( .A1(SerClk), .A2(SerValid), .Z(SerClock) );
endmodule


module SerialRx_0 ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;
  wire   n2;

  PLLTop_3 PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid3_0 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [2:0] ReadAddr;
  output [2:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n1411, n1412, StateClockRaw, StateClock, N46, N47, N48, N49, N63, N64,
         N65, N66, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n115, n121, n122,
         n124, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n140, n141, n142, n143, n144, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n53,
         n70, n71, n91, n114, n116, n117, n118, n119, n120, n123, n125, n126,
         n139, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1410;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [2:0] OldReadAr;
  wire   [2:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n165), .CPN(StateClock), .Q(FullFIFO), .QN(n115) );
  DFND1 EmptyFIFOr_reg ( .D(n8), .CPN(StateClock), .Q(EmptyFIFO) );
  IAO21D1 U6 ( .A1(n39), .A2(n40), .B(Reset), .ZN(n38) );
  MOAI22D1 U7 ( .A1(n142), .A2(n41), .B1(n41), .B2(n1338), .ZN(n129) );
  MOAI22D1 U11 ( .A1(n144), .A2(n42), .B1(n42), .B2(OldWriteAr[0]), .ZN(n133)
         );
  MOAI22D1 U70 ( .A1(n143), .A2(n41), .B1(n41), .B2(n1399), .ZN(n140) );
  DFNCND1 \NextState_reg[0]  ( .D(n285), .CPN(StateClock), .CDN(n1410), .Q(
        NextState[0]), .QN(n124) );
  DFNCND1 \NextState_reg[1]  ( .D(n347), .CPN(StateClock), .CDN(n1410), .Q(
        NextState[1]), .QN(n122) );
  DFNCND1 \NextState_reg[2]  ( .D(n411), .CPN(StateClock), .CDN(n1410), .Q(
        NextState[2]), .QN(n121) );
  DFCNQD1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n1410), 
        .Q(CurState[2]) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n1410), 
        .Q(CurState[1]) );
  EDFCNQD1 \WriteAr_reg[2]  ( .D(n470), .E(n858), .CP(StateClock), .CDN(n1410), 
        .Q(WriteAddr[2]) );
  DFCNQD1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n1410), 
        .Q(CurState[0]) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(n527), .E(n858), .CP(StateClock), .CDN(n1410), 
        .Q(WriteAddr[1]) );
  EDFCND1 \ReadAr_reg[2]  ( .D(n587), .E(n797), .CP(StateClock), .CDN(n1410), 
        .Q(ReadAddr[2]), .QN(n141) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n645), .E(n797), .CP(StateClock), .CDN(n1410), 
        .Q(ReadAddr[1]), .QN(n142) );
  EDFCND1 \ReadAr_reg[0]  ( .D(n699), .E(n797), .CP(StateClock), .CDN(n1410), 
        .Q(ReadAddr[0]), .QN(n143) );
  EDFCND1 \WriteAr_reg[0]  ( .D(n798), .E(n858), .CP(StateClock), .CDN(n1410), 
        .Q(WriteAddr[0]), .QN(n144) );
  DFNCND1 WriteCmdr_reg ( .D(n912), .CPN(StateClock), .CDN(n1410), .Q(n1412), 
        .QN(n85) );
  DFNCND1 ReadCmdr_reg ( .D(n970), .CPN(StateClock), .CDN(n1410), .Q(n1411), 
        .QN(n7) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n1031), .CPN(StateClock), .CDN(n1410), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n1093), .CPN(StateClock), .CDN(n1410), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n1155), .CPN(StateClock), .CDN(n1410), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n1218), .CPN(StateClock), .CDN(n1410), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n1280), .CPN(StateClock), .CDN(n1410), .Q(
        OldReadAr[1]) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n1342), .CPN(StateClock), .CDN(n1410), .Q(
        OldReadAr[0]) );
  AOI21D0 U3 ( .A1(WriteReq), .A2(n40), .B(n105), .ZN(n104) );
  OA21D0 U4 ( .A1(n46), .A2(n414), .B(n47), .Z(n4) );
  BUFFD0 U5 ( .I(n6), .Z(n1) );
  BUFFD0 U8 ( .I(n754), .Z(n2) );
  AN3D8 U9 ( .A1(n894), .A2(n906), .A3(n112), .Z(n5) );
  BUFFD0 U10 ( .I(n5), .Z(n3) );
  INVD1 U12 ( .I(n4), .ZN(n134) );
  INVD1 U13 ( .I(n3), .ZN(N66) );
  AN2D1 U14 ( .A1(n7), .A2(n2), .Z(n6) );
  INVD1 U15 ( .I(n1), .ZN(N48) );
  BUFFD0 U16 ( .I(n11), .Z(n8) );
  BUFFD0 U17 ( .I(n127), .Z(n9) );
  BUFFD0 U18 ( .I(n36), .Z(n10) );
  BUFFD0 U19 ( .I(n12), .Z(n11) );
  BUFFD0 U20 ( .I(n13), .Z(n12) );
  BUFFD0 U21 ( .I(n14), .Z(n13) );
  BUFFD0 U22 ( .I(n15), .Z(n14) );
  BUFFD0 U23 ( .I(n16), .Z(n15) );
  BUFFD0 U24 ( .I(n17), .Z(n16) );
  BUFFD0 U25 ( .I(n18), .Z(n17) );
  BUFFD0 U26 ( .I(n19), .Z(n18) );
  BUFFD0 U27 ( .I(n20), .Z(n19) );
  BUFFD0 U28 ( .I(n21), .Z(n20) );
  BUFFD0 U29 ( .I(n22), .Z(n21) );
  BUFFD0 U30 ( .I(n23), .Z(n22) );
  BUFFD0 U31 ( .I(n24), .Z(n23) );
  BUFFD0 U32 ( .I(n25), .Z(n24) );
  BUFFD0 U33 ( .I(n26), .Z(n25) );
  BUFFD0 U34 ( .I(n27), .Z(n26) );
  BUFFD0 U35 ( .I(n28), .Z(n27) );
  BUFFD0 U36 ( .I(n29), .Z(n28) );
  BUFFD0 U37 ( .I(n30), .Z(n29) );
  BUFFD0 U38 ( .I(n31), .Z(n30) );
  BUFFD0 U39 ( .I(n32), .Z(n31) );
  BUFFD0 U40 ( .I(n33), .Z(n32) );
  BUFFD0 U41 ( .I(n34), .Z(n33) );
  BUFFD0 U42 ( .I(n53), .Z(n34) );
  BUFFD0 U43 ( .I(n70), .Z(n53) );
  BUFFD0 U44 ( .I(n71), .Z(n70) );
  BUFFD0 U45 ( .I(n91), .Z(n71) );
  BUFFD0 U46 ( .I(n114), .Z(n91) );
  BUFFD0 U47 ( .I(n116), .Z(n114) );
  BUFFD0 U48 ( .I(n117), .Z(n116) );
  BUFFD0 U49 ( .I(n118), .Z(n117) );
  BUFFD0 U50 ( .I(n119), .Z(n118) );
  BUFFD0 U51 ( .I(n120), .Z(n119) );
  BUFFD0 U52 ( .I(n123), .Z(n120) );
  BUFFD0 U53 ( .I(n125), .Z(n123) );
  BUFFD0 U54 ( .I(n126), .Z(n125) );
  BUFFD0 U55 ( .I(n139), .Z(n126) );
  BUFFD0 U56 ( .I(n145), .Z(n139) );
  BUFFD0 U57 ( .I(n146), .Z(n145) );
  BUFFD0 U58 ( .I(n147), .Z(n146) );
  BUFFD0 U59 ( .I(n148), .Z(n147) );
  BUFFD0 U60 ( .I(n149), .Z(n148) );
  BUFFD0 U61 ( .I(n150), .Z(n149) );
  BUFFD0 U62 ( .I(n151), .Z(n150) );
  BUFFD0 U63 ( .I(n152), .Z(n151) );
  BUFFD0 U64 ( .I(n153), .Z(n152) );
  BUFFD0 U65 ( .I(n154), .Z(n153) );
  BUFFD0 U66 ( .I(n155), .Z(n154) );
  BUFFD0 U67 ( .I(n156), .Z(n155) );
  BUFFD0 U68 ( .I(n157), .Z(n156) );
  BUFFD0 U69 ( .I(n158), .Z(n157) );
  BUFFD0 U71 ( .I(n159), .Z(n158) );
  BUFFD0 U72 ( .I(n160), .Z(n159) );
  BUFFD0 U73 ( .I(n161), .Z(n160) );
  BUFFD0 U74 ( .I(n162), .Z(n161) );
  BUFFD0 U75 ( .I(n163), .Z(n162) );
  BUFFD0 U76 ( .I(n164), .Z(n163) );
  BUFFD0 U77 ( .I(n9), .Z(n164) );
  BUFFD0 U78 ( .I(n170), .Z(n165) );
  BUFFD0 U79 ( .I(n167), .Z(n166) );
  BUFFD0 U80 ( .I(n168), .Z(n167) );
  BUFFD0 U81 ( .I(n169), .Z(n168) );
  BUFFD0 U82 ( .I(n115), .Z(n169) );
  BUFFD0 U83 ( .I(n171), .Z(n170) );
  BUFFD0 U84 ( .I(n172), .Z(n171) );
  BUFFD0 U85 ( .I(n173), .Z(n172) );
  BUFFD0 U86 ( .I(n174), .Z(n173) );
  BUFFD0 U87 ( .I(n175), .Z(n174) );
  BUFFD0 U88 ( .I(n176), .Z(n175) );
  BUFFD0 U89 ( .I(n177), .Z(n176) );
  BUFFD0 U90 ( .I(n178), .Z(n177) );
  BUFFD0 U91 ( .I(n179), .Z(n178) );
  BUFFD0 U92 ( .I(n180), .Z(n179) );
  BUFFD0 U93 ( .I(n181), .Z(n180) );
  BUFFD0 U94 ( .I(n182), .Z(n181) );
  BUFFD0 U95 ( .I(n183), .Z(n182) );
  BUFFD0 U96 ( .I(n184), .Z(n183) );
  BUFFD0 U97 ( .I(n185), .Z(n184) );
  BUFFD0 U98 ( .I(n186), .Z(n185) );
  BUFFD0 U99 ( .I(n187), .Z(n186) );
  BUFFD0 U100 ( .I(n188), .Z(n187) );
  BUFFD0 U101 ( .I(n189), .Z(n188) );
  BUFFD0 U102 ( .I(n190), .Z(n189) );
  BUFFD0 U103 ( .I(n191), .Z(n190) );
  BUFFD0 U104 ( .I(n192), .Z(n191) );
  BUFFD0 U105 ( .I(n193), .Z(n192) );
  BUFFD0 U106 ( .I(n194), .Z(n193) );
  BUFFD0 U107 ( .I(n195), .Z(n194) );
  BUFFD0 U108 ( .I(n196), .Z(n195) );
  BUFFD0 U109 ( .I(n197), .Z(n196) );
  BUFFD0 U110 ( .I(n198), .Z(n197) );
  BUFFD0 U111 ( .I(n199), .Z(n198) );
  BUFFD0 U112 ( .I(n200), .Z(n199) );
  BUFFD0 U113 ( .I(n201), .Z(n200) );
  BUFFD0 U114 ( .I(n202), .Z(n201) );
  BUFFD0 U115 ( .I(n203), .Z(n202) );
  BUFFD0 U116 ( .I(n204), .Z(n203) );
  BUFFD0 U117 ( .I(n205), .Z(n204) );
  BUFFD0 U118 ( .I(n206), .Z(n205) );
  BUFFD0 U119 ( .I(n207), .Z(n206) );
  BUFFD0 U120 ( .I(n208), .Z(n207) );
  BUFFD0 U121 ( .I(n209), .Z(n208) );
  BUFFD0 U122 ( .I(n210), .Z(n209) );
  BUFFD0 U123 ( .I(n211), .Z(n210) );
  BUFFD0 U124 ( .I(n212), .Z(n211) );
  BUFFD0 U125 ( .I(n213), .Z(n212) );
  BUFFD0 U126 ( .I(n214), .Z(n213) );
  BUFFD0 U127 ( .I(n215), .Z(n214) );
  BUFFD0 U128 ( .I(n216), .Z(n215) );
  BUFFD0 U129 ( .I(n217), .Z(n216) );
  BUFFD0 U130 ( .I(n218), .Z(n217) );
  BUFFD0 U131 ( .I(n219), .Z(n218) );
  BUFFD0 U132 ( .I(n220), .Z(n219) );
  BUFFD0 U133 ( .I(n221), .Z(n220) );
  BUFFD0 U134 ( .I(n222), .Z(n221) );
  BUFFD0 U135 ( .I(n223), .Z(n222) );
  BUFFD0 U136 ( .I(n224), .Z(n223) );
  BUFFD0 U137 ( .I(n225), .Z(n224) );
  BUFFD0 U138 ( .I(n226), .Z(n225) );
  BUFFD0 U139 ( .I(n227), .Z(n226) );
  BUFFD0 U140 ( .I(n128), .Z(n227) );
  BUFFD0 U141 ( .I(n1412), .Z(n228) );
  BUFFD0 U142 ( .I(n228), .Z(n229) );
  BUFFD0 U143 ( .I(n229), .Z(n230) );
  BUFFD0 U144 ( .I(n230), .Z(n231) );
  BUFFD0 U145 ( .I(n231), .Z(n232) );
  BUFFD0 U146 ( .I(n232), .Z(n233) );
  BUFFD0 U147 ( .I(n233), .Z(n234) );
  BUFFD0 U148 ( .I(n234), .Z(n235) );
  BUFFD0 U149 ( .I(n235), .Z(n236) );
  BUFFD0 U150 ( .I(n236), .Z(n237) );
  BUFFD0 U151 ( .I(n237), .Z(n238) );
  BUFFD0 U152 ( .I(n238), .Z(n239) );
  BUFFD0 U153 ( .I(n239), .Z(n240) );
  BUFFD0 U154 ( .I(n240), .Z(n241) );
  BUFFD0 U155 ( .I(n241), .Z(n242) );
  BUFFD0 U156 ( .I(n242), .Z(n243) );
  BUFFD0 U157 ( .I(n243), .Z(n244) );
  BUFFD0 U158 ( .I(n244), .Z(n245) );
  BUFFD0 U159 ( .I(n245), .Z(n246) );
  BUFFD0 U160 ( .I(n246), .Z(n247) );
  BUFFD0 U161 ( .I(n247), .Z(n248) );
  BUFFD0 U162 ( .I(n248), .Z(n249) );
  BUFFD0 U163 ( .I(n249), .Z(n250) );
  BUFFD0 U164 ( .I(n250), .Z(n251) );
  BUFFD0 U165 ( .I(n251), .Z(n252) );
  BUFFD0 U166 ( .I(n252), .Z(n253) );
  BUFFD0 U167 ( .I(n253), .Z(n254) );
  BUFFD0 U168 ( .I(n254), .Z(n255) );
  BUFFD0 U169 ( .I(n255), .Z(n256) );
  BUFFD0 U170 ( .I(n256), .Z(n257) );
  BUFFD0 U171 ( .I(n257), .Z(n258) );
  BUFFD0 U172 ( .I(n258), .Z(n259) );
  BUFFD0 U173 ( .I(n259), .Z(n260) );
  BUFFD0 U174 ( .I(n260), .Z(n261) );
  BUFFD0 U175 ( .I(n261), .Z(n262) );
  BUFFD0 U176 ( .I(n262), .Z(n263) );
  BUFFD0 U177 ( .I(n263), .Z(n264) );
  BUFFD0 U178 ( .I(n264), .Z(n265) );
  BUFFD0 U179 ( .I(n265), .Z(n266) );
  BUFFD0 U180 ( .I(n266), .Z(n267) );
  BUFFD0 U181 ( .I(n267), .Z(n268) );
  BUFFD0 U182 ( .I(n268), .Z(n269) );
  BUFFD0 U183 ( .I(n269), .Z(n270) );
  BUFFD0 U184 ( .I(n270), .Z(n271) );
  BUFFD0 U185 ( .I(n271), .Z(n272) );
  BUFFD0 U186 ( .I(n272), .Z(n273) );
  BUFFD0 U187 ( .I(n273), .Z(n274) );
  BUFFD0 U188 ( .I(n274), .Z(n275) );
  BUFFD0 U189 ( .I(n275), .Z(n276) );
  BUFFD0 U190 ( .I(n276), .Z(n277) );
  BUFFD0 U191 ( .I(n277), .Z(n278) );
  BUFFD0 U192 ( .I(n278), .Z(n279) );
  BUFFD0 U193 ( .I(n279), .Z(n280) );
  BUFFD0 U194 ( .I(n280), .Z(n281) );
  BUFFD0 U195 ( .I(n281), .Z(n282) );
  BUFFD0 U196 ( .I(n282), .Z(n283) );
  CKBD0 U197 ( .CLK(n283), .C(WriteCmd) );
  BUFFD0 U198 ( .I(n288), .Z(n285) );
  BUFFD0 U199 ( .I(n137), .Z(n286) );
  BUFFD0 U200 ( .I(n286), .Z(n287) );
  BUFFD0 U201 ( .I(n289), .Z(n288) );
  BUFFD0 U202 ( .I(n290), .Z(n289) );
  BUFFD0 U203 ( .I(n297), .Z(n290) );
  BUFFD0 U204 ( .I(n292), .Z(n291) );
  BUFFD0 U205 ( .I(n293), .Z(n292) );
  BUFFD0 U206 ( .I(n294), .Z(n293) );
  BUFFD0 U207 ( .I(n295), .Z(n294) );
  BUFFD0 U208 ( .I(n296), .Z(n295) );
  BUFFD0 U209 ( .I(n124), .Z(n296) );
  BUFFD0 U210 ( .I(n298), .Z(n297) );
  BUFFD0 U211 ( .I(n299), .Z(n298) );
  BUFFD0 U212 ( .I(n300), .Z(n299) );
  BUFFD0 U213 ( .I(n301), .Z(n300) );
  BUFFD0 U214 ( .I(n302), .Z(n301) );
  BUFFD0 U215 ( .I(n303), .Z(n302) );
  BUFFD0 U216 ( .I(n304), .Z(n303) );
  BUFFD0 U217 ( .I(n305), .Z(n304) );
  BUFFD0 U218 ( .I(n306), .Z(n305) );
  BUFFD0 U219 ( .I(n307), .Z(n306) );
  BUFFD0 U220 ( .I(n308), .Z(n307) );
  BUFFD0 U221 ( .I(n309), .Z(n308) );
  BUFFD0 U222 ( .I(n310), .Z(n309) );
  BUFFD0 U223 ( .I(n311), .Z(n310) );
  BUFFD0 U224 ( .I(n312), .Z(n311) );
  BUFFD0 U225 ( .I(n313), .Z(n312) );
  BUFFD0 U226 ( .I(n314), .Z(n313) );
  BUFFD0 U227 ( .I(n315), .Z(n314) );
  BUFFD0 U228 ( .I(n316), .Z(n315) );
  BUFFD0 U229 ( .I(n317), .Z(n316) );
  BUFFD0 U230 ( .I(n318), .Z(n317) );
  BUFFD0 U231 ( .I(n319), .Z(n318) );
  BUFFD0 U232 ( .I(n320), .Z(n319) );
  BUFFD0 U233 ( .I(n321), .Z(n320) );
  BUFFD0 U234 ( .I(n322), .Z(n321) );
  BUFFD0 U235 ( .I(n323), .Z(n322) );
  BUFFD0 U236 ( .I(n324), .Z(n323) );
  BUFFD0 U237 ( .I(n325), .Z(n324) );
  BUFFD0 U238 ( .I(n326), .Z(n325) );
  BUFFD0 U239 ( .I(n327), .Z(n326) );
  BUFFD0 U240 ( .I(n328), .Z(n327) );
  BUFFD0 U241 ( .I(n329), .Z(n328) );
  BUFFD0 U242 ( .I(n330), .Z(n329) );
  BUFFD0 U243 ( .I(n331), .Z(n330) );
  BUFFD0 U244 ( .I(n332), .Z(n331) );
  BUFFD0 U245 ( .I(n333), .Z(n332) );
  BUFFD0 U246 ( .I(n334), .Z(n333) );
  BUFFD0 U247 ( .I(n335), .Z(n334) );
  BUFFD0 U248 ( .I(n336), .Z(n335) );
  BUFFD0 U249 ( .I(n337), .Z(n336) );
  BUFFD0 U250 ( .I(n338), .Z(n337) );
  BUFFD0 U251 ( .I(n339), .Z(n338) );
  BUFFD0 U252 ( .I(n340), .Z(n339) );
  BUFFD0 U253 ( .I(n341), .Z(n340) );
  BUFFD0 U254 ( .I(n342), .Z(n341) );
  BUFFD0 U255 ( .I(n343), .Z(n342) );
  BUFFD0 U256 ( .I(n344), .Z(n343) );
  BUFFD0 U257 ( .I(n345), .Z(n344) );
  BUFFD0 U258 ( .I(n346), .Z(n345) );
  BUFFD0 U259 ( .I(n287), .Z(n346) );
  BUFFD0 U260 ( .I(n350), .Z(n347) );
  BUFFD0 U261 ( .I(n135), .Z(n348) );
  BUFFD0 U262 ( .I(n348), .Z(n349) );
  BUFFD0 U263 ( .I(n351), .Z(n350) );
  BUFFD0 U264 ( .I(n358), .Z(n351) );
  BUFFD0 U265 ( .I(n353), .Z(n352) );
  OAI211D0 U266 ( .A1(CurState[1]), .A2(n79), .B(n83), .C(n104), .ZN(n46) );
  BUFFD0 U267 ( .I(n354), .Z(n353) );
  BUFFD0 U268 ( .I(n355), .Z(n354) );
  BUFFD0 U269 ( .I(n356), .Z(n355) );
  BUFFD0 U270 ( .I(n357), .Z(n356) );
  BUFFD0 U271 ( .I(n122), .Z(n357) );
  BUFFD0 U272 ( .I(n359), .Z(n358) );
  BUFFD0 U273 ( .I(n360), .Z(n359) );
  BUFFD0 U274 ( .I(n361), .Z(n360) );
  BUFFD0 U275 ( .I(n362), .Z(n361) );
  BUFFD0 U276 ( .I(n363), .Z(n362) );
  BUFFD0 U277 ( .I(n364), .Z(n363) );
  BUFFD0 U278 ( .I(n365), .Z(n364) );
  BUFFD0 U279 ( .I(n366), .Z(n365) );
  BUFFD0 U280 ( .I(n367), .Z(n366) );
  BUFFD0 U281 ( .I(n368), .Z(n367) );
  BUFFD0 U282 ( .I(n369), .Z(n368) );
  BUFFD0 U283 ( .I(n370), .Z(n369) );
  BUFFD0 U284 ( .I(n371), .Z(n370) );
  BUFFD0 U285 ( .I(n372), .Z(n371) );
  BUFFD0 U286 ( .I(n373), .Z(n372) );
  BUFFD0 U287 ( .I(n374), .Z(n373) );
  BUFFD0 U288 ( .I(n375), .Z(n374) );
  BUFFD0 U289 ( .I(n376), .Z(n375) );
  BUFFD0 U290 ( .I(n377), .Z(n376) );
  BUFFD0 U291 ( .I(n378), .Z(n377) );
  BUFFD0 U292 ( .I(n379), .Z(n378) );
  BUFFD0 U293 ( .I(n380), .Z(n379) );
  BUFFD0 U294 ( .I(n381), .Z(n380) );
  BUFFD0 U295 ( .I(n382), .Z(n381) );
  BUFFD0 U296 ( .I(n383), .Z(n382) );
  BUFFD0 U297 ( .I(n384), .Z(n383) );
  BUFFD0 U298 ( .I(n385), .Z(n384) );
  BUFFD0 U299 ( .I(n386), .Z(n385) );
  BUFFD0 U300 ( .I(n387), .Z(n386) );
  BUFFD0 U301 ( .I(n388), .Z(n387) );
  BUFFD0 U302 ( .I(n389), .Z(n388) );
  BUFFD0 U303 ( .I(n390), .Z(n389) );
  BUFFD0 U304 ( .I(n391), .Z(n390) );
  BUFFD0 U305 ( .I(n392), .Z(n391) );
  BUFFD0 U306 ( .I(n393), .Z(n392) );
  BUFFD0 U307 ( .I(n394), .Z(n393) );
  BUFFD0 U308 ( .I(n395), .Z(n394) );
  BUFFD0 U309 ( .I(n396), .Z(n395) );
  BUFFD0 U310 ( .I(n397), .Z(n396) );
  BUFFD0 U311 ( .I(n398), .Z(n397) );
  BUFFD0 U312 ( .I(n399), .Z(n398) );
  BUFFD0 U313 ( .I(n400), .Z(n399) );
  BUFFD0 U314 ( .I(n401), .Z(n400) );
  BUFFD0 U315 ( .I(n402), .Z(n401) );
  BUFFD0 U316 ( .I(n403), .Z(n402) );
  BUFFD0 U317 ( .I(n404), .Z(n403) );
  BUFFD0 U318 ( .I(n405), .Z(n404) );
  BUFFD0 U319 ( .I(n406), .Z(n405) );
  BUFFD0 U320 ( .I(n407), .Z(n406) );
  BUFFD0 U321 ( .I(n408), .Z(n407) );
  BUFFD0 U322 ( .I(n349), .Z(n408) );
  BUFFD0 U323 ( .I(n134), .Z(n409) );
  BUFFD0 U324 ( .I(n409), .Z(n410) );
  BUFFD0 U325 ( .I(n412), .Z(n411) );
  BUFFD0 U326 ( .I(n413), .Z(n412) );
  BUFFD0 U327 ( .I(n418), .Z(n413) );
  BUFFD0 U328 ( .I(n415), .Z(n414) );
  BUFFD0 U329 ( .I(n416), .Z(n415) );
  BUFFD0 U330 ( .I(n417), .Z(n416) );
  BUFFD0 U331 ( .I(n121), .Z(n417) );
  BUFFD0 U332 ( .I(n419), .Z(n418) );
  BUFFD0 U333 ( .I(n420), .Z(n419) );
  BUFFD0 U334 ( .I(n421), .Z(n420) );
  BUFFD0 U335 ( .I(n422), .Z(n421) );
  BUFFD0 U336 ( .I(n423), .Z(n422) );
  BUFFD0 U337 ( .I(n424), .Z(n423) );
  BUFFD0 U338 ( .I(n425), .Z(n424) );
  BUFFD0 U339 ( .I(n426), .Z(n425) );
  BUFFD0 U340 ( .I(n427), .Z(n426) );
  BUFFD0 U341 ( .I(n428), .Z(n427) );
  BUFFD0 U342 ( .I(n429), .Z(n428) );
  BUFFD0 U343 ( .I(n430), .Z(n429) );
  BUFFD0 U344 ( .I(n431), .Z(n430) );
  BUFFD0 U345 ( .I(n432), .Z(n431) );
  BUFFD0 U346 ( .I(n433), .Z(n432) );
  BUFFD0 U347 ( .I(n434), .Z(n433) );
  BUFFD0 U348 ( .I(n435), .Z(n434) );
  BUFFD0 U349 ( .I(n436), .Z(n435) );
  BUFFD0 U350 ( .I(n437), .Z(n436) );
  BUFFD0 U351 ( .I(n438), .Z(n437) );
  BUFFD0 U352 ( .I(n439), .Z(n438) );
  BUFFD0 U353 ( .I(n440), .Z(n439) );
  BUFFD0 U354 ( .I(n441), .Z(n440) );
  BUFFD0 U355 ( .I(n442), .Z(n441) );
  BUFFD0 U356 ( .I(n443), .Z(n442) );
  BUFFD0 U357 ( .I(n444), .Z(n443) );
  BUFFD0 U358 ( .I(n445), .Z(n444) );
  BUFFD0 U359 ( .I(n446), .Z(n445) );
  BUFFD0 U360 ( .I(n447), .Z(n446) );
  BUFFD0 U361 ( .I(n448), .Z(n447) );
  BUFFD0 U362 ( .I(n449), .Z(n448) );
  BUFFD0 U363 ( .I(n450), .Z(n449) );
  BUFFD0 U364 ( .I(n451), .Z(n450) );
  BUFFD0 U365 ( .I(n452), .Z(n451) );
  BUFFD0 U366 ( .I(n453), .Z(n452) );
  BUFFD0 U367 ( .I(n454), .Z(n453) );
  BUFFD0 U368 ( .I(n455), .Z(n454) );
  BUFFD0 U369 ( .I(n456), .Z(n455) );
  BUFFD0 U370 ( .I(n457), .Z(n456) );
  BUFFD0 U371 ( .I(n458), .Z(n457) );
  BUFFD0 U372 ( .I(n459), .Z(n458) );
  BUFFD0 U373 ( .I(n460), .Z(n459) );
  BUFFD0 U374 ( .I(n461), .Z(n460) );
  BUFFD0 U375 ( .I(n462), .Z(n461) );
  BUFFD0 U376 ( .I(n463), .Z(n462) );
  BUFFD0 U377 ( .I(n464), .Z(n463) );
  BUFFD0 U378 ( .I(n465), .Z(n464) );
  BUFFD0 U379 ( .I(n466), .Z(n465) );
  BUFFD0 U380 ( .I(n467), .Z(n466) );
  BUFFD0 U381 ( .I(n468), .Z(n467) );
  BUFFD0 U382 ( .I(n469), .Z(n468) );
  BUFFD0 U383 ( .I(n410), .Z(n469) );
  BUFFD0 U384 ( .I(n474), .Z(n470) );
  BUFFD0 U385 ( .I(N65), .Z(n471) );
  BUFFD0 U386 ( .I(n471), .Z(n472) );
  BUFFD0 U387 ( .I(n472), .Z(n473) );
  BUFFD0 U388 ( .I(n475), .Z(n474) );
  BUFFD0 U389 ( .I(n476), .Z(n475) );
  BUFFD0 U390 ( .I(n477), .Z(n476) );
  BUFFD0 U391 ( .I(n478), .Z(n477) );
  BUFFD0 U392 ( .I(n479), .Z(n478) );
  BUFFD0 U393 ( .I(n480), .Z(n479) );
  BUFFD0 U394 ( .I(n481), .Z(n480) );
  BUFFD0 U395 ( .I(n482), .Z(n481) );
  BUFFD0 U396 ( .I(n483), .Z(n482) );
  BUFFD0 U397 ( .I(n484), .Z(n483) );
  BUFFD0 U398 ( .I(n485), .Z(n484) );
  BUFFD0 U399 ( .I(n486), .Z(n485) );
  BUFFD0 U400 ( .I(n487), .Z(n486) );
  BUFFD0 U401 ( .I(n488), .Z(n487) );
  BUFFD0 U402 ( .I(n489), .Z(n488) );
  BUFFD0 U403 ( .I(n490), .Z(n489) );
  BUFFD0 U404 ( .I(n491), .Z(n490) );
  BUFFD0 U405 ( .I(n492), .Z(n491) );
  BUFFD0 U406 ( .I(n493), .Z(n492) );
  BUFFD0 U407 ( .I(n494), .Z(n493) );
  BUFFD0 U408 ( .I(n495), .Z(n494) );
  BUFFD0 U409 ( .I(n496), .Z(n495) );
  BUFFD0 U410 ( .I(n497), .Z(n496) );
  BUFFD0 U411 ( .I(n498), .Z(n497) );
  BUFFD0 U412 ( .I(n499), .Z(n498) );
  BUFFD0 U413 ( .I(n500), .Z(n499) );
  BUFFD0 U414 ( .I(n501), .Z(n500) );
  BUFFD0 U415 ( .I(n502), .Z(n501) );
  BUFFD0 U416 ( .I(n503), .Z(n502) );
  BUFFD0 U417 ( .I(n504), .Z(n503) );
  BUFFD0 U418 ( .I(n505), .Z(n504) );
  BUFFD0 U419 ( .I(n506), .Z(n505) );
  BUFFD0 U420 ( .I(n507), .Z(n506) );
  BUFFD0 U421 ( .I(n508), .Z(n507) );
  BUFFD0 U422 ( .I(n509), .Z(n508) );
  BUFFD0 U423 ( .I(n510), .Z(n509) );
  BUFFD0 U424 ( .I(n511), .Z(n510) );
  BUFFD0 U425 ( .I(n512), .Z(n511) );
  BUFFD0 U426 ( .I(n513), .Z(n512) );
  BUFFD0 U427 ( .I(n514), .Z(n513) );
  BUFFD0 U428 ( .I(n515), .Z(n514) );
  BUFFD0 U429 ( .I(n516), .Z(n515) );
  BUFFD0 U430 ( .I(n517), .Z(n516) );
  BUFFD0 U431 ( .I(n518), .Z(n517) );
  BUFFD0 U432 ( .I(n519), .Z(n518) );
  BUFFD0 U433 ( .I(n520), .Z(n519) );
  BUFFD0 U434 ( .I(n521), .Z(n520) );
  BUFFD0 U435 ( .I(n522), .Z(n521) );
  BUFFD0 U436 ( .I(n523), .Z(n522) );
  BUFFD0 U437 ( .I(n524), .Z(n523) );
  BUFFD0 U438 ( .I(n525), .Z(n524) );
  BUFFD0 U439 ( .I(n473), .Z(n525) );
  BUFFD0 U440 ( .I(n141), .Z(n526) );
  BUFFD0 U441 ( .I(n532), .Z(n527) );
  BUFFD0 U442 ( .I(N64), .Z(n528) );
  BUFFD0 U443 ( .I(n528), .Z(n529) );
  BUFFD0 U444 ( .I(n529), .Z(n530) );
  BUFFD0 U445 ( .I(n530), .Z(n531) );
  BUFFD0 U446 ( .I(n533), .Z(n532) );
  BUFFD0 U447 ( .I(n534), .Z(n533) );
  BUFFD0 U448 ( .I(n535), .Z(n534) );
  BUFFD0 U449 ( .I(n536), .Z(n535) );
  BUFFD0 U450 ( .I(n537), .Z(n536) );
  BUFFD0 U451 ( .I(n538), .Z(n537) );
  BUFFD0 U452 ( .I(n539), .Z(n538) );
  BUFFD0 U453 ( .I(n540), .Z(n539) );
  BUFFD0 U454 ( .I(n541), .Z(n540) );
  BUFFD0 U455 ( .I(n542), .Z(n541) );
  BUFFD0 U456 ( .I(n543), .Z(n542) );
  BUFFD0 U457 ( .I(n544), .Z(n543) );
  BUFFD0 U458 ( .I(n545), .Z(n544) );
  BUFFD0 U459 ( .I(n546), .Z(n545) );
  BUFFD0 U460 ( .I(n547), .Z(n546) );
  BUFFD0 U461 ( .I(n548), .Z(n547) );
  BUFFD0 U462 ( .I(n549), .Z(n548) );
  BUFFD0 U463 ( .I(n550), .Z(n549) );
  BUFFD0 U464 ( .I(n551), .Z(n550) );
  BUFFD0 U465 ( .I(n552), .Z(n551) );
  BUFFD0 U466 ( .I(n553), .Z(n552) );
  BUFFD0 U467 ( .I(n554), .Z(n553) );
  BUFFD0 U468 ( .I(n555), .Z(n554) );
  BUFFD0 U469 ( .I(n556), .Z(n555) );
  BUFFD0 U470 ( .I(n557), .Z(n556) );
  BUFFD0 U471 ( .I(n558), .Z(n557) );
  BUFFD0 U472 ( .I(n559), .Z(n558) );
  BUFFD0 U473 ( .I(n560), .Z(n559) );
  BUFFD0 U474 ( .I(n561), .Z(n560) );
  BUFFD0 U475 ( .I(n562), .Z(n561) );
  BUFFD0 U476 ( .I(n563), .Z(n562) );
  BUFFD0 U477 ( .I(n564), .Z(n563) );
  BUFFD0 U478 ( .I(n565), .Z(n564) );
  BUFFD0 U479 ( .I(n566), .Z(n565) );
  BUFFD0 U480 ( .I(n567), .Z(n566) );
  BUFFD0 U481 ( .I(n568), .Z(n567) );
  BUFFD0 U482 ( .I(n569), .Z(n568) );
  BUFFD0 U483 ( .I(n570), .Z(n569) );
  BUFFD0 U484 ( .I(n571), .Z(n570) );
  BUFFD0 U485 ( .I(n572), .Z(n571) );
  BUFFD0 U486 ( .I(n573), .Z(n572) );
  BUFFD0 U487 ( .I(n574), .Z(n573) );
  BUFFD0 U488 ( .I(n575), .Z(n574) );
  BUFFD0 U489 ( .I(n576), .Z(n575) );
  BUFFD0 U490 ( .I(n577), .Z(n576) );
  BUFFD0 U491 ( .I(n578), .Z(n577) );
  BUFFD0 U492 ( .I(n579), .Z(n578) );
  BUFFD0 U493 ( .I(n580), .Z(n579) );
  BUFFD0 U494 ( .I(n581), .Z(n580) );
  BUFFD0 U495 ( .I(n582), .Z(n581) );
  BUFFD0 U496 ( .I(n583), .Z(n582) );
  BUFFD0 U497 ( .I(n531), .Z(n583) );
  CKBD0 U498 ( .CLK(WriteAddr[0]), .C(n857) );
  BUFFD0 U499 ( .I(n142), .Z(n584) );
  OAI21D0 U500 ( .A1(WriteAddr[1]), .A2(n857), .B(n81), .ZN(n100) );
  BUFFD0 U501 ( .I(n1411), .Z(n585) );
  BUFFD0 U502 ( .I(n585), .Z(n586) );
  BUFFD0 U503 ( .I(n588), .Z(n587) );
  BUFFD0 U504 ( .I(n589), .Z(n588) );
  BUFFD0 U505 ( .I(n590), .Z(n589) );
  BUFFD0 U506 ( .I(n591), .Z(n590) );
  BUFFD0 U507 ( .I(n592), .Z(n591) );
  BUFFD0 U508 ( .I(n593), .Z(n592) );
  BUFFD0 U509 ( .I(n595), .Z(n593) );
  BUFFD0 U510 ( .I(n596), .Z(n594) );
  BUFFD0 U511 ( .I(n597), .Z(n595) );
  BUFFD0 U512 ( .I(n598), .Z(n596) );
  BUFFD0 U513 ( .I(n599), .Z(n597) );
  BUFFD0 U514 ( .I(n600), .Z(n598) );
  BUFFD0 U515 ( .I(n601), .Z(n599) );
  BUFFD0 U516 ( .I(n602), .Z(n600) );
  BUFFD0 U517 ( .I(n603), .Z(n601) );
  BUFFD0 U518 ( .I(n604), .Z(n602) );
  BUFFD0 U519 ( .I(n605), .Z(n603) );
  BUFFD0 U520 ( .I(n606), .Z(n604) );
  BUFFD0 U521 ( .I(n607), .Z(n605) );
  BUFFD0 U522 ( .I(n608), .Z(n606) );
  BUFFD0 U523 ( .I(n609), .Z(n607) );
  BUFFD0 U524 ( .I(n610), .Z(n608) );
  BUFFD0 U525 ( .I(n611), .Z(n609) );
  BUFFD0 U526 ( .I(n612), .Z(n610) );
  BUFFD0 U527 ( .I(n613), .Z(n611) );
  BUFFD0 U528 ( .I(n614), .Z(n612) );
  BUFFD0 U529 ( .I(n615), .Z(n613) );
  BUFFD0 U530 ( .I(n616), .Z(n614) );
  BUFFD0 U531 ( .I(n617), .Z(n615) );
  BUFFD0 U532 ( .I(n618), .Z(n616) );
  BUFFD0 U533 ( .I(n619), .Z(n617) );
  BUFFD0 U534 ( .I(n620), .Z(n618) );
  BUFFD0 U535 ( .I(N49), .Z(n619) );
  BUFFD0 U536 ( .I(n621), .Z(n620) );
  BUFFD0 U537 ( .I(n622), .Z(n621) );
  BUFFD0 U538 ( .I(n623), .Z(n622) );
  BUFFD0 U539 ( .I(n624), .Z(n623) );
  BUFFD0 U540 ( .I(n625), .Z(n624) );
  BUFFD0 U541 ( .I(n626), .Z(n625) );
  BUFFD0 U542 ( .I(n627), .Z(n626) );
  BUFFD0 U543 ( .I(n628), .Z(n627) );
  BUFFD0 U544 ( .I(n629), .Z(n628) );
  BUFFD0 U545 ( .I(n630), .Z(n629) );
  BUFFD0 U546 ( .I(n631), .Z(n630) );
  BUFFD0 U547 ( .I(n632), .Z(n631) );
  BUFFD0 U548 ( .I(n633), .Z(n632) );
  BUFFD0 U549 ( .I(n634), .Z(n633) );
  BUFFD0 U550 ( .I(n635), .Z(n634) );
  BUFFD0 U551 ( .I(n636), .Z(n635) );
  BUFFD0 U552 ( .I(n637), .Z(n636) );
  BUFFD0 U553 ( .I(n638), .Z(n637) );
  BUFFD0 U554 ( .I(n639), .Z(n638) );
  BUFFD0 U555 ( .I(n640), .Z(n639) );
  BUFFD0 U556 ( .I(n643), .Z(n640) );
  BUFFD0 U557 ( .I(n584), .Z(n641) );
  BUFFD0 U558 ( .I(n644), .Z(n642) );
  BUFFD0 U559 ( .I(n99), .Z(n643) );
  BUFFD0 U560 ( .I(n526), .Z(n644) );
  BUFFD0 U561 ( .I(n646), .Z(n645) );
  BUFFD0 U562 ( .I(n647), .Z(n646) );
  BUFFD0 U563 ( .I(n648), .Z(n647) );
  BUFFD0 U564 ( .I(n649), .Z(n648) );
  BUFFD0 U565 ( .I(n651), .Z(n649) );
  BUFFD0 U566 ( .I(n652), .Z(n650) );
  BUFFD0 U567 ( .I(n653), .Z(n651) );
  BUFFD0 U568 ( .I(n654), .Z(n652) );
  BUFFD0 U569 ( .I(n655), .Z(n653) );
  BUFFD0 U570 ( .I(n656), .Z(n654) );
  BUFFD0 U571 ( .I(n657), .Z(n655) );
  BUFFD0 U572 ( .I(n658), .Z(n656) );
  BUFFD0 U573 ( .I(n659), .Z(n657) );
  BUFFD0 U574 ( .I(n661), .Z(n658) );
  BUFFD0 U575 ( .I(n660), .Z(n659) );
  BUFFD0 U576 ( .I(n662), .Z(n660) );
  BUFFD0 U577 ( .I(n663), .Z(n661) );
  BUFFD0 U578 ( .I(n664), .Z(n662) );
  BUFFD0 U579 ( .I(n665), .Z(n663) );
  BUFFD0 U580 ( .I(n666), .Z(n664) );
  BUFFD0 U581 ( .I(n667), .Z(n665) );
  BUFFD0 U582 ( .I(n668), .Z(n666) );
  BUFFD0 U583 ( .I(n669), .Z(n667) );
  BUFFD0 U584 ( .I(n670), .Z(n668) );
  BUFFD0 U585 ( .I(n671), .Z(n669) );
  BUFFD0 U586 ( .I(n672), .Z(n670) );
  BUFFD0 U587 ( .I(n673), .Z(n671) );
  BUFFD0 U588 ( .I(n674), .Z(n672) );
  BUFFD0 U589 ( .I(n675), .Z(n673) );
  BUFFD0 U590 ( .I(n676), .Z(n674) );
  BUFFD0 U591 ( .I(n677), .Z(n675) );
  BUFFD0 U592 ( .I(n678), .Z(n676) );
  BUFFD0 U593 ( .I(n679), .Z(n677) );
  BUFFD0 U594 ( .I(N47), .Z(n678) );
  BUFFD0 U595 ( .I(n680), .Z(n679) );
  BUFFD0 U596 ( .I(n681), .Z(n680) );
  BUFFD0 U597 ( .I(n682), .Z(n681) );
  BUFFD0 U598 ( .I(n683), .Z(n682) );
  BUFFD0 U599 ( .I(n684), .Z(n683) );
  BUFFD0 U600 ( .I(n685), .Z(n684) );
  BUFFD0 U601 ( .I(n686), .Z(n685) );
  BUFFD0 U602 ( .I(n687), .Z(n686) );
  BUFFD0 U603 ( .I(n688), .Z(n687) );
  BUFFD0 U604 ( .I(n689), .Z(n688) );
  BUFFD0 U605 ( .I(n690), .Z(n689) );
  BUFFD0 U606 ( .I(n691), .Z(n690) );
  BUFFD0 U607 ( .I(n692), .Z(n691) );
  BUFFD0 U608 ( .I(n693), .Z(n692) );
  BUFFD0 U609 ( .I(n694), .Z(n693) );
  BUFFD0 U610 ( .I(n695), .Z(n694) );
  BUFFD0 U611 ( .I(n696), .Z(n695) );
  BUFFD0 U612 ( .I(n697), .Z(n696) );
  BUFFD0 U613 ( .I(n698), .Z(n697) );
  BUFFD0 U614 ( .I(n113), .Z(n698) );
  XNR2D0 U615 ( .A1(n700), .A2(ReadAddr[1]), .ZN(n113) );
  BUFFD0 U616 ( .I(n701), .Z(n699) );
  BUFFD0 U617 ( .I(n702), .Z(n700) );
  BUFFD0 U618 ( .I(n703), .Z(n701) );
  BUFFD0 U619 ( .I(n704), .Z(n702) );
  BUFFD0 U620 ( .I(n705), .Z(n703) );
  BUFFD0 U621 ( .I(n706), .Z(n704) );
  BUFFD0 U622 ( .I(n707), .Z(n705) );
  BUFFD0 U623 ( .I(n708), .Z(n706) );
  BUFFD0 U624 ( .I(n709), .Z(n707) );
  BUFFD0 U625 ( .I(n710), .Z(n708) );
  BUFFD0 U626 ( .I(n711), .Z(n709) );
  BUFFD0 U627 ( .I(n712), .Z(n710) );
  BUFFD0 U628 ( .I(n713), .Z(n711) );
  BUFFD0 U629 ( .I(n714), .Z(n712) );
  BUFFD0 U630 ( .I(n715), .Z(n713) );
  BUFFD0 U631 ( .I(n716), .Z(n714) );
  BUFFD0 U632 ( .I(n717), .Z(n715) );
  BUFFD0 U633 ( .I(n718), .Z(n716) );
  BUFFD0 U634 ( .I(n719), .Z(n717) );
  BUFFD0 U635 ( .I(n720), .Z(n718) );
  BUFFD0 U636 ( .I(n721), .Z(n719) );
  BUFFD0 U637 ( .I(n722), .Z(n720) );
  BUFFD0 U638 ( .I(n723), .Z(n721) );
  BUFFD0 U639 ( .I(n724), .Z(n722) );
  BUFFD0 U640 ( .I(n725), .Z(n723) );
  BUFFD0 U641 ( .I(n726), .Z(n724) );
  BUFFD0 U642 ( .I(n727), .Z(n725) );
  BUFFD0 U643 ( .I(n728), .Z(n726) );
  BUFFD0 U644 ( .I(n729), .Z(n727) );
  BUFFD0 U645 ( .I(n730), .Z(n728) );
  BUFFD0 U646 ( .I(n731), .Z(n729) );
  BUFFD0 U647 ( .I(n732), .Z(n730) );
  BUFFD0 U648 ( .I(n733), .Z(n731) );
  BUFFD0 U649 ( .I(n734), .Z(n732) );
  BUFFD0 U650 ( .I(n735), .Z(n733) );
  BUFFD0 U651 ( .I(n736), .Z(n734) );
  BUFFD0 U652 ( .I(n737), .Z(n735) );
  BUFFD0 U653 ( .I(n738), .Z(n736) );
  BUFFD0 U654 ( .I(n739), .Z(n737) );
  BUFFD0 U655 ( .I(n740), .Z(n738) );
  BUFFD0 U656 ( .I(N46), .Z(n739) );
  BUFFD0 U657 ( .I(n741), .Z(n740) );
  BUFFD0 U658 ( .I(n742), .Z(n741) );
  BUFFD0 U659 ( .I(n743), .Z(n742) );
  BUFFD0 U660 ( .I(n744), .Z(n743) );
  BUFFD0 U661 ( .I(n745), .Z(n744) );
  BUFFD0 U662 ( .I(n746), .Z(n745) );
  BUFFD0 U663 ( .I(n747), .Z(n746) );
  BUFFD0 U664 ( .I(n748), .Z(n747) );
  BUFFD0 U665 ( .I(n749), .Z(n748) );
  BUFFD0 U666 ( .I(n750), .Z(n749) );
  BUFFD0 U667 ( .I(n751), .Z(n750) );
  BUFFD0 U668 ( .I(n752), .Z(n751) );
  BUFFD0 U669 ( .I(ReadAddr[0]), .Z(n752) );
  BUFFD0 U670 ( .I(N48), .Z(n753) );
  BUFFD0 U671 ( .I(n756), .Z(n754) );
  BUFFD0 U672 ( .I(n753), .Z(n755) );
  BUFFD0 U673 ( .I(n758), .Z(n756) );
  BUFFD0 U674 ( .I(n755), .Z(n757) );
  BUFFD0 U675 ( .I(n760), .Z(n758) );
  BUFFD0 U676 ( .I(n757), .Z(n759) );
  BUFFD0 U677 ( .I(n762), .Z(n760) );
  BUFFD0 U678 ( .I(n759), .Z(n761) );
  BUFFD0 U679 ( .I(n764), .Z(n762) );
  BUFFD0 U680 ( .I(n761), .Z(n763) );
  BUFFD0 U681 ( .I(n766), .Z(n764) );
  BUFFD0 U682 ( .I(n763), .Z(n765) );
  BUFFD0 U683 ( .I(n768), .Z(n766) );
  BUFFD0 U684 ( .I(n765), .Z(n767) );
  BUFFD0 U685 ( .I(n770), .Z(n768) );
  BUFFD0 U686 ( .I(n767), .Z(n769) );
  BUFFD0 U687 ( .I(n772), .Z(n770) );
  BUFFD0 U688 ( .I(n769), .Z(n771) );
  BUFFD0 U689 ( .I(n774), .Z(n772) );
  BUFFD0 U690 ( .I(n771), .Z(n773) );
  BUFFD0 U691 ( .I(n776), .Z(n774) );
  BUFFD0 U692 ( .I(n773), .Z(n775) );
  BUFFD0 U693 ( .I(n778), .Z(n776) );
  BUFFD0 U694 ( .I(n775), .Z(n777) );
  BUFFD0 U695 ( .I(n780), .Z(n778) );
  BUFFD0 U696 ( .I(n777), .Z(n779) );
  BUFFD0 U697 ( .I(n782), .Z(n780) );
  BUFFD0 U698 ( .I(n779), .Z(n781) );
  BUFFD0 U699 ( .I(n784), .Z(n782) );
  BUFFD0 U700 ( .I(n781), .Z(n783) );
  BUFFD0 U701 ( .I(n785), .Z(n784) );
  BUFFD0 U702 ( .I(n786), .Z(n785) );
  BUFFD0 U703 ( .I(n787), .Z(n786) );
  BUFFD0 U704 ( .I(n789), .Z(n787) );
  BUFFD0 U705 ( .I(n35), .Z(n788) );
  BUFFD0 U706 ( .I(n791), .Z(n789) );
  BUFFD0 U707 ( .I(n788), .Z(n790) );
  BUFFD0 U708 ( .I(n793), .Z(n791) );
  BUFFD0 U709 ( .I(n790), .Z(n792) );
  BUFFD0 U710 ( .I(n795), .Z(n793) );
  BUFFD0 U711 ( .I(n792), .Z(n794) );
  BUFFD0 U712 ( .I(n796), .Z(n795) );
  BUFFD0 U713 ( .I(n906), .Z(n796) );
  CKBXD0 U714 ( .I(n783), .Z(n797) );
  BUFFD0 U715 ( .I(n802), .Z(n798) );
  BUFFD0 U716 ( .I(N63), .Z(n799) );
  BUFFD0 U717 ( .I(n799), .Z(n800) );
  BUFFD0 U718 ( .I(n800), .Z(n801) );
  BUFFD0 U719 ( .I(n803), .Z(n802) );
  BUFFD0 U720 ( .I(n804), .Z(n803) );
  BUFFD0 U721 ( .I(n805), .Z(n804) );
  BUFFD0 U722 ( .I(n806), .Z(n805) );
  BUFFD0 U723 ( .I(n807), .Z(n806) );
  BUFFD0 U724 ( .I(n808), .Z(n807) );
  BUFFD0 U725 ( .I(n809), .Z(n808) );
  BUFFD0 U726 ( .I(n810), .Z(n809) );
  BUFFD0 U727 ( .I(n811), .Z(n810) );
  BUFFD0 U728 ( .I(n812), .Z(n811) );
  BUFFD0 U729 ( .I(n813), .Z(n812) );
  BUFFD0 U730 ( .I(n814), .Z(n813) );
  BUFFD0 U731 ( .I(n815), .Z(n814) );
  BUFFD0 U732 ( .I(n816), .Z(n815) );
  BUFFD0 U733 ( .I(n817), .Z(n816) );
  BUFFD0 U734 ( .I(n818), .Z(n817) );
  BUFFD0 U735 ( .I(n819), .Z(n818) );
  BUFFD0 U736 ( .I(n820), .Z(n819) );
  BUFFD0 U737 ( .I(n821), .Z(n820) );
  BUFFD0 U738 ( .I(n822), .Z(n821) );
  BUFFD0 U739 ( .I(n823), .Z(n822) );
  BUFFD0 U740 ( .I(n824), .Z(n823) );
  BUFFD0 U741 ( .I(n825), .Z(n824) );
  BUFFD0 U742 ( .I(n826), .Z(n825) );
  BUFFD0 U743 ( .I(n827), .Z(n826) );
  BUFFD0 U744 ( .I(n828), .Z(n827) );
  BUFFD0 U745 ( .I(n829), .Z(n828) );
  BUFFD0 U746 ( .I(n830), .Z(n829) );
  BUFFD0 U747 ( .I(n831), .Z(n830) );
  BUFFD0 U748 ( .I(n832), .Z(n831) );
  BUFFD0 U749 ( .I(n833), .Z(n832) );
  BUFFD0 U750 ( .I(n834), .Z(n833) );
  BUFFD0 U751 ( .I(n835), .Z(n834) );
  BUFFD0 U752 ( .I(n836), .Z(n835) );
  BUFFD0 U753 ( .I(n837), .Z(n836) );
  BUFFD0 U754 ( .I(n838), .Z(n837) );
  BUFFD0 U755 ( .I(n839), .Z(n838) );
  BUFFD0 U756 ( .I(n840), .Z(n839) );
  BUFFD0 U757 ( .I(n841), .Z(n840) );
  BUFFD0 U758 ( .I(n842), .Z(n841) );
  BUFFD0 U759 ( .I(n843), .Z(n842) );
  BUFFD0 U760 ( .I(n844), .Z(n843) );
  BUFFD0 U761 ( .I(n845), .Z(n844) );
  BUFFD0 U762 ( .I(n846), .Z(n845) );
  BUFFD0 U763 ( .I(n847), .Z(n846) );
  BUFFD0 U764 ( .I(n848), .Z(n847) );
  BUFFD0 U765 ( .I(n849), .Z(n848) );
  BUFFD0 U766 ( .I(n850), .Z(n849) );
  BUFFD0 U767 ( .I(n851), .Z(n850) );
  BUFFD0 U768 ( .I(n852), .Z(n851) );
  BUFFD0 U769 ( .I(n853), .Z(n852) );
  BUFFD0 U770 ( .I(n854), .Z(n853) );
  BUFFD0 U771 ( .I(n855), .Z(n854) );
  BUFFD0 U772 ( .I(n856), .Z(n855) );
  BUFFD0 U773 ( .I(n801), .Z(n856) );
  BUFFD0 U774 ( .I(n907), .Z(n858) );
  CKBD0 U775 ( .CLK(N66), .C(n859) );
  CKBD0 U776 ( .CLK(n859), .C(n860) );
  CKBD0 U777 ( .CLK(n860), .C(n861) );
  CKBD0 U778 ( .CLK(n861), .C(n862) );
  CKBD0 U779 ( .CLK(n862), .C(n863) );
  CKBD0 U780 ( .CLK(n863), .C(n864) );
  CKBD0 U781 ( .CLK(n864), .C(n865) );
  CKBD0 U782 ( .CLK(n865), .C(n866) );
  CKBD0 U783 ( .CLK(n866), .C(n867) );
  CKBD0 U784 ( .CLK(n867), .C(n868) );
  CKBD0 U785 ( .CLK(n868), .C(n869) );
  CKBD0 U786 ( .CLK(n869), .C(n870) );
  CKBD0 U787 ( .CLK(n870), .C(n871) );
  CKBD0 U788 ( .CLK(n871), .C(n872) );
  CKBD0 U789 ( .CLK(n872), .C(n873) );
  CKBD0 U790 ( .CLK(n873), .C(n874) );
  CKBD0 U791 ( .CLK(n874), .C(n875) );
  CKBD0 U792 ( .CLK(n875), .C(n876) );
  CKBD0 U793 ( .CLK(n876), .C(n877) );
  CKBD0 U794 ( .CLK(n877), .C(n878) );
  CKBD0 U795 ( .CLK(n878), .C(n879) );
  CKBD0 U796 ( .CLK(n879), .C(n880) );
  CKBD0 U797 ( .CLK(n880), .C(n881) );
  CKBD0 U798 ( .CLK(n881), .C(n882) );
  CKBD0 U799 ( .CLK(n882), .C(n883) );
  CKBD0 U800 ( .CLK(n883), .C(n884) );
  CKBD0 U801 ( .CLK(n884), .C(n885) );
  CKBD0 U802 ( .CLK(n885), .C(n886) );
  CKBD0 U803 ( .CLK(n886), .C(n887) );
  CKBD0 U804 ( .CLK(n887), .C(n888) );
  CKBD0 U805 ( .CLK(n888), .C(n889) );
  CKBD0 U806 ( .CLK(n889), .C(n890) );
  CKBD0 U807 ( .CLK(n890), .C(n891) );
  CKBD0 U808 ( .CLK(n891), .C(n892) );
  CKBD0 U809 ( .CLK(n892), .C(n893) );
  BUFFD0 U810 ( .I(n37), .Z(n894) );
  BUFFD0 U811 ( .I(n893), .Z(n895) );
  BUFFD0 U812 ( .I(n895), .Z(n896) );
  BUFFD0 U813 ( .I(n896), .Z(n897) );
  BUFFD0 U814 ( .I(n897), .Z(n898) );
  BUFFD0 U815 ( .I(n898), .Z(n899) );
  BUFFD0 U816 ( .I(n899), .Z(n900) );
  BUFFD0 U817 ( .I(n900), .Z(n901) );
  BUFFD0 U818 ( .I(CurState[2]), .Z(n902) );
  INVD0 U819 ( .I(n40), .ZN(n35) );
  BUFFD0 U820 ( .I(CurState[1]), .Z(n903) );
  BUFFD0 U821 ( .I(n901), .Z(n904) );
  CKBD0 U822 ( .CLK(n903), .C(n905) );
  BUFFD0 U823 ( .I(n794), .Z(n906) );
  CKBD0 U824 ( .CLK(n904), .C(n907) );
  CKND2D0 U825 ( .A1(n905), .A2(n39), .ZN(n37) );
  OAI33XD4 U826 ( .A1(n915), .A2(n40), .A3(n86), .B1(n87), .B2(n88), .B3(n89), 
        .ZN(n136) );
  BUFFD0 U827 ( .I(n136), .Z(n908) );
  BUFFD0 U828 ( .I(n908), .Z(n909) );
  BUFFD0 U829 ( .I(n909), .Z(n910) );
  BUFFD0 U830 ( .I(n910), .Z(n911) );
  BUFFD0 U831 ( .I(n913), .Z(n912) );
  BUFFD0 U832 ( .I(n914), .Z(n913) );
  BUFFD0 U833 ( .I(n916), .Z(n914) );
  BUFFD0 U834 ( .I(n85), .Z(n915) );
  BUFFD0 U835 ( .I(n917), .Z(n916) );
  BUFFD0 U836 ( .I(n918), .Z(n917) );
  BUFFD0 U837 ( .I(n919), .Z(n918) );
  BUFFD0 U838 ( .I(n920), .Z(n919) );
  BUFFD0 U839 ( .I(n921), .Z(n920) );
  BUFFD0 U840 ( .I(n922), .Z(n921) );
  BUFFD0 U841 ( .I(n923), .Z(n922) );
  BUFFD0 U842 ( .I(n924), .Z(n923) );
  BUFFD0 U843 ( .I(n925), .Z(n924) );
  BUFFD0 U844 ( .I(n926), .Z(n925) );
  BUFFD0 U845 ( .I(n927), .Z(n926) );
  BUFFD0 U846 ( .I(n928), .Z(n927) );
  BUFFD0 U847 ( .I(n929), .Z(n928) );
  BUFFD0 U848 ( .I(n930), .Z(n929) );
  BUFFD0 U849 ( .I(n931), .Z(n930) );
  BUFFD0 U850 ( .I(n932), .Z(n931) );
  BUFFD0 U851 ( .I(n933), .Z(n932) );
  BUFFD0 U852 ( .I(n934), .Z(n933) );
  BUFFD0 U853 ( .I(n935), .Z(n934) );
  BUFFD0 U854 ( .I(n936), .Z(n935) );
  BUFFD0 U855 ( .I(n937), .Z(n936) );
  BUFFD0 U856 ( .I(n938), .Z(n937) );
  BUFFD0 U857 ( .I(n939), .Z(n938) );
  BUFFD0 U858 ( .I(n940), .Z(n939) );
  BUFFD0 U859 ( .I(n941), .Z(n940) );
  BUFFD0 U860 ( .I(n942), .Z(n941) );
  BUFFD0 U861 ( .I(n943), .Z(n942) );
  BUFFD0 U862 ( .I(n944), .Z(n943) );
  BUFFD0 U863 ( .I(n945), .Z(n944) );
  BUFFD0 U864 ( .I(n946), .Z(n945) );
  BUFFD0 U865 ( .I(n947), .Z(n946) );
  BUFFD0 U866 ( .I(n948), .Z(n947) );
  BUFFD0 U867 ( .I(n949), .Z(n948) );
  BUFFD0 U868 ( .I(n950), .Z(n949) );
  BUFFD0 U869 ( .I(n951), .Z(n950) );
  BUFFD0 U870 ( .I(n952), .Z(n951) );
  BUFFD0 U871 ( .I(n953), .Z(n952) );
  BUFFD0 U872 ( .I(n954), .Z(n953) );
  BUFFD0 U873 ( .I(n955), .Z(n954) );
  BUFFD0 U874 ( .I(n956), .Z(n955) );
  BUFFD0 U875 ( .I(n957), .Z(n956) );
  BUFFD0 U876 ( .I(n958), .Z(n957) );
  BUFFD0 U877 ( .I(n959), .Z(n958) );
  BUFFD0 U878 ( .I(n960), .Z(n959) );
  BUFFD0 U879 ( .I(n961), .Z(n960) );
  BUFFD0 U880 ( .I(n962), .Z(n961) );
  BUFFD0 U881 ( .I(n963), .Z(n962) );
  BUFFD0 U882 ( .I(n964), .Z(n963) );
  BUFFD0 U883 ( .I(n965), .Z(n964) );
  BUFFD0 U884 ( .I(n966), .Z(n965) );
  BUFFD0 U885 ( .I(n967), .Z(n966) );
  BUFFD0 U886 ( .I(n968), .Z(n967) );
  BUFFD0 U887 ( .I(n969), .Z(n968) );
  BUFFD0 U888 ( .I(n911), .Z(n969) );
  BUFFD0 U889 ( .I(n974), .Z(n970) );
  BUFFD0 U890 ( .I(n138), .Z(n971) );
  BUFFD0 U891 ( .I(n971), .Z(n972) );
  BUFFD0 U892 ( .I(n972), .Z(n973) );
  BUFFD0 U893 ( .I(n975), .Z(n974) );
  BUFFD0 U894 ( .I(n976), .Z(n975) );
  BUFFD0 U895 ( .I(n977), .Z(n976) );
  BUFFD0 U896 ( .I(n978), .Z(n977) );
  BUFFD0 U897 ( .I(n979), .Z(n978) );
  BUFFD0 U898 ( .I(n980), .Z(n979) );
  BUFFD0 U899 ( .I(n981), .Z(n980) );
  BUFFD0 U900 ( .I(n982), .Z(n981) );
  BUFFD0 U901 ( .I(n983), .Z(n982) );
  BUFFD0 U902 ( .I(n984), .Z(n983) );
  BUFFD0 U903 ( .I(n985), .Z(n984) );
  BUFFD0 U904 ( .I(n986), .Z(n985) );
  BUFFD0 U905 ( .I(n987), .Z(n986) );
  BUFFD0 U906 ( .I(n988), .Z(n987) );
  BUFFD0 U907 ( .I(n989), .Z(n988) );
  BUFFD0 U908 ( .I(n990), .Z(n989) );
  BUFFD0 U909 ( .I(n991), .Z(n990) );
  BUFFD0 U910 ( .I(n992), .Z(n991) );
  BUFFD0 U911 ( .I(n993), .Z(n992) );
  BUFFD0 U912 ( .I(n994), .Z(n993) );
  BUFFD0 U913 ( .I(n995), .Z(n994) );
  BUFFD0 U914 ( .I(n996), .Z(n995) );
  BUFFD0 U915 ( .I(n997), .Z(n996) );
  BUFFD0 U916 ( .I(n998), .Z(n997) );
  BUFFD0 U917 ( .I(n999), .Z(n998) );
  BUFFD0 U918 ( .I(n1000), .Z(n999) );
  BUFFD0 U919 ( .I(n1001), .Z(n1000) );
  BUFFD0 U920 ( .I(n1002), .Z(n1001) );
  BUFFD0 U921 ( .I(n1003), .Z(n1002) );
  BUFFD0 U922 ( .I(n1004), .Z(n1003) );
  BUFFD0 U923 ( .I(n1005), .Z(n1004) );
  BUFFD0 U924 ( .I(n1006), .Z(n1005) );
  BUFFD0 U925 ( .I(n1007), .Z(n1006) );
  BUFFD0 U926 ( .I(n1008), .Z(n1007) );
  BUFFD0 U927 ( .I(n1009), .Z(n1008) );
  BUFFD0 U928 ( .I(n1010), .Z(n1009) );
  BUFFD0 U929 ( .I(n1011), .Z(n1010) );
  BUFFD0 U930 ( .I(n1012), .Z(n1011) );
  BUFFD0 U931 ( .I(n1013), .Z(n1012) );
  BUFFD0 U932 ( .I(n1014), .Z(n1013) );
  BUFFD0 U933 ( .I(n1015), .Z(n1014) );
  BUFFD0 U934 ( .I(n1016), .Z(n1015) );
  BUFFD0 U935 ( .I(n1017), .Z(n1016) );
  BUFFD0 U936 ( .I(n1018), .Z(n1017) );
  BUFFD0 U937 ( .I(n1019), .Z(n1018) );
  BUFFD0 U938 ( .I(n1020), .Z(n1019) );
  BUFFD0 U939 ( .I(n1021), .Z(n1020) );
  BUFFD0 U940 ( .I(n1022), .Z(n1021) );
  BUFFD0 U941 ( .I(n1023), .Z(n1022) );
  BUFFD0 U942 ( .I(n1024), .Z(n1023) );
  BUFFD0 U943 ( .I(n1025), .Z(n1024) );
  BUFFD0 U944 ( .I(n1026), .Z(n1025) );
  BUFFD0 U945 ( .I(n1027), .Z(n1026) );
  BUFFD0 U946 ( .I(n1028), .Z(n1027) );
  BUFFD0 U947 ( .I(n973), .Z(n1028) );
  BUFFD0 U948 ( .I(n586), .Z(n1029) );
  CKBD0 U949 ( .CLK(n1029), .C(ReadCmd) );
  BUFFD0 U950 ( .I(n1032), .Z(n1031) );
  BUFFD0 U951 ( .I(n1033), .Z(n1032) );
  BUFFD0 U952 ( .I(n1034), .Z(n1033) );
  BUFFD0 U953 ( .I(n1035), .Z(n1034) );
  BUFFD0 U954 ( .I(n1036), .Z(n1035) );
  BUFFD0 U955 ( .I(n1037), .Z(n1036) );
  BUFFD0 U956 ( .I(n1039), .Z(n1037) );
  BUFFD0 U957 ( .I(OldWriteAr[1]), .Z(n1038) );
  BUFFD0 U958 ( .I(n1041), .Z(n1039) );
  CKBD0 U959 ( .CLK(n1038), .C(n1040) );
  BUFFD0 U960 ( .I(n1042), .Z(n1041) );
  BUFFD0 U961 ( .I(n1043), .Z(n1042) );
  BUFFD0 U962 ( .I(n1044), .Z(n1043) );
  BUFFD0 U963 ( .I(n1045), .Z(n1044) );
  BUFFD0 U964 ( .I(n1046), .Z(n1045) );
  BUFFD0 U965 ( .I(n1047), .Z(n1046) );
  BUFFD0 U966 ( .I(n1048), .Z(n1047) );
  BUFFD0 U967 ( .I(n1049), .Z(n1048) );
  BUFFD0 U968 ( .I(n1050), .Z(n1049) );
  BUFFD0 U969 ( .I(n1051), .Z(n1050) );
  BUFFD0 U970 ( .I(n1052), .Z(n1051) );
  BUFFD0 U971 ( .I(n1053), .Z(n1052) );
  BUFFD0 U972 ( .I(n1054), .Z(n1053) );
  BUFFD0 U973 ( .I(n1055), .Z(n1054) );
  BUFFD0 U974 ( .I(n1056), .Z(n1055) );
  BUFFD0 U975 ( .I(n1057), .Z(n1056) );
  BUFFD0 U976 ( .I(n1058), .Z(n1057) );
  BUFFD0 U977 ( .I(n1059), .Z(n1058) );
  BUFFD0 U978 ( .I(n1060), .Z(n1059) );
  BUFFD0 U979 ( .I(n1061), .Z(n1060) );
  BUFFD0 U980 ( .I(n1062), .Z(n1061) );
  BUFFD0 U981 ( .I(n1063), .Z(n1062) );
  BUFFD0 U982 ( .I(n1064), .Z(n1063) );
  BUFFD0 U983 ( .I(n1065), .Z(n1064) );
  BUFFD0 U984 ( .I(n1066), .Z(n1065) );
  BUFFD0 U985 ( .I(n1067), .Z(n1066) );
  BUFFD0 U986 ( .I(n1068), .Z(n1067) );
  BUFFD0 U987 ( .I(n1069), .Z(n1068) );
  BUFFD0 U988 ( .I(n1070), .Z(n1069) );
  BUFFD0 U989 ( .I(n1071), .Z(n1070) );
  BUFFD0 U990 ( .I(n1072), .Z(n1071) );
  BUFFD0 U991 ( .I(n1073), .Z(n1072) );
  BUFFD0 U992 ( .I(n1074), .Z(n1073) );
  BUFFD0 U993 ( .I(n1075), .Z(n1074) );
  BUFFD0 U994 ( .I(n1076), .Z(n1075) );
  BUFFD0 U995 ( .I(n1077), .Z(n1076) );
  BUFFD0 U996 ( .I(n1078), .Z(n1077) );
  BUFFD0 U997 ( .I(n1079), .Z(n1078) );
  BUFFD0 U998 ( .I(n1080), .Z(n1079) );
  BUFFD0 U999 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1000 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1001 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1002 ( .I(n1084), .Z(n1083) );
  BUFFD0 U1003 ( .I(n1085), .Z(n1084) );
  BUFFD0 U1004 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1005 ( .I(n1087), .Z(n1086) );
  BUFFD0 U1006 ( .I(n1088), .Z(n1087) );
  BUFFD0 U1007 ( .I(n1089), .Z(n1088) );
  BUFFD0 U1008 ( .I(n1090), .Z(n1089) );
  BUFFD0 U1009 ( .I(n1091), .Z(n1090) );
  BUFFD0 U1010 ( .I(n1092), .Z(n1091) );
  BUFFD0 U1011 ( .I(n131), .Z(n1092) );
  MOAI22D0 U1012 ( .A1(n42), .A2(n43), .B1(n42), .B2(n1040), .ZN(n131) );
  BUFFD0 U1013 ( .I(n1094), .Z(n1093) );
  BUFFD0 U1014 ( .I(n1095), .Z(n1094) );
  BUFFD0 U1015 ( .I(n1096), .Z(n1095) );
  BUFFD0 U1016 ( .I(n1097), .Z(n1096) );
  BUFFD0 U1017 ( .I(n1098), .Z(n1097) );
  BUFFD0 U1018 ( .I(n1099), .Z(n1098) );
  BUFFD0 U1019 ( .I(n1101), .Z(n1099) );
  BUFFD0 U1020 ( .I(OldWriteAr[2]), .Z(n1100) );
  BUFFD0 U1021 ( .I(n1103), .Z(n1101) );
  CKBD0 U1022 ( .CLK(n1100), .C(n1102) );
  BUFFD0 U1023 ( .I(n1104), .Z(n1103) );
  BUFFD0 U1024 ( .I(n1105), .Z(n1104) );
  BUFFD0 U1025 ( .I(n1106), .Z(n1105) );
  BUFFD0 U1026 ( .I(n1107), .Z(n1106) );
  BUFFD0 U1027 ( .I(n1108), .Z(n1107) );
  BUFFD0 U1028 ( .I(n1109), .Z(n1108) );
  BUFFD0 U1029 ( .I(n1110), .Z(n1109) );
  BUFFD0 U1030 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1031 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1032 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1033 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1034 ( .I(n1115), .Z(n1114) );
  BUFFD0 U1035 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1036 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1037 ( .I(n1118), .Z(n1117) );
  BUFFD0 U1038 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1039 ( .I(n1120), .Z(n1119) );
  BUFFD0 U1040 ( .I(n1121), .Z(n1120) );
  BUFFD0 U1041 ( .I(n1122), .Z(n1121) );
  BUFFD0 U1042 ( .I(n1123), .Z(n1122) );
  BUFFD0 U1043 ( .I(n1124), .Z(n1123) );
  BUFFD0 U1044 ( .I(n1125), .Z(n1124) );
  BUFFD0 U1045 ( .I(n1126), .Z(n1125) );
  BUFFD0 U1046 ( .I(n1127), .Z(n1126) );
  BUFFD0 U1047 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1048 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1049 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1050 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1051 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1052 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1053 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1054 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1055 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1056 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1057 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1058 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1059 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1060 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1061 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1062 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1063 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1064 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1065 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1066 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1067 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1068 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1069 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1070 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1071 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1072 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1073 ( .I(n1154), .Z(n1153) );
  MOAI22D0 U1074 ( .A1(n42), .A2(n44), .B1(n42), .B2(n1102), .ZN(n132) );
  BUFFD0 U1075 ( .I(n132), .Z(n1154) );
  BUFFD0 U1076 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1077 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1078 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1079 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1080 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1081 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1082 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1083 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1084 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1085 ( .I(n1165), .Z(n1164) );
  BUFFD0 U1086 ( .I(n1166), .Z(n1165) );
  BUFFD0 U1087 ( .I(n1167), .Z(n1166) );
  BUFFD0 U1088 ( .I(n1168), .Z(n1167) );
  BUFFD0 U1089 ( .I(n1169), .Z(n1168) );
  BUFFD0 U1090 ( .I(n1170), .Z(n1169) );
  BUFFD0 U1091 ( .I(n1171), .Z(n1170) );
  BUFFD0 U1092 ( .I(n1172), .Z(n1171) );
  BUFFD0 U1093 ( .I(n1173), .Z(n1172) );
  BUFFD0 U1094 ( .I(n1174), .Z(n1173) );
  BUFFD0 U1095 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1096 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1097 ( .I(n1177), .Z(n1176) );
  BUFFD0 U1098 ( .I(n1178), .Z(n1177) );
  BUFFD0 U1099 ( .I(n1179), .Z(n1178) );
  BUFFD0 U1100 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1101 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1102 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1103 ( .I(n1183), .Z(n1182) );
  BUFFD0 U1104 ( .I(n1184), .Z(n1183) );
  BUFFD0 U1105 ( .I(n1185), .Z(n1184) );
  BUFFD0 U1106 ( .I(n1186), .Z(n1185) );
  BUFFD0 U1107 ( .I(n1187), .Z(n1186) );
  BUFFD0 U1108 ( .I(n1188), .Z(n1187) );
  BUFFD0 U1109 ( .I(n1189), .Z(n1188) );
  BUFFD0 U1110 ( .I(n1190), .Z(n1189) );
  BUFFD0 U1111 ( .I(n1191), .Z(n1190) );
  BUFFD0 U1112 ( .I(n1192), .Z(n1191) );
  BUFFD0 U1113 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1114 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1115 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1116 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1117 ( .I(n1197), .Z(n1196) );
  BUFFD0 U1118 ( .I(n1198), .Z(n1197) );
  BUFFD0 U1119 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1120 ( .I(n1200), .Z(n1199) );
  BUFFD0 U1121 ( .I(n1201), .Z(n1200) );
  BUFFD0 U1122 ( .I(n1202), .Z(n1201) );
  BUFFD0 U1123 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1124 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1125 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1126 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1127 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1128 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1129 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1130 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1131 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1132 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1133 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1134 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1135 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1136 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1137 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1138 ( .I(n133), .Z(n1217) );
  BUFFD0 U1139 ( .I(n1222), .Z(n1218) );
  BUFFD0 U1140 ( .I(n130), .Z(n1219) );
  BUFFD0 U1141 ( .I(n1219), .Z(n1220) );
  BUFFD0 U1142 ( .I(n1220), .Z(n1221) );
  BUFFD0 U1143 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1144 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1145 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1146 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1147 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1148 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1149 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1150 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1151 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1152 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1153 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1154 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1155 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1156 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1157 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1158 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1159 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1160 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1161 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1162 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1163 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1164 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1165 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1166 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1167 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1168 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1169 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1170 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1171 ( .I(n1251), .Z(n1250) );
  BUFFD0 U1172 ( .I(n1252), .Z(n1251) );
  BUFFD0 U1173 ( .I(n1253), .Z(n1252) );
  BUFFD0 U1174 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1175 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1176 ( .I(n1256), .Z(n1255) );
  BUFFD0 U1177 ( .I(n1257), .Z(n1256) );
  BUFFD0 U1178 ( .I(n1258), .Z(n1257) );
  BUFFD0 U1179 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1180 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1181 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1182 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1183 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1184 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1185 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1186 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1187 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1188 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1189 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1190 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1191 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1192 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1193 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1194 ( .I(n1276), .Z(n1273) );
  BUFFD0 U1195 ( .I(OldReadAr[2]), .Z(n1274) );
  CKBD0 U1196 ( .CLK(n1274), .C(n1275) );
  BUFFD0 U1197 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1198 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1199 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1200 ( .I(n1221), .Z(n1279) );
  MOAI22D0 U1201 ( .A1(n141), .A2(n41), .B1(n41), .B2(n1275), .ZN(n130) );
  BUFFD0 U1202 ( .I(n1283), .Z(n1280) );
  BUFFD0 U1203 ( .I(n129), .Z(n1281) );
  BUFFD0 U1204 ( .I(n1281), .Z(n1282) );
  BUFFD0 U1205 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1206 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1207 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1208 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1209 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1210 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1211 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1212 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1213 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1214 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1215 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1216 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1217 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1218 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1219 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1220 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1221 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1222 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1223 ( .I(n1302), .Z(n1301) );
  BUFFD0 U1224 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1225 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1226 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1227 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1228 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1229 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1230 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1231 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1232 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1233 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1234 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1235 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1236 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1237 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1238 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1239 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1240 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1241 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1242 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1243 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1244 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1245 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1246 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1247 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1248 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1249 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1250 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1251 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1252 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1253 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1254 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1255 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1256 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1257 ( .I(n1337), .Z(n1335) );
  BUFFD0 U1258 ( .I(OldReadAr[1]), .Z(n1336) );
  BUFFD0 U1259 ( .I(n1339), .Z(n1337) );
  CKBD0 U1260 ( .CLK(n1336), .C(n1338) );
  BUFFD0 U1261 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1262 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1263 ( .I(n1282), .Z(n1341) );
  BUFFD0 U1264 ( .I(n1345), .Z(n1342) );
  BUFFD0 U1265 ( .I(n140), .Z(n1343) );
  BUFFD0 U1266 ( .I(n1343), .Z(n1344) );
  BUFFD0 U1267 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1268 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1269 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1270 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1271 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1272 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1273 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1274 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1275 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1276 ( .I(n1355), .Z(n1354) );
  BUFFD0 U1277 ( .I(n1356), .Z(n1355) );
  BUFFD0 U1278 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1279 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1280 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1281 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1282 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1283 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1284 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1285 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1286 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1287 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1288 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1289 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1290 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1291 ( .I(n1370), .Z(n1369) );
  BUFFD0 U1292 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1293 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1294 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1295 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1296 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1297 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1298 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1299 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1300 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1301 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1302 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1303 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1304 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1305 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1306 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1307 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1308 ( .I(n1387), .Z(n1386) );
  BUFFD0 U1309 ( .I(n1388), .Z(n1387) );
  BUFFD0 U1310 ( .I(n1389), .Z(n1388) );
  BUFFD0 U1311 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1312 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1313 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1314 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1315 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1316 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1317 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1318 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1319 ( .I(n1400), .Z(n1397) );
  BUFFD0 U1320 ( .I(OldReadAr[0]), .Z(n1398) );
  CKBD0 U1321 ( .CLK(n1398), .C(n1399) );
  BUFFD0 U1322 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1323 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1324 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1325 ( .I(n1344), .Z(n1403) );
  INVD1 U1326 ( .I(Reset), .ZN(n1410) );
  INVD1 U1327 ( .I(n77), .ZN(n84) );
  MAOI22D0 U1328 ( .A1(ReadAddr[0]), .A2(n75), .B1(n43), .B2(n98), .ZN(n101)
         );
  ND2D1 U1329 ( .A1(n83), .A2(n37), .ZN(n86) );
  ND2D1 U1330 ( .A1(WriteReq), .A2(n45), .ZN(n42) );
  ND2D1 U1331 ( .A1(ReadReq), .A2(n86), .ZN(n41) );
  INVD1 U1332 ( .I(n46), .ZN(n52) );
  NR2D1 U1333 ( .A1(n68), .A2(n79), .ZN(n39) );
  ND2D1 U1334 ( .A1(n83), .A2(n35), .ZN(n45) );
  XNR2D1 U1335 ( .A1(n44), .A2(n75), .ZN(n77) );
  INVD1 U1336 ( .I(n75), .ZN(n81) );
  XNR2D1 U1337 ( .A1(n84), .A2(ReadAddr[2]), .ZN(n56) );
  NR2D1 U1338 ( .A1(n700), .A2(n109), .ZN(N46) );
  NR2D1 U1339 ( .A1(n594), .A2(n109), .ZN(N49) );
  NR2D1 U1340 ( .A1(n650), .A2(n109), .ZN(N47) );
  INVD1 U1341 ( .I(ReadReq), .ZN(n106) );
  MAOI22D0 U1342 ( .A1(WriteAddr[0]), .A2(n103), .B1(n142), .B2(n98), .ZN(n102) );
  OAI222D0 U1343 ( .A1(n44), .A2(ReadAddr[2]), .B1(n43), .B2(ReadAddr[1]), 
        .C1(n144), .C2(ReadAddr[0]), .ZN(n73) );
  OAI33D1 U1344 ( .A1(ReadAddr[1]), .A2(WriteAddr[2]), .A3(n101), .B1(n44), 
        .B2(WriteAddr[1]), .B3(n102), .ZN(n54) );
  OAI33D1 U1345 ( .A1(ReadAddr[1]), .A2(n101), .A3(n44), .B1(n102), .B2(
        WriteAddr[2]), .B3(WriteAddr[1]), .ZN(n55) );
  AOI22D0 U1346 ( .A1(n68), .A2(CurState[1]), .B1(n51), .B2(n39), .ZN(n83) );
  NR3D0 U1347 ( .A1(n905), .A2(n902), .A3(CurState[0]), .ZN(n40) );
  AOI21D1 U1348 ( .A1(CurState[0]), .A2(n106), .B(n68), .ZN(n105) );
  INVD1 U1349 ( .I(WriteAddr[2]), .ZN(n44) );
  XNR2D1 U1350 ( .A1(n44), .A2(n1102), .ZN(n89) );
  XNR2D1 U1351 ( .A1(n43), .A2(n1040), .ZN(n88) );
  INVD1 U1352 ( .I(WriteAddr[1]), .ZN(n43) );
  NR2D1 U1353 ( .A1(n43), .A2(n144), .ZN(n75) );
  OAI211D1 U1354 ( .A1(n144), .A2(ReadAddr[1]), .B(n80), .C(n81), .ZN(n78) );
  OAI21D1 U1355 ( .A1(WriteAddr[1]), .A2(n142), .B(n143), .ZN(n80) );
  INVD1 U1356 ( .I(CurState[0]), .ZN(n79) );
  OAI32D1 U1357 ( .A1(n107), .A2(n108), .A3(n106), .B1(n86), .B2(n109), .ZN(
        n138) );
  XNR2D1 U1358 ( .A1(n142), .A2(n1338), .ZN(n108) );
  ND3D1 U1359 ( .A1(n110), .A2(n86), .A3(n111), .ZN(n107) );
  XNR2D1 U1360 ( .A1(ReadAddr[2]), .A2(n1275), .ZN(n110) );
  XOR2D1 U1361 ( .A1(n100), .A2(n142), .Z(n57) );
  INVD1 U1362 ( .I(n902), .ZN(n68) );
  ND2D1 U1363 ( .A1(n144), .A2(n143), .ZN(n98) );
  AOI31D0 U1364 ( .A1(n65), .A2(n66), .A3(n67), .B(n68), .ZN(n64) );
  AOI22D0 U1365 ( .A1(n69), .A2(ReadAddr[1]), .B1(n144), .B2(ReadAddr[0]), 
        .ZN(n67) );
  OAI21D1 U1366 ( .A1(n69), .A2(n73), .B(n43), .ZN(n65) );
  OAI21D1 U1367 ( .A1(ReadAddr[1]), .A2(n72), .B(n73), .ZN(n66) );
  OAI22D0 U1368 ( .A1(n46), .A2(n352), .B1(n52), .B2(n59), .ZN(n135) );
  AOI31D0 U1369 ( .A1(n60), .A2(n61), .A3(n62), .B(n40), .ZN(n59) );
  IIND4D1 U1370 ( .A1(n69), .A2(n73), .B1(n78), .B2(n79), .ZN(n61) );
  AOI31D0 U1371 ( .A1(n143), .A2(CurState[0]), .A3(n63), .B(n64), .ZN(n62) );
  OAI22D0 U1372 ( .A1(n46), .A2(n291), .B1(n52), .B2(n92), .ZN(n137) );
  AOI21D1 U1373 ( .A1(CurState[1]), .A2(n93), .B(n39), .ZN(n92) );
  OAI21D1 U1374 ( .A1(CurState[2]), .A2(n94), .B(n95), .ZN(n93) );
  AOI22D0 U1375 ( .A1(n55), .A2(ReadAddr[2]), .B1(n141), .B2(n54), .ZN(n94) );
  OAI31D0 U1376 ( .A1(n96), .A2(n97), .A3(n58), .B(CurState[0]), .ZN(n95) );
  XNR2D1 U1377 ( .A1(WriteAddr[2]), .A2(n99), .ZN(n97) );
  INVD1 U1378 ( .I(n57), .ZN(n96) );
  OAI211D1 U1379 ( .A1(CurState[2]), .A2(n48), .B(CurState[0]), .C(n49), .ZN(
        n47) );
  AOI21D1 U1380 ( .A1(n50), .A2(n51), .B(n52), .ZN(n49) );
  NR4D0 U1381 ( .A1(n56), .A2(n57), .A3(n51), .A4(n58), .ZN(n48) );
  INVD1 U1382 ( .I(CurState[1]), .ZN(n51) );
  NR3D0 U1383 ( .A1(n57), .A2(n144), .A3(n74), .ZN(n63) );
  AOI21D1 U1384 ( .A1(n69), .A2(n75), .B(n76), .ZN(n74) );
  OAI32D1 U1385 ( .A1(n44), .A2(n141), .A3(n75), .B1(ReadAddr[2]), .B2(n77), 
        .ZN(n76) );
  AOI31D0 U1386 ( .A1(n144), .A2(CurState[0]), .A3(n82), .B(n83), .ZN(n60) );
  NR3D0 U1387 ( .A1(n57), .A2(n143), .A3(n56), .ZN(n82) );
  NR2D1 U1388 ( .A1(n143), .A2(n641), .ZN(n103) );
  XOR2D1 U1389 ( .A1(n103), .A2(n642), .Z(n99) );
  AO22D0 U1390 ( .A1(ReadAddr[2]), .A2(n54), .B1(n55), .B2(n141), .Z(n50) );
  XNR2D1 U1391 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n72) );
  ND2D1 U1392 ( .A1(ReadCmd), .A2(n2), .ZN(n109) );
  OAI21D1 U1393 ( .A1(n144), .A2(n143), .B(n98), .ZN(n58) );
  OAI32D1 U1394 ( .A1(n37), .A2(Reset), .A3(ReadReq), .B1(n38), .B2(n166), 
        .ZN(n128) );
  ND2D1 U1395 ( .A1(n1412), .A2(n894), .ZN(n112) );
  NR2D1 U1396 ( .A1(WriteAddr[2]), .A2(n141), .ZN(n69) );
  OAI22D0 U1397 ( .A1(n143), .A2(n894), .B1(n857), .B2(n112), .ZN(N63) );
  OAI22D0 U1398 ( .A1(n642), .A2(n894), .B1(n84), .B2(n112), .ZN(N65) );
  OAI22D0 U1399 ( .A1(n641), .A2(n894), .B1(n100), .B2(n112), .ZN(N64) );
  OAI31D0 U1400 ( .A1(n35), .A2(WriteReq), .A3(Reset), .B(n10), .ZN(n127) );
  OAI31D0 U1401 ( .A1(CurState[0]), .A2(Reset), .A3(CurState[2]), .B(EmptyFIFO), .ZN(n36) );
  ND3D1 U1402 ( .A1(n90), .A2(n45), .A3(WriteReq), .ZN(n87) );
  XNR2D1 U1403 ( .A1(WriteAddr[0]), .A2(OldWriteAr[0]), .ZN(n90) );
  XNR2D1 U1404 ( .A1(ReadAddr[0]), .A2(n1399), .ZN(n111) );
  ND2D1 U1405 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
endmodule


module DPMem1kx32_AWid3_DWid32_0 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [2:0] AddrR;
  input [2:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N48, N49, N50, ClockW, Dreadyr, \Storage[7][32] , \Storage[7][31] ,
         \Storage[7][30] , \Storage[7][29] , \Storage[7][28] ,
         \Storage[7][27] , \Storage[7][26] , \Storage[7][25] ,
         \Storage[7][24] , \Storage[7][23] , \Storage[7][22] ,
         \Storage[7][21] , \Storage[7][20] , \Storage[7][19] ,
         \Storage[7][18] , \Storage[7][17] , \Storage[7][16] ,
         \Storage[7][15] , \Storage[7][14] , \Storage[7][13] ,
         \Storage[7][12] , \Storage[7][11] , \Storage[7][10] , \Storage[7][9] ,
         \Storage[7][8] , \Storage[7][7] , \Storage[7][6] , \Storage[7][5] ,
         \Storage[7][4] , \Storage[7][3] , \Storage[7][2] , \Storage[7][1] ,
         \Storage[7][0] , \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N87, N194, N293, N326, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854;
  wire   [31:0] DataOr;
  assign N48 = AddrR[0];
  assign N49 = AddrR[1];
  assign N50 = AddrR[2];

  XNR4D1 U13 ( .A1(n1223), .A2(n3744), .A3(n3747), .A4(n1208), .ZN(n78) );
  XOR4D1 U14 ( .A1(n1174), .A2(n3748), .A3(n3751), .A4(n1159), .Z(n77) );
  XOR4D1 U15 ( .A1(n3742), .A2(n3741), .A3(DataI[23]), .A4(n3743), .Z(n74) );
  XOR4D1 U16 ( .A1(n3736), .A2(DataI[13]), .A3(DataI[16]), .A4(n3737), .Z(n71)
         );
  XOR4D1 U21 ( .A1(n83), .A2(N74), .A3(n84), .A4(N77), .Z(n82) );
  XNR4D1 U22 ( .A1(N71), .A2(N70), .A3(N73), .A4(N72), .ZN(n84) );
  XNR4D1 U27 ( .A1(N53), .A2(N52), .A3(N55), .A4(N54), .ZN(n90) );
  XOR4D1 U28 ( .A1(N57), .A2(N56), .A3(N59), .A4(N58), .Z(n89) );
  XNR4D1 U29 ( .A1(N64), .A2(N63), .A3(N66), .A4(N65), .ZN(n86) );
  XNR4D1 U30 ( .A1(N82), .A2(N80), .A3(N84), .A4(N83), .ZN(n80) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n12), .E(n3766), .CP(n3811), .CDN(n3828), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n147), .E(n3766), .CP(n3778), .CDN(n3828), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n203), .E(n3766), .CP(n3778), .CDN(n3827), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n205), .E(n3766), .CP(n3777), .CDN(n3827), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n312), .E(n3766), .CP(n3807), .CDN(n3827), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n368), .E(n3766), .CP(n3808), .CDN(n3827), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n370), .E(n3766), .CP(n3806), .CDN(n3827), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n423), .E(n3766), .CP(n3805), .CDN(n3827), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n530), .E(n3766), .CP(n3804), .CDN(n3827), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n586), .E(n3764), .CP(n3809), .CDN(n3827), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n589), .E(n3766), .CP(n3774), .CDN(n3826), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n696), .E(N194), .CP(n3803), .CDN(n3826), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n752), .E(N194), .CP(ClockW), .CDN(n3826), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n754), .E(N194), .CP(n3802), .CDN(n3826), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n807), .E(N194), .CP(ClockW), .CDN(n3826), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n915), .E(N194), .CP(n3776), .CDN(n3826), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n971), .E(N194), .CP(n3775), .CDN(n3826), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n973), .E(n3764), .CP(n3809), .CDN(n3826), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n975), .E(N194), .CP(n3773), .CDN(n3826), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n1024), .E(n3764), .CP(n3774), .CDN(n3826), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n12), .E(n3770), .CP(n3798), .CDN(n3822), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n147), .E(n3771), .CP(n3798), .CDN(n3822), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n203), .E(n3771), .CP(n3799), .CDN(n3821), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n205), .E(n3771), .CP(n3799), .CDN(n3821), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n312), .E(n3771), .CP(n3799), .CDN(n3821), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n368), .E(n3771), .CP(n3799), .CDN(n3821), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n370), .E(n3771), .CP(n3799), .CDN(n3821), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n423), .E(n3769), .CP(n3799), .CDN(n3821), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n530), .E(n3771), .CP(n3800), .CDN(n3821), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n586), .E(n3770), .CP(n3800), .CDN(n3821), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n589), .E(n3769), .CP(n3800), .CDN(n3820), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n696), .E(n3769), .CP(n3800), .CDN(n3820), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n752), .E(n3769), .CP(n3800), .CDN(n3820), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n754), .E(n3769), .CP(n3800), .CDN(n3820), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n807), .E(n3769), .CP(n3800), .CDN(n3820), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n915), .E(n3769), .CP(n3800), .CDN(n3820), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n971), .E(n3769), .CP(n3800), .CDN(n3820), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n3728), .E(n3769), .CP(n3801), .CDN(n3820), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n9), .E(n3769), .CP(n3801), .CDN(n3820), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n3726), .E(n3769), .CP(n3801), .CDN(n3820), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n12), .E(n3754), .CP(n3783), .CDN(n3840), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n147), .E(n3755), .CP(n3783), .CDN(n3840), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n203), .E(n3755), .CP(n3784), .CDN(n3839), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n205), .E(n3755), .CP(n3784), .CDN(n3839), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n312), .E(n3755), .CP(n3784), .CDN(n3839), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n368), .E(n3755), .CP(n3784), .CDN(n3839), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n370), .E(n3755), .CP(n3784), .CDN(n3839), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n423), .E(N326), .CP(n3784), .CDN(n3839), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n530), .E(n3754), .CP(n3785), .CDN(n3839), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n586), .E(n3755), .CP(n3785), .CDN(n3839), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n589), .E(n3754), .CP(n3785), .CDN(n3838), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n696), .E(n3755), .CP(n3785), .CDN(n3838), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n752), .E(N326), .CP(n3785), .CDN(n3838), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n754), .E(N326), .CP(n3785), .CDN(n3838), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n807), .E(N326), .CP(n3785), .CDN(n3838), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n915), .E(N326), .CP(n3785), .CDN(n3838), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n971), .E(N326), .CP(n3785), .CDN(n3838), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n973), .E(n3755), .CP(n3786), .CDN(n3838), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n975), .E(n3755), .CP(n3786), .CDN(n3838), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n1024), .E(n3755), .CP(n3786), .CDN(n3838), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n12), .E(n3757), .CP(n3787), .CDN(n3837), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n147), .E(n3758), .CP(n3787), .CDN(n3837), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n203), .E(n3758), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n205), .E(n3758), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n312), .E(n3758), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n368), .E(n3758), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n370), .E(n3758), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n423), .E(N293), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n530), .E(n3757), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n586), .E(n3758), .CP(n3788), .CDN(n3836), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n589), .E(n3757), .CP(n3788), .CDN(n3835), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n696), .E(n3758), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n752), .E(N293), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n754), .E(N293), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n807), .E(N293), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n915), .E(N293), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n971), .E(N293), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n973), .E(n3758), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n975), .E(n3758), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n1024), .E(n3758), .CP(n3789), .CDN(n3835), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n12), .E(n3760), .CP(n3791), .CDN(n3834), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n147), .E(n3760), .CP(n3791), .CDN(n3834), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n203), .E(n3760), .CP(n3791), .CDN(n3833), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n205), .E(n3760), .CP(n3791), .CDN(n3833), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n312), .E(n3760), .CP(n3791), .CDN(n3833), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n368), .E(n3760), .CP(n3792), .CDN(n3833), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n370), .E(n3760), .CP(n3792), .CDN(n3833), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n423), .E(n3761), .CP(n3792), .CDN(n3833), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n530), .E(n3761), .CP(n3792), .CDN(n3833), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n586), .E(n3761), .CP(n3792), .CDN(n3833), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n589), .E(n3761), .CP(n3792), .CDN(n3832), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n696), .E(n3761), .CP(n3792), .CDN(n3832), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n752), .E(n3761), .CP(n3792), .CDN(n3832), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n754), .E(n3761), .CP(n3792), .CDN(n3832), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n807), .E(n3761), .CP(n3793), .CDN(n3832), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n915), .E(n3761), .CP(n3793), .CDN(n3832), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n971), .E(n3761), .CP(n3793), .CDN(n3832), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n973), .E(n3761), .CP(n3793), .CDN(n3832), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n975), .E(n3760), .CP(n3793), .CDN(n3832), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n1024), .E(n3761), .CP(n3793), .CDN(n3832), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n12), .E(n3763), .CP(n3794), .CDN(n3831), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n147), .E(n3762), .CP(n3794), .CDN(n3831), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n203), .E(n3762), .CP(n3795), .CDN(n3830), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n205), .E(n3763), .CP(n3795), .CDN(n3830), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n312), .E(n3762), .CP(n3795), .CDN(n3830), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n368), .E(n3763), .CP(n3795), .CDN(n3830), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n370), .E(n3762), .CP(n3795), .CDN(n3830), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n423), .E(n3762), .CP(n3795), .CDN(n3830), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n530), .E(n3762), .CP(n3796), .CDN(n3830), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n586), .E(n3762), .CP(n3796), .CDN(n3830), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n589), .E(n3762), .CP(n3796), .CDN(n3829), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n696), .E(n3762), .CP(n3796), .CDN(n3829), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n752), .E(n3762), .CP(n3796), .CDN(n3829), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n754), .E(n3762), .CP(n3796), .CDN(n3829), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n807), .E(n3762), .CP(n3796), .CDN(n3829), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n915), .E(n3762), .CP(n3796), .CDN(n3829), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n971), .E(n3762), .CP(n3796), .CDN(n3829), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n973), .E(n3763), .CP(n3797), .CDN(n3829), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n975), .E(n3763), .CP(n3797), .CDN(n3829), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n1024), .E(n3763), .CP(n3797), .CDN(n3829), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n12), .E(n3767), .CP(n3773), .CDN(n3825), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n147), .E(n3768), .CP(n3807), .CDN(n3825), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n203), .E(n3768), .CP(n3806), .CDN(n3824), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n205), .E(n3768), .CP(n3805), .CDN(n3824), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n312), .E(n3768), .CP(n3777), .CDN(n3824), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n368), .E(n3768), .CP(n3778), .CDN(n3824), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n370), .E(n3768), .CP(n3808), .CDN(n3824), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n423), .E(n3768), .CP(n3810), .CDN(n3824), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n530), .E(n3767), .CP(n3811), .CDN(n3824), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n586), .E(n3767), .CP(n3812), .CDN(n3824), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n589), .E(n3768), .CP(n3804), .CDN(n3823), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n696), .E(n3767), .CP(n3805), .CDN(n3823), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n752), .E(n3768), .CP(n3806), .CDN(n3823), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n754), .E(n3767), .CP(n3810), .CDN(n3823), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n807), .E(n3768), .CP(n3777), .CDN(n3823), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n915), .E(n3767), .CP(n3808), .CDN(n3823), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n971), .E(n3768), .CP(n3801), .CDN(n3823), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n973), .E(n3768), .CP(n3773), .CDN(n3823), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n975), .E(n3768), .CP(n3809), .CDN(n3823), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n1024), .E(n3768), .CP(n3774), .CDN(n3823), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n12), .E(n3752), .CP(n3780), .CDN(n3843), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n147), .E(n3752), .CP(n3780), .CDN(n3843), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n203), .E(n3752), .CP(n3780), .CDN(n3842), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n205), .E(n3752), .CP(n3780), .CDN(n3842), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n312), .E(n3752), .CP(n3780), .CDN(n3842), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n368), .E(n3752), .CP(n3781), .CDN(n3842), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n370), .E(n3752), .CP(n3781), .CDN(n3842), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n423), .E(n3752), .CP(n3781), .CDN(n3842), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n530), .E(n3752), .CP(n3781), .CDN(n3842), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n586), .E(n3752), .CP(n3781), .CDN(n3842), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n589), .E(n3752), .CP(n3781), .CDN(n3841), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n696), .E(n3752), .CP(n3781), .CDN(n3841), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n752), .E(n3753), .CP(n3781), .CDN(n3841), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n754), .E(n3752), .CP(n3781), .CDN(n3841), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n807), .E(n3753), .CP(n3782), .CDN(n3841), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n915), .E(n3752), .CP(n3782), .CDN(n3841), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n971), .E(n3753), .CP(n3782), .CDN(n3841), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n973), .E(n3753), .CP(n3782), .CDN(n3841), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n975), .E(n3753), .CP(n3782), .CDN(n3841), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n1024), .E(n3753), .CP(n3782), .CDN(n3841), 
        .Q(\Storage[7][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n1025), .CP(n3813), .CDN(n3820), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(n1137), .E(n3764), .CP(n3797), .CDN(n3829), .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n1138), .E(n3764), .CP(n3797), .CDN(n3828), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n1162), .E(n3764), .CP(n3797), .CDN(n3828), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n1177), .E(n3766), .CP(n3797), .CDN(n3828), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n1178), .E(n3766), .CP(n3797), .CDN(n3828), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n1188), .E(n3764), .CP(n3797), .CDN(n3828), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n1212), .E(n3766), .CP(n3810), .CDN(n3828), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n1227), .E(n3766), .CP(n3802), .CDN(n3828), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n1229), .E(n3764), .CP(n3807), .CDN(n3828), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n1243), .E(n3766), .CP(n3803), .CDN(n3828), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n1245), .E(n3766), .CP(n3802), .CDN(n3827), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n1252), .E(n3766), .CP(n3777), .CDN(n3827), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n1266), .E(n3766), .CP(n3812), .CDN(n3827), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(n1137), .E(n3770), .CP(n3775), .CDN(n3823), .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n1138), .E(n3770), .CP(n3776), .CDN(n3822), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n1162), .E(n3770), .CP(ClockW), .CDN(
        n3822), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n1177), .E(n3770), .CP(n3798), .CDN(n3822), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n1178), .E(n3770), .CP(n3798), .CDN(n3822), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n1188), .E(n3770), .CP(n3798), .CDN(n3822), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n1212), .E(n3770), .CP(n3798), .CDN(n3822), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n1227), .E(n3770), .CP(n3798), .CDN(n3822), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n1229), .E(n3770), .CP(n3798), .CDN(n3822), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n1243), .E(n3771), .CP(n3798), .CDN(n3822), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n1245), .E(n3771), .CP(n3799), .CDN(n3821), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n1252), .E(n3771), .CP(n3799), .CDN(n3821), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n1266), .E(n3771), .CP(n3799), .CDN(n3821), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(n1137), .E(n3754), .CP(n3782), .CDN(n3841), .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n1138), .E(n3754), .CP(n3782), .CDN(n3840), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n1162), .E(n3754), .CP(n3782), .CDN(n3840), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n1177), .E(n3754), .CP(n3783), .CDN(n3840), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n1178), .E(n3754), .CP(n3783), .CDN(n3840), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n1188), .E(n3754), .CP(n3783), .CDN(n3840), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n1212), .E(n3754), .CP(n3783), .CDN(n3840), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n1227), .E(n3754), .CP(n3783), .CDN(n3840), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n1229), .E(n3754), .CP(n3783), .CDN(n3840), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n1243), .E(n3755), .CP(n3783), .CDN(n3840), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n1245), .E(n3755), .CP(n3784), .CDN(n3839), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n1252), .E(N326), .CP(n3784), .CDN(n3839), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n1266), .E(n3754), .CP(n3784), .CDN(n3839), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(n1137), .E(n3757), .CP(n3786), .CDN(n3838), .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n1138), .E(n3757), .CP(n3786), .CDN(n3837), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n1162), .E(n3757), .CP(n3786), .CDN(n3837), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n1177), .E(n3757), .CP(n3786), .CDN(n3837), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n1178), .E(n3757), .CP(n3786), .CDN(n3837), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n1188), .E(n3757), .CP(n3786), .CDN(n3837), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n1212), .E(n3757), .CP(n3787), .CDN(n3837), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n1227), .E(n3757), .CP(n3787), .CDN(n3837), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n1229), .E(n3757), .CP(n3787), .CDN(n3837), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n1243), .E(n3758), .CP(n3787), .CDN(n3837), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n1245), .E(n3758), .CP(n3787), .CDN(n3836), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n1252), .E(N293), .CP(n3787), .CDN(n3836), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n1266), .E(n3757), .CP(n3787), .CDN(n3836), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(n1137), .E(n3760), .CP(n3790), .CDN(n3835), .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n1138), .E(n3761), .CP(n3790), .CDN(n3834), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n1162), .E(n3760), .CP(n3790), .CDN(n3834), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n1177), .E(n3761), .CP(n3790), .CDN(n3834), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n1178), .E(n3760), .CP(n3790), .CDN(n3834), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n1188), .E(n3761), .CP(n3790), .CDN(n3834), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n1212), .E(n3760), .CP(n3790), .CDN(n3834), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n1227), .E(n3761), .CP(n3790), .CDN(n3834), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n1229), .E(n3760), .CP(n3790), .CDN(n3834), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n1243), .E(n3760), .CP(n3791), .CDN(n3834), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n1245), .E(n3760), .CP(n3791), .CDN(n3833), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n1252), .E(n3760), .CP(n3791), .CDN(n3833), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n1266), .E(n3760), .CP(n3791), .CDN(n3833), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(n1137), .E(n3763), .CP(n3793), .CDN(n3832), .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n1138), .E(n3763), .CP(n3793), .CDN(n3831), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n1162), .E(n3763), .CP(n3793), .CDN(n3831), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n1177), .E(n3763), .CP(n3794), .CDN(n3831), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n1178), .E(n3763), .CP(n3794), .CDN(n3831), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n1188), .E(n3763), .CP(n3794), .CDN(n3831), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n1212), .E(n3763), .CP(n3794), .CDN(n3831), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n1227), .E(n3762), .CP(n3794), .CDN(n3831), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n1229), .E(n3763), .CP(n3794), .CDN(n3831), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n1243), .E(n3763), .CP(n3794), .CDN(n3831), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n1245), .E(n3762), .CP(n3795), .CDN(n3830), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n1252), .E(n3763), .CP(n3795), .CDN(n3830), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n1266), .E(n3762), .CP(n3795), .CDN(n3830), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(n1137), .E(n3767), .CP(n3804), .CDN(n3826), .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n1138), .E(n3767), .CP(n3775), .CDN(n3825), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n1162), .E(n3767), .CP(n3803), .CDN(n3825), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n1177), .E(n3767), .CP(n3811), .CDN(n3825), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n1178), .E(n3767), .CP(n3808), .CDN(n3825), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n1188), .E(n3767), .CP(n3807), .CDN(n3825), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n1212), .E(n3767), .CP(n3810), .CDN(n3825), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n1227), .E(n3767), .CP(n3812), .CDN(n3825), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n1229), .E(n3767), .CP(n3811), .CDN(n3825), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n1243), .E(n3768), .CP(n3778), .CDN(n3825), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n1245), .E(n3768), .CP(n3776), .CDN(n3824), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n1252), .E(n3767), .CP(n3801), .CDN(n3824), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n1266), .E(n3768), .CP(ClockW), .CDN(
        n3824), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(n1137), .E(n3753), .CP(n3779), .CDN(n3844), .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n1138), .E(n3753), .CP(n3779), .CDN(n3843), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n1162), .E(n3753), .CP(n3779), .CDN(n3843), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n1177), .E(n3753), .CP(n3779), .CDN(n3843), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n1178), .E(n3753), .CP(n3779), .CDN(n3843), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n1188), .E(n3752), .CP(n3779), .CDN(n3843), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n1212), .E(n3753), .CP(n3779), .CDN(n3843), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n1227), .E(n3752), .CP(n3779), .CDN(n3843), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n1229), .E(n3753), .CP(n3779), .CDN(n3843), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n1243), .E(n3752), .CP(n3780), .CDN(n3843), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n1245), .E(n3752), .CP(n3780), .CDN(n3842), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n1252), .E(n3752), .CP(n3780), .CDN(n3842), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n1266), .E(n3753), .CP(n3780), .CDN(n3842), .Q(\Storage[7][18] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n1268), .E(n3816), .CP(n3813), .CDN(n3852), 
        .Q(DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n1338), .E(n3816), .CP(n3813), .CDN(n3825), 
        .Q(DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n1408), .E(n3816), .CP(n3814), .CDN(n3849), 
        .Q(DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n1478), .E(n3816), .CP(n3813), .CDN(n3853), 
        .Q(DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n1548), .E(n3816), .CP(n3814), .CDN(n3849), 
        .Q(DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n1618), .E(n3816), .CP(n3814), .CDN(n3846), 
        .Q(DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n1688), .E(n3816), .CP(n3814), .CDN(n3831), 
        .Q(DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n1758), .E(n3816), .CP(n3813), .CDN(n3841), 
        .Q(DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n1828), .E(n3816), .CP(n3814), .CDN(n3823), 
        .Q(DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n1898), .E(n3816), .CP(n3813), .CDN(n3840), 
        .Q(DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n1968), .E(n3816), .CP(n3813), .CDN(n3822), 
        .Q(DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n2038), .E(n3816), .CP(n3813), .CDN(n3821), 
        .Q(DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n2108), .E(n3816), .CP(n3813), .CDN(n3824), 
        .Q(DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n2178), .E(n3816), .CP(n3813), .CDN(n3835), 
        .Q(DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n2248), .E(n3816), .CP(n3813), .CDN(n3831), 
        .Q(DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n2318), .E(n3816), .CP(n3813), .CDN(n3853), 
        .Q(DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n2388), .E(n3816), .CP(n3813), .CDN(n3824), 
        .Q(DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n2458), .E(n3815), .CP(n3813), .CDN(n3831), 
        .Q(DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n2528), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n2598), .E(n3815), .CP(n3814), .CDN(n3821), 
        .Q(DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n2668), .E(n3815), .CP(n3814), .CDN(n3835), 
        .Q(DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n2738), .E(n3815), .CP(n3814), .CDN(n3831), 
        .Q(DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n2808), .E(n3815), .CP(n3814), .CDN(n3820), 
        .Q(DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n2878), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n2947), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n3017), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n3087), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n3157), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n1), .E(n3815), .CP(n3813), .CDN(n3844), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n3294), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n3363), .E(n3815), .CP(n3814), .CDN(n3844), 
        .Q(DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n3432), .E(n3815), .CP(n3813), .CDN(n3844), 
        .Q(DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(n3503), .E(n3815), .CP(n3813), .CDN(n3844), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  BUFFD0 U3 ( .I(n3226), .Z(n1) );
  BUFFD0 U4 ( .I(n3569), .Z(n2) );
  CKBD0 U5 ( .CLK(DataI[0]), .C(n3726) );
  INVD0 U6 ( .I(n1023), .ZN(n1024) );
  CKBD0 U7 ( .CLK(DataI[2]), .C(n3728) );
  INVD0 U8 ( .I(n972), .ZN(n973) );
  CKBD0 U9 ( .CLK(n1246), .C(n1245) );
  CKBD0 U10 ( .CLK(n1230), .C(n1229) );
  CKBD0 U11 ( .CLK(n1253), .C(n1252) );
  CKBD0 U12 ( .CLK(n1139), .C(n1138) );
  CKBD0 U17 ( .CLK(n1189), .C(n1188) );
  CKBD0 U18 ( .CLK(n1179), .C(n1178) );
  CKBD0 U19 ( .CLK(n590), .C(n589) );
  CKBD0 U20 ( .CLK(n371), .C(n370) );
  CKBD0 U23 ( .CLK(n13), .C(n12) );
  CKBD0 U24 ( .CLK(n808), .C(n807) );
  CKBD0 U25 ( .CLK(n755), .C(n754) );
  CKBD0 U26 ( .CLK(n206), .C(n205) );
  CKBD0 U31 ( .CLK(n424), .C(n423) );
  OR3D1 U32 ( .A1(n1267), .A2(AddrW[1]), .A3(AddrW[0]), .Z(n3) );
  OR3D1 U33 ( .A1(n93), .A2(AddrW[1]), .A3(n10), .Z(n4) );
  CKND2D0 U34 ( .A1(ClkR), .A2(ChipEna), .ZN(n5) );
  OR3D1 U35 ( .A1(n91), .A2(n10), .A3(n93), .Z(n6) );
  INVD0 U36 ( .I(n8), .ZN(n3769) );
  OR3D1 U37 ( .A1(n91), .A2(n1267), .A3(n93), .Z(n7) );
  INVD0 U38 ( .I(n3765), .ZN(n3764) );
  OR3D1 U39 ( .A1(n66), .A2(AddrW[1]), .A3(AddrW[0]), .Z(n8) );
  XNR4D0 U40 ( .A1(n3732), .A2(n3731), .A3(DataI[9]), .A4(n3733), .ZN(n68) );
  BUFFD0 U41 ( .I(n974), .Z(n9) );
  BUFFD0 U42 ( .I(n66), .Z(n10) );
  CKBD0 U43 ( .CLK(DataI[23]), .C(n11) );
  BUFFD0 U44 ( .I(n14), .Z(n13) );
  BUFFD0 U45 ( .I(n15), .Z(n14) );
  BUFFD0 U46 ( .I(n16), .Z(n15) );
  BUFFD0 U47 ( .I(n17), .Z(n16) );
  BUFFD0 U48 ( .I(n18), .Z(n17) );
  BUFFD0 U49 ( .I(n19), .Z(n18) );
  BUFFD0 U50 ( .I(n20), .Z(n19) );
  BUFFD0 U51 ( .I(n21), .Z(n20) );
  BUFFD0 U52 ( .I(n22), .Z(n21) );
  BUFFD0 U53 ( .I(n23), .Z(n22) );
  BUFFD0 U54 ( .I(n24), .Z(n23) );
  BUFFD0 U55 ( .I(n25), .Z(n24) );
  BUFFD0 U56 ( .I(n26), .Z(n25) );
  BUFFD0 U57 ( .I(n27), .Z(n26) );
  BUFFD0 U58 ( .I(n28), .Z(n27) );
  BUFFD0 U59 ( .I(n29), .Z(n28) );
  BUFFD0 U60 ( .I(n30), .Z(n29) );
  BUFFD0 U61 ( .I(n31), .Z(n30) );
  BUFFD0 U62 ( .I(n32), .Z(n31) );
  BUFFD0 U63 ( .I(n33), .Z(n32) );
  BUFFD0 U64 ( .I(n34), .Z(n33) );
  BUFFD0 U65 ( .I(n35), .Z(n34) );
  BUFFD0 U66 ( .I(n36), .Z(n35) );
  BUFFD0 U67 ( .I(n37), .Z(n36) );
  BUFFD0 U68 ( .I(n38), .Z(n37) );
  BUFFD0 U69 ( .I(n39), .Z(n38) );
  BUFFD0 U70 ( .I(n40), .Z(n39) );
  BUFFD0 U71 ( .I(n41), .Z(n40) );
  BUFFD0 U72 ( .I(n42), .Z(n41) );
  BUFFD0 U73 ( .I(n43), .Z(n42) );
  BUFFD0 U74 ( .I(n44), .Z(n43) );
  BUFFD0 U75 ( .I(n45), .Z(n44) );
  BUFFD0 U76 ( .I(n46), .Z(n45) );
  BUFFD0 U77 ( .I(n47), .Z(n46) );
  BUFFD0 U78 ( .I(n48), .Z(n47) );
  BUFFD0 U79 ( .I(n49), .Z(n48) );
  BUFFD0 U80 ( .I(n50), .Z(n49) );
  BUFFD0 U81 ( .I(n51), .Z(n50) );
  BUFFD0 U82 ( .I(n52), .Z(n51) );
  BUFFD0 U83 ( .I(n53), .Z(n52) );
  BUFFD0 U84 ( .I(n54), .Z(n53) );
  BUFFD0 U85 ( .I(n55), .Z(n54) );
  BUFFD0 U86 ( .I(n56), .Z(n55) );
  BUFFD0 U87 ( .I(n57), .Z(n56) );
  BUFFD0 U88 ( .I(n58), .Z(n57) );
  BUFFD0 U89 ( .I(n59), .Z(n58) );
  BUFFD0 U90 ( .I(n60), .Z(n59) );
  BUFFD0 U91 ( .I(n61), .Z(n60) );
  BUFFD0 U92 ( .I(n63), .Z(n61) );
  INVD0 U93 ( .I(n62), .ZN(n63) );
  CKNXD16 U94 ( .I(n11), .ZN(n62) );
  BUFFD0 U95 ( .I(n3743), .Z(n64) );
  BUFFD0 U96 ( .I(n64), .Z(n65) );
  BUFFD0 U97 ( .I(n65), .Z(n94) );
  BUFFD0 U98 ( .I(n94), .Z(n95) );
  BUFFD0 U99 ( .I(n95), .Z(n96) );
  BUFFD0 U100 ( .I(n96), .Z(n97) );
  BUFFD0 U101 ( .I(n97), .Z(n98) );
  BUFFD0 U102 ( .I(n98), .Z(n99) );
  BUFFD0 U103 ( .I(n99), .Z(n100) );
  BUFFD0 U104 ( .I(n100), .Z(n101) );
  BUFFD0 U105 ( .I(n101), .Z(n102) );
  BUFFD0 U106 ( .I(n102), .Z(n103) );
  BUFFD0 U107 ( .I(n103), .Z(n104) );
  BUFFD0 U108 ( .I(n104), .Z(n105) );
  BUFFD0 U109 ( .I(n105), .Z(n106) );
  BUFFD0 U110 ( .I(n106), .Z(n107) );
  BUFFD0 U111 ( .I(n107), .Z(n108) );
  BUFFD0 U112 ( .I(n108), .Z(n109) );
  BUFFD0 U113 ( .I(n109), .Z(n110) );
  BUFFD0 U114 ( .I(n110), .Z(n111) );
  BUFFD0 U115 ( .I(n111), .Z(n112) );
  BUFFD0 U116 ( .I(n112), .Z(n113) );
  BUFFD0 U117 ( .I(n113), .Z(n114) );
  BUFFD0 U118 ( .I(n114), .Z(n115) );
  BUFFD0 U119 ( .I(n115), .Z(n116) );
  BUFFD0 U120 ( .I(n116), .Z(n117) );
  BUFFD0 U121 ( .I(n117), .Z(n118) );
  BUFFD0 U122 ( .I(n118), .Z(n119) );
  BUFFD0 U123 ( .I(n119), .Z(n120) );
  BUFFD0 U124 ( .I(n120), .Z(n121) );
  BUFFD0 U125 ( .I(n121), .Z(n122) );
  BUFFD0 U126 ( .I(n122), .Z(n123) );
  BUFFD0 U127 ( .I(n123), .Z(n124) );
  BUFFD0 U128 ( .I(n124), .Z(n125) );
  BUFFD0 U129 ( .I(n125), .Z(n126) );
  BUFFD0 U130 ( .I(n126), .Z(n127) );
  BUFFD0 U131 ( .I(n127), .Z(n128) );
  BUFFD0 U132 ( .I(n128), .Z(n129) );
  BUFFD0 U133 ( .I(n129), .Z(n130) );
  BUFFD0 U134 ( .I(n130), .Z(n131) );
  BUFFD0 U135 ( .I(n131), .Z(n132) );
  BUFFD0 U136 ( .I(n132), .Z(n133) );
  BUFFD0 U137 ( .I(n133), .Z(n134) );
  BUFFD0 U138 ( .I(n134), .Z(n135) );
  BUFFD0 U139 ( .I(n135), .Z(n136) );
  BUFFD0 U140 ( .I(n136), .Z(n137) );
  BUFFD0 U141 ( .I(n137), .Z(n138) );
  BUFFD0 U142 ( .I(n138), .Z(n139) );
  BUFFD0 U143 ( .I(n139), .Z(n140) );
  BUFFD0 U144 ( .I(n140), .Z(n141) );
  BUFFD0 U145 ( .I(n141), .Z(n142) );
  BUFFD0 U146 ( .I(n142), .Z(n143) );
  BUFFD0 U147 ( .I(n143), .Z(n144) );
  BUFFD0 U148 ( .I(n144), .Z(n145) );
  BUFFD0 U149 ( .I(n145), .Z(n146) );
  CKBD0 U150 ( .CLK(n146), .C(n147) );
  CKBD0 U151 ( .CLK(n3738), .C(n148) );
  BUFFD0 U152 ( .I(n148), .Z(n149) );
  BUFFD0 U153 ( .I(n149), .Z(n150) );
  BUFFD0 U154 ( .I(n150), .Z(n151) );
  BUFFD0 U155 ( .I(n151), .Z(n152) );
  BUFFD0 U156 ( .I(n152), .Z(n153) );
  BUFFD0 U157 ( .I(n153), .Z(n154) );
  BUFFD0 U158 ( .I(n154), .Z(n155) );
  BUFFD0 U159 ( .I(n155), .Z(n156) );
  BUFFD0 U160 ( .I(n156), .Z(n157) );
  BUFFD0 U161 ( .I(n157), .Z(n158) );
  BUFFD0 U162 ( .I(n158), .Z(n159) );
  BUFFD0 U163 ( .I(n159), .Z(n160) );
  BUFFD0 U164 ( .I(n160), .Z(n161) );
  BUFFD0 U165 ( .I(n161), .Z(n162) );
  BUFFD0 U166 ( .I(n162), .Z(n163) );
  BUFFD0 U167 ( .I(n163), .Z(n164) );
  BUFFD0 U168 ( .I(n164), .Z(n165) );
  BUFFD0 U169 ( .I(n165), .Z(n166) );
  BUFFD0 U170 ( .I(n166), .Z(n167) );
  BUFFD0 U171 ( .I(n167), .Z(n168) );
  BUFFD0 U172 ( .I(n168), .Z(n169) );
  BUFFD0 U173 ( .I(n169), .Z(n170) );
  BUFFD0 U174 ( .I(n170), .Z(n171) );
  BUFFD0 U175 ( .I(n171), .Z(n172) );
  BUFFD0 U176 ( .I(n172), .Z(n173) );
  BUFFD0 U177 ( .I(n173), .Z(n174) );
  BUFFD0 U178 ( .I(n174), .Z(n175) );
  BUFFD0 U179 ( .I(n175), .Z(n176) );
  BUFFD0 U180 ( .I(n176), .Z(n177) );
  BUFFD0 U181 ( .I(n177), .Z(n178) );
  BUFFD0 U182 ( .I(n178), .Z(n179) );
  BUFFD0 U183 ( .I(n179), .Z(n180) );
  BUFFD0 U184 ( .I(n180), .Z(n181) );
  BUFFD0 U185 ( .I(n181), .Z(n182) );
  BUFFD0 U186 ( .I(n182), .Z(n183) );
  BUFFD0 U187 ( .I(n183), .Z(n184) );
  BUFFD0 U188 ( .I(n184), .Z(n185) );
  BUFFD0 U189 ( .I(n185), .Z(n186) );
  BUFFD0 U190 ( .I(n186), .Z(n187) );
  BUFFD0 U191 ( .I(n187), .Z(n188) );
  BUFFD0 U192 ( .I(n188), .Z(n189) );
  BUFFD0 U193 ( .I(n189), .Z(n190) );
  BUFFD0 U194 ( .I(n190), .Z(n191) );
  BUFFD0 U195 ( .I(n191), .Z(n192) );
  BUFFD0 U196 ( .I(n192), .Z(n193) );
  BUFFD0 U197 ( .I(n193), .Z(n194) );
  BUFFD0 U198 ( .I(n194), .Z(n195) );
  BUFFD0 U199 ( .I(n195), .Z(n196) );
  BUFFD0 U200 ( .I(n196), .Z(n197) );
  BUFFD0 U201 ( .I(n197), .Z(n198) );
  BUFFD0 U202 ( .I(n198), .Z(n199) );
  BUFFD0 U203 ( .I(n199), .Z(n200) );
  BUFFD0 U204 ( .I(n200), .Z(n201) );
  BUFFD0 U205 ( .I(n201), .Z(n202) );
  CKBD0 U206 ( .CLK(n202), .C(n203) );
  CKBD0 U207 ( .CLK(DataI[16]), .C(n204) );
  BUFFD0 U208 ( .I(n207), .Z(n206) );
  BUFFD0 U209 ( .I(n208), .Z(n207) );
  BUFFD0 U210 ( .I(n209), .Z(n208) );
  BUFFD0 U211 ( .I(n210), .Z(n209) );
  BUFFD0 U212 ( .I(n211), .Z(n210) );
  BUFFD0 U213 ( .I(n212), .Z(n211) );
  BUFFD0 U214 ( .I(n213), .Z(n212) );
  BUFFD0 U215 ( .I(n214), .Z(n213) );
  BUFFD0 U216 ( .I(n215), .Z(n214) );
  BUFFD0 U217 ( .I(n216), .Z(n215) );
  BUFFD0 U218 ( .I(n217), .Z(n216) );
  BUFFD0 U219 ( .I(n218), .Z(n217) );
  BUFFD0 U220 ( .I(n219), .Z(n218) );
  BUFFD0 U221 ( .I(n220), .Z(n219) );
  BUFFD0 U222 ( .I(n221), .Z(n220) );
  BUFFD0 U223 ( .I(n222), .Z(n221) );
  BUFFD0 U224 ( .I(n223), .Z(n222) );
  BUFFD0 U225 ( .I(n224), .Z(n223) );
  BUFFD0 U226 ( .I(n225), .Z(n224) );
  BUFFD0 U227 ( .I(n226), .Z(n225) );
  BUFFD0 U228 ( .I(n227), .Z(n226) );
  BUFFD0 U229 ( .I(n228), .Z(n227) );
  BUFFD0 U230 ( .I(n229), .Z(n228) );
  BUFFD0 U231 ( .I(n230), .Z(n229) );
  BUFFD0 U232 ( .I(n231), .Z(n230) );
  BUFFD0 U233 ( .I(n232), .Z(n231) );
  BUFFD0 U234 ( .I(n233), .Z(n232) );
  BUFFD0 U235 ( .I(n234), .Z(n233) );
  BUFFD0 U236 ( .I(n235), .Z(n234) );
  BUFFD0 U237 ( .I(n236), .Z(n235) );
  BUFFD0 U238 ( .I(n237), .Z(n236) );
  BUFFD0 U239 ( .I(n238), .Z(n237) );
  BUFFD0 U240 ( .I(n239), .Z(n238) );
  BUFFD0 U241 ( .I(n240), .Z(n239) );
  BUFFD0 U242 ( .I(n241), .Z(n240) );
  BUFFD0 U243 ( .I(n242), .Z(n241) );
  BUFFD0 U244 ( .I(n243), .Z(n242) );
  BUFFD0 U245 ( .I(n244), .Z(n243) );
  BUFFD0 U246 ( .I(n245), .Z(n244) );
  BUFFD0 U247 ( .I(n246), .Z(n245) );
  BUFFD0 U248 ( .I(n247), .Z(n246) );
  BUFFD0 U249 ( .I(n248), .Z(n247) );
  BUFFD0 U250 ( .I(n249), .Z(n248) );
  BUFFD0 U251 ( .I(n250), .Z(n249) );
  BUFFD0 U252 ( .I(n251), .Z(n250) );
  BUFFD0 U253 ( .I(n252), .Z(n251) );
  BUFFD0 U254 ( .I(n253), .Z(n252) );
  BUFFD0 U255 ( .I(n254), .Z(n253) );
  BUFFD0 U256 ( .I(n256), .Z(n254) );
  INVD0 U257 ( .I(n255), .ZN(n256) );
  CKNXD16 U258 ( .I(n204), .ZN(n255) );
  BUFFD0 U259 ( .I(n3737), .Z(n257) );
  BUFFD0 U260 ( .I(n257), .Z(n258) );
  BUFFD0 U261 ( .I(n258), .Z(n259) );
  BUFFD0 U262 ( .I(n259), .Z(n260) );
  BUFFD0 U263 ( .I(n260), .Z(n261) );
  BUFFD0 U264 ( .I(n261), .Z(n262) );
  BUFFD0 U265 ( .I(n262), .Z(n263) );
  BUFFD0 U266 ( .I(n263), .Z(n264) );
  BUFFD0 U267 ( .I(n264), .Z(n265) );
  BUFFD0 U268 ( .I(n265), .Z(n266) );
  BUFFD0 U269 ( .I(n266), .Z(n267) );
  BUFFD0 U270 ( .I(n267), .Z(n268) );
  BUFFD0 U271 ( .I(n268), .Z(n269) );
  BUFFD0 U272 ( .I(n269), .Z(n270) );
  BUFFD0 U273 ( .I(n270), .Z(n271) );
  BUFFD0 U274 ( .I(n271), .Z(n272) );
  BUFFD0 U275 ( .I(n272), .Z(n273) );
  BUFFD0 U276 ( .I(n273), .Z(n274) );
  BUFFD0 U277 ( .I(n274), .Z(n275) );
  BUFFD0 U278 ( .I(n275), .Z(n276) );
  BUFFD0 U279 ( .I(n276), .Z(n277) );
  BUFFD0 U280 ( .I(n277), .Z(n278) );
  BUFFD0 U281 ( .I(n278), .Z(n279) );
  BUFFD0 U282 ( .I(n279), .Z(n280) );
  BUFFD0 U283 ( .I(n280), .Z(n281) );
  BUFFD0 U284 ( .I(n281), .Z(n282) );
  BUFFD0 U285 ( .I(n282), .Z(n283) );
  BUFFD0 U286 ( .I(n283), .Z(n284) );
  BUFFD0 U287 ( .I(n284), .Z(n285) );
  BUFFD0 U288 ( .I(n285), .Z(n286) );
  BUFFD0 U289 ( .I(n286), .Z(n287) );
  BUFFD0 U290 ( .I(n287), .Z(n288) );
  BUFFD0 U291 ( .I(n288), .Z(n289) );
  BUFFD0 U292 ( .I(n289), .Z(n290) );
  BUFFD0 U293 ( .I(n290), .Z(n291) );
  BUFFD0 U294 ( .I(n291), .Z(n292) );
  BUFFD0 U295 ( .I(n292), .Z(n293) );
  BUFFD0 U296 ( .I(n293), .Z(n294) );
  BUFFD0 U297 ( .I(n294), .Z(n295) );
  BUFFD0 U298 ( .I(n295), .Z(n296) );
  BUFFD0 U299 ( .I(n296), .Z(n297) );
  BUFFD0 U300 ( .I(n297), .Z(n298) );
  BUFFD0 U301 ( .I(n298), .Z(n299) );
  BUFFD0 U302 ( .I(n299), .Z(n300) );
  BUFFD0 U303 ( .I(n300), .Z(n301) );
  BUFFD0 U304 ( .I(n301), .Z(n302) );
  BUFFD0 U305 ( .I(n302), .Z(n303) );
  BUFFD0 U306 ( .I(n303), .Z(n304) );
  BUFFD0 U307 ( .I(n304), .Z(n305) );
  BUFFD0 U308 ( .I(n305), .Z(n306) );
  BUFFD0 U309 ( .I(n306), .Z(n307) );
  BUFFD0 U310 ( .I(n307), .Z(n308) );
  BUFFD0 U311 ( .I(n308), .Z(n309) );
  BUFFD0 U312 ( .I(n309), .Z(n310) );
  BUFFD0 U313 ( .I(n310), .Z(n311) );
  CKBD0 U314 ( .CLK(n311), .C(n312) );
  BUFFD0 U315 ( .I(n3736), .Z(n313) );
  BUFFD0 U316 ( .I(n313), .Z(n314) );
  BUFFD0 U317 ( .I(n314), .Z(n315) );
  BUFFD0 U318 ( .I(n315), .Z(n316) );
  BUFFD0 U319 ( .I(n316), .Z(n317) );
  BUFFD0 U320 ( .I(n317), .Z(n318) );
  BUFFD0 U321 ( .I(n318), .Z(n319) );
  BUFFD0 U322 ( .I(n319), .Z(n320) );
  BUFFD0 U323 ( .I(n320), .Z(n321) );
  BUFFD0 U324 ( .I(n321), .Z(n322) );
  BUFFD0 U325 ( .I(n322), .Z(n323) );
  BUFFD0 U326 ( .I(n323), .Z(n324) );
  BUFFD0 U327 ( .I(n324), .Z(n325) );
  BUFFD0 U328 ( .I(n325), .Z(n326) );
  BUFFD0 U329 ( .I(n326), .Z(n327) );
  BUFFD0 U330 ( .I(n327), .Z(n328) );
  BUFFD0 U331 ( .I(n328), .Z(n329) );
  BUFFD0 U332 ( .I(n329), .Z(n330) );
  BUFFD0 U333 ( .I(n330), .Z(n331) );
  BUFFD0 U334 ( .I(n331), .Z(n332) );
  BUFFD0 U335 ( .I(n332), .Z(n333) );
  BUFFD0 U336 ( .I(n333), .Z(n334) );
  BUFFD0 U337 ( .I(n334), .Z(n335) );
  BUFFD0 U338 ( .I(n335), .Z(n336) );
  BUFFD0 U339 ( .I(n336), .Z(n337) );
  BUFFD0 U340 ( .I(n337), .Z(n338) );
  BUFFD0 U341 ( .I(n338), .Z(n339) );
  BUFFD0 U342 ( .I(n339), .Z(n340) );
  BUFFD0 U343 ( .I(n340), .Z(n341) );
  BUFFD0 U344 ( .I(n341), .Z(n342) );
  BUFFD0 U345 ( .I(n342), .Z(n343) );
  BUFFD0 U346 ( .I(n343), .Z(n344) );
  BUFFD0 U347 ( .I(n344), .Z(n345) );
  BUFFD0 U348 ( .I(n345), .Z(n346) );
  BUFFD0 U349 ( .I(n346), .Z(n347) );
  BUFFD0 U350 ( .I(n347), .Z(n348) );
  BUFFD0 U351 ( .I(n348), .Z(n349) );
  BUFFD0 U352 ( .I(n349), .Z(n350) );
  BUFFD0 U353 ( .I(n350), .Z(n351) );
  BUFFD0 U354 ( .I(n351), .Z(n352) );
  BUFFD0 U355 ( .I(n352), .Z(n353) );
  BUFFD0 U356 ( .I(n353), .Z(n354) );
  BUFFD0 U357 ( .I(n354), .Z(n355) );
  BUFFD0 U358 ( .I(n355), .Z(n356) );
  BUFFD0 U359 ( .I(n356), .Z(n357) );
  BUFFD0 U360 ( .I(n357), .Z(n358) );
  BUFFD0 U361 ( .I(n358), .Z(n359) );
  BUFFD0 U362 ( .I(n359), .Z(n360) );
  BUFFD0 U363 ( .I(n360), .Z(n361) );
  BUFFD0 U364 ( .I(n361), .Z(n362) );
  BUFFD0 U365 ( .I(n362), .Z(n363) );
  BUFFD0 U366 ( .I(n363), .Z(n364) );
  BUFFD0 U367 ( .I(n364), .Z(n365) );
  BUFFD0 U368 ( .I(n365), .Z(n366) );
  BUFFD0 U369 ( .I(n366), .Z(n367) );
  CKBD0 U370 ( .CLK(n367), .C(n368) );
  CKBD0 U371 ( .CLK(DataI[13]), .C(n369) );
  BUFFD0 U372 ( .I(n372), .Z(n371) );
  BUFFD0 U373 ( .I(n373), .Z(n372) );
  BUFFD0 U374 ( .I(n374), .Z(n373) );
  BUFFD0 U375 ( .I(n375), .Z(n374) );
  BUFFD0 U376 ( .I(n376), .Z(n375) );
  BUFFD0 U377 ( .I(n377), .Z(n376) );
  BUFFD0 U378 ( .I(n378), .Z(n377) );
  BUFFD0 U379 ( .I(n379), .Z(n378) );
  BUFFD0 U380 ( .I(n380), .Z(n379) );
  BUFFD0 U381 ( .I(n381), .Z(n380) );
  BUFFD0 U382 ( .I(n382), .Z(n381) );
  BUFFD0 U383 ( .I(n383), .Z(n382) );
  BUFFD0 U384 ( .I(n384), .Z(n383) );
  BUFFD0 U385 ( .I(n385), .Z(n384) );
  BUFFD0 U386 ( .I(n386), .Z(n385) );
  BUFFD0 U387 ( .I(n387), .Z(n386) );
  BUFFD0 U388 ( .I(n388), .Z(n387) );
  BUFFD0 U389 ( .I(n389), .Z(n388) );
  BUFFD0 U390 ( .I(n390), .Z(n389) );
  BUFFD0 U391 ( .I(n391), .Z(n390) );
  BUFFD0 U392 ( .I(n392), .Z(n391) );
  BUFFD0 U393 ( .I(n393), .Z(n392) );
  BUFFD0 U394 ( .I(n394), .Z(n393) );
  BUFFD0 U395 ( .I(n395), .Z(n394) );
  BUFFD0 U396 ( .I(n396), .Z(n395) );
  BUFFD0 U397 ( .I(n397), .Z(n396) );
  BUFFD0 U398 ( .I(n398), .Z(n397) );
  BUFFD0 U399 ( .I(n399), .Z(n398) );
  BUFFD0 U400 ( .I(n400), .Z(n399) );
  BUFFD0 U401 ( .I(n401), .Z(n400) );
  BUFFD0 U402 ( .I(n402), .Z(n401) );
  BUFFD0 U403 ( .I(n403), .Z(n402) );
  BUFFD0 U404 ( .I(n404), .Z(n403) );
  BUFFD0 U405 ( .I(n405), .Z(n404) );
  BUFFD0 U406 ( .I(n406), .Z(n405) );
  BUFFD0 U407 ( .I(n407), .Z(n406) );
  BUFFD0 U408 ( .I(n408), .Z(n407) );
  BUFFD0 U409 ( .I(n409), .Z(n408) );
  BUFFD0 U410 ( .I(n410), .Z(n409) );
  BUFFD0 U411 ( .I(n411), .Z(n410) );
  BUFFD0 U412 ( .I(n412), .Z(n411) );
  BUFFD0 U413 ( .I(n413), .Z(n412) );
  BUFFD0 U414 ( .I(n414), .Z(n413) );
  BUFFD0 U415 ( .I(n415), .Z(n414) );
  BUFFD0 U416 ( .I(n416), .Z(n415) );
  BUFFD0 U417 ( .I(n417), .Z(n416) );
  BUFFD0 U418 ( .I(n418), .Z(n417) );
  BUFFD0 U419 ( .I(n419), .Z(n418) );
  BUFFD0 U420 ( .I(n421), .Z(n419) );
  INVD0 U421 ( .I(n420), .ZN(n421) );
  CKNXD16 U422 ( .I(n369), .ZN(n420) );
  CKBD0 U423 ( .CLK(DataI[12]), .C(n422) );
  BUFFD0 U424 ( .I(n425), .Z(n424) );
  BUFFD0 U425 ( .I(n426), .Z(n425) );
  BUFFD0 U426 ( .I(n427), .Z(n426) );
  BUFFD0 U427 ( .I(n428), .Z(n427) );
  BUFFD0 U428 ( .I(n429), .Z(n428) );
  BUFFD0 U429 ( .I(n430), .Z(n429) );
  BUFFD0 U430 ( .I(n431), .Z(n430) );
  BUFFD0 U431 ( .I(n432), .Z(n431) );
  BUFFD0 U432 ( .I(n433), .Z(n432) );
  BUFFD0 U433 ( .I(n434), .Z(n433) );
  BUFFD0 U434 ( .I(n435), .Z(n434) );
  BUFFD0 U435 ( .I(n436), .Z(n435) );
  BUFFD0 U436 ( .I(n437), .Z(n436) );
  BUFFD0 U437 ( .I(n438), .Z(n437) );
  BUFFD0 U438 ( .I(n439), .Z(n438) );
  BUFFD0 U439 ( .I(n440), .Z(n439) );
  BUFFD0 U440 ( .I(n441), .Z(n440) );
  BUFFD0 U441 ( .I(n442), .Z(n441) );
  BUFFD0 U442 ( .I(n443), .Z(n442) );
  BUFFD0 U443 ( .I(n444), .Z(n443) );
  BUFFD0 U444 ( .I(n445), .Z(n444) );
  BUFFD0 U445 ( .I(n446), .Z(n445) );
  BUFFD0 U446 ( .I(n447), .Z(n446) );
  BUFFD0 U447 ( .I(n448), .Z(n447) );
  BUFFD0 U448 ( .I(n449), .Z(n448) );
  BUFFD0 U449 ( .I(n450), .Z(n449) );
  BUFFD0 U450 ( .I(n451), .Z(n450) );
  BUFFD0 U451 ( .I(n452), .Z(n451) );
  BUFFD0 U452 ( .I(n453), .Z(n452) );
  BUFFD0 U453 ( .I(n454), .Z(n453) );
  BUFFD0 U454 ( .I(n455), .Z(n454) );
  BUFFD0 U455 ( .I(n456), .Z(n455) );
  BUFFD0 U456 ( .I(n457), .Z(n456) );
  BUFFD0 U457 ( .I(n458), .Z(n457) );
  BUFFD0 U458 ( .I(n459), .Z(n458) );
  BUFFD0 U459 ( .I(n460), .Z(n459) );
  BUFFD0 U460 ( .I(n461), .Z(n460) );
  BUFFD0 U461 ( .I(n462), .Z(n461) );
  BUFFD0 U462 ( .I(n463), .Z(n462) );
  BUFFD0 U463 ( .I(n464), .Z(n463) );
  BUFFD0 U464 ( .I(n465), .Z(n464) );
  BUFFD0 U465 ( .I(n466), .Z(n465) );
  BUFFD0 U466 ( .I(n467), .Z(n466) );
  BUFFD0 U467 ( .I(n468), .Z(n467) );
  BUFFD0 U468 ( .I(n469), .Z(n468) );
  BUFFD0 U469 ( .I(n470), .Z(n469) );
  BUFFD0 U470 ( .I(n471), .Z(n470) );
  BUFFD0 U471 ( .I(n472), .Z(n471) );
  BUFFD0 U472 ( .I(n474), .Z(n472) );
  INVD0 U473 ( .I(n473), .ZN(n474) );
  CKNXD16 U474 ( .I(n422), .ZN(n473) );
  CKBD0 U475 ( .CLK(n3735), .C(n475) );
  BUFFD0 U476 ( .I(n475), .Z(n476) );
  BUFFD0 U477 ( .I(n476), .Z(n477) );
  BUFFD0 U478 ( .I(n477), .Z(n478) );
  BUFFD0 U479 ( .I(n478), .Z(n479) );
  BUFFD0 U480 ( .I(n479), .Z(n480) );
  BUFFD0 U481 ( .I(n480), .Z(n481) );
  BUFFD0 U482 ( .I(n481), .Z(n482) );
  BUFFD0 U483 ( .I(n482), .Z(n483) );
  BUFFD0 U484 ( .I(n483), .Z(n484) );
  BUFFD0 U485 ( .I(n484), .Z(n485) );
  BUFFD0 U486 ( .I(n485), .Z(n486) );
  BUFFD0 U487 ( .I(n486), .Z(n487) );
  BUFFD0 U488 ( .I(n487), .Z(n488) );
  BUFFD0 U489 ( .I(n488), .Z(n489) );
  BUFFD0 U490 ( .I(n489), .Z(n490) );
  BUFFD0 U491 ( .I(n490), .Z(n491) );
  BUFFD0 U492 ( .I(n491), .Z(n492) );
  BUFFD0 U493 ( .I(n492), .Z(n493) );
  BUFFD0 U494 ( .I(n493), .Z(n494) );
  BUFFD0 U495 ( .I(n494), .Z(n495) );
  BUFFD0 U496 ( .I(n495), .Z(n496) );
  BUFFD0 U497 ( .I(n496), .Z(n497) );
  BUFFD0 U498 ( .I(n497), .Z(n498) );
  BUFFD0 U499 ( .I(n498), .Z(n499) );
  BUFFD0 U500 ( .I(n499), .Z(n500) );
  BUFFD0 U501 ( .I(n500), .Z(n501) );
  BUFFD0 U502 ( .I(n501), .Z(n502) );
  BUFFD0 U503 ( .I(n502), .Z(n503) );
  BUFFD0 U504 ( .I(n503), .Z(n504) );
  BUFFD0 U505 ( .I(n504), .Z(n505) );
  BUFFD0 U506 ( .I(n505), .Z(n506) );
  BUFFD0 U507 ( .I(n506), .Z(n507) );
  BUFFD0 U508 ( .I(n507), .Z(n508) );
  BUFFD0 U509 ( .I(n508), .Z(n509) );
  BUFFD0 U510 ( .I(n509), .Z(n510) );
  BUFFD0 U511 ( .I(n510), .Z(n511) );
  BUFFD0 U512 ( .I(n511), .Z(n512) );
  BUFFD0 U513 ( .I(n512), .Z(n513) );
  BUFFD0 U514 ( .I(n513), .Z(n514) );
  BUFFD0 U515 ( .I(n514), .Z(n515) );
  BUFFD0 U516 ( .I(n515), .Z(n516) );
  BUFFD0 U517 ( .I(n516), .Z(n517) );
  BUFFD0 U518 ( .I(n517), .Z(n518) );
  BUFFD0 U519 ( .I(n518), .Z(n519) );
  BUFFD0 U520 ( .I(n519), .Z(n520) );
  BUFFD0 U521 ( .I(n520), .Z(n521) );
  BUFFD0 U522 ( .I(n521), .Z(n522) );
  BUFFD0 U523 ( .I(n522), .Z(n523) );
  BUFFD0 U524 ( .I(n523), .Z(n524) );
  BUFFD0 U525 ( .I(n524), .Z(n525) );
  BUFFD0 U526 ( .I(n525), .Z(n526) );
  BUFFD0 U527 ( .I(n526), .Z(n527) );
  BUFFD0 U528 ( .I(n527), .Z(n528) );
  BUFFD0 U529 ( .I(n528), .Z(n529) );
  CKBD0 U530 ( .CLK(n529), .C(n530) );
  CKBD0 U531 ( .CLK(n3734), .C(n531) );
  BUFFD0 U532 ( .I(n531), .Z(n532) );
  BUFFD0 U533 ( .I(n532), .Z(n533) );
  BUFFD0 U534 ( .I(n533), .Z(n534) );
  BUFFD0 U535 ( .I(n534), .Z(n535) );
  BUFFD0 U536 ( .I(n535), .Z(n536) );
  BUFFD0 U537 ( .I(n536), .Z(n537) );
  BUFFD0 U538 ( .I(n537), .Z(n538) );
  BUFFD0 U539 ( .I(n538), .Z(n539) );
  BUFFD0 U540 ( .I(n539), .Z(n540) );
  BUFFD0 U541 ( .I(n540), .Z(n541) );
  BUFFD0 U542 ( .I(n541), .Z(n542) );
  BUFFD0 U543 ( .I(n542), .Z(n543) );
  BUFFD0 U544 ( .I(n543), .Z(n544) );
  BUFFD0 U545 ( .I(n544), .Z(n545) );
  BUFFD0 U546 ( .I(n545), .Z(n546) );
  BUFFD0 U547 ( .I(n546), .Z(n547) );
  BUFFD0 U548 ( .I(n547), .Z(n548) );
  BUFFD0 U549 ( .I(n548), .Z(n549) );
  BUFFD0 U550 ( .I(n549), .Z(n550) );
  BUFFD0 U551 ( .I(n550), .Z(n551) );
  BUFFD0 U552 ( .I(n551), .Z(n552) );
  BUFFD0 U553 ( .I(n552), .Z(n553) );
  BUFFD0 U554 ( .I(n553), .Z(n554) );
  BUFFD0 U555 ( .I(n554), .Z(n555) );
  BUFFD0 U556 ( .I(n555), .Z(n556) );
  BUFFD0 U557 ( .I(n556), .Z(n557) );
  BUFFD0 U558 ( .I(n557), .Z(n558) );
  BUFFD0 U559 ( .I(n558), .Z(n559) );
  BUFFD0 U560 ( .I(n559), .Z(n560) );
  BUFFD0 U561 ( .I(n560), .Z(n561) );
  BUFFD0 U562 ( .I(n561), .Z(n562) );
  BUFFD0 U563 ( .I(n562), .Z(n563) );
  BUFFD0 U564 ( .I(n563), .Z(n564) );
  BUFFD0 U565 ( .I(n564), .Z(n565) );
  BUFFD0 U566 ( .I(n565), .Z(n566) );
  BUFFD0 U567 ( .I(n566), .Z(n567) );
  BUFFD0 U568 ( .I(n567), .Z(n568) );
  BUFFD0 U569 ( .I(n568), .Z(n569) );
  BUFFD0 U570 ( .I(n569), .Z(n570) );
  BUFFD0 U571 ( .I(n570), .Z(n571) );
  BUFFD0 U572 ( .I(n571), .Z(n572) );
  BUFFD0 U573 ( .I(n572), .Z(n573) );
  BUFFD0 U574 ( .I(n573), .Z(n574) );
  BUFFD0 U575 ( .I(n574), .Z(n575) );
  BUFFD0 U576 ( .I(n575), .Z(n576) );
  BUFFD0 U577 ( .I(n576), .Z(n577) );
  BUFFD0 U578 ( .I(n577), .Z(n578) );
  BUFFD0 U579 ( .I(n578), .Z(n579) );
  BUFFD0 U580 ( .I(n579), .Z(n580) );
  BUFFD0 U581 ( .I(n580), .Z(n581) );
  BUFFD0 U582 ( .I(n581), .Z(n582) );
  BUFFD0 U583 ( .I(n582), .Z(n583) );
  BUFFD0 U584 ( .I(n583), .Z(n584) );
  BUFFD0 U585 ( .I(n584), .Z(n585) );
  CKBD0 U586 ( .CLK(n585), .C(n586) );
  INVD0 U587 ( .I(n587), .ZN(n588) );
  INVD16 U588 ( .I(DataI[9]), .ZN(n587) );
  BUFFD0 U589 ( .I(n591), .Z(n590) );
  BUFFD0 U590 ( .I(n592), .Z(n591) );
  BUFFD0 U591 ( .I(n593), .Z(n592) );
  BUFFD0 U592 ( .I(n594), .Z(n593) );
  BUFFD0 U593 ( .I(n595), .Z(n594) );
  BUFFD0 U594 ( .I(n596), .Z(n595) );
  BUFFD0 U595 ( .I(n597), .Z(n596) );
  BUFFD0 U596 ( .I(n598), .Z(n597) );
  BUFFD0 U597 ( .I(n599), .Z(n598) );
  BUFFD0 U598 ( .I(n600), .Z(n599) );
  BUFFD0 U599 ( .I(n601), .Z(n600) );
  BUFFD0 U600 ( .I(n602), .Z(n601) );
  BUFFD0 U601 ( .I(n603), .Z(n602) );
  BUFFD0 U602 ( .I(n604), .Z(n603) );
  BUFFD0 U603 ( .I(n605), .Z(n604) );
  BUFFD0 U604 ( .I(n606), .Z(n605) );
  BUFFD0 U605 ( .I(n607), .Z(n606) );
  BUFFD0 U606 ( .I(n608), .Z(n607) );
  BUFFD0 U607 ( .I(n609), .Z(n608) );
  BUFFD0 U608 ( .I(n610), .Z(n609) );
  BUFFD0 U609 ( .I(n611), .Z(n610) );
  BUFFD0 U610 ( .I(n612), .Z(n611) );
  BUFFD0 U611 ( .I(n613), .Z(n612) );
  BUFFD0 U612 ( .I(n614), .Z(n613) );
  BUFFD0 U613 ( .I(n615), .Z(n614) );
  BUFFD0 U614 ( .I(n616), .Z(n615) );
  BUFFD0 U615 ( .I(n617), .Z(n616) );
  BUFFD0 U616 ( .I(n618), .Z(n617) );
  BUFFD0 U617 ( .I(n619), .Z(n618) );
  BUFFD0 U618 ( .I(n620), .Z(n619) );
  BUFFD0 U619 ( .I(n621), .Z(n620) );
  BUFFD0 U620 ( .I(n622), .Z(n621) );
  BUFFD0 U621 ( .I(n623), .Z(n622) );
  BUFFD0 U622 ( .I(n624), .Z(n623) );
  BUFFD0 U623 ( .I(n625), .Z(n624) );
  BUFFD0 U624 ( .I(n626), .Z(n625) );
  BUFFD0 U625 ( .I(n627), .Z(n626) );
  BUFFD0 U626 ( .I(n628), .Z(n627) );
  BUFFD0 U627 ( .I(n629), .Z(n628) );
  BUFFD0 U628 ( .I(n630), .Z(n629) );
  BUFFD0 U629 ( .I(n631), .Z(n630) );
  BUFFD0 U630 ( .I(n632), .Z(n631) );
  BUFFD0 U631 ( .I(n633), .Z(n632) );
  BUFFD0 U632 ( .I(n634), .Z(n633) );
  BUFFD0 U633 ( .I(n635), .Z(n634) );
  BUFFD0 U634 ( .I(n636), .Z(n635) );
  BUFFD0 U635 ( .I(n637), .Z(n636) );
  BUFFD0 U636 ( .I(n638), .Z(n637) );
  BUFFD0 U637 ( .I(n640), .Z(n638) );
  INVD0 U638 ( .I(n639), .ZN(n640) );
  CKNXD16 U639 ( .I(n588), .ZN(n639) );
  BUFFD0 U640 ( .I(n3733), .Z(n641) );
  BUFFD0 U641 ( .I(n641), .Z(n642) );
  BUFFD0 U642 ( .I(n642), .Z(n643) );
  BUFFD0 U643 ( .I(n643), .Z(n644) );
  BUFFD0 U644 ( .I(n644), .Z(n645) );
  BUFFD0 U645 ( .I(n645), .Z(n646) );
  BUFFD0 U646 ( .I(n646), .Z(n647) );
  BUFFD0 U647 ( .I(n647), .Z(n648) );
  BUFFD0 U648 ( .I(n648), .Z(n649) );
  BUFFD0 U649 ( .I(n649), .Z(n650) );
  BUFFD0 U650 ( .I(n650), .Z(n651) );
  BUFFD0 U651 ( .I(n651), .Z(n652) );
  BUFFD0 U652 ( .I(n652), .Z(n653) );
  BUFFD0 U653 ( .I(n653), .Z(n654) );
  BUFFD0 U654 ( .I(n654), .Z(n655) );
  BUFFD0 U655 ( .I(n655), .Z(n656) );
  BUFFD0 U656 ( .I(n656), .Z(n657) );
  BUFFD0 U657 ( .I(n657), .Z(n658) );
  BUFFD0 U658 ( .I(n658), .Z(n659) );
  BUFFD0 U659 ( .I(n659), .Z(n660) );
  BUFFD0 U660 ( .I(n660), .Z(n661) );
  BUFFD0 U661 ( .I(n661), .Z(n662) );
  BUFFD0 U662 ( .I(n662), .Z(n663) );
  BUFFD0 U663 ( .I(n663), .Z(n664) );
  BUFFD0 U664 ( .I(n664), .Z(n665) );
  BUFFD0 U665 ( .I(n665), .Z(n666) );
  BUFFD0 U666 ( .I(n666), .Z(n667) );
  BUFFD0 U667 ( .I(n667), .Z(n668) );
  BUFFD0 U668 ( .I(n668), .Z(n669) );
  BUFFD0 U669 ( .I(n669), .Z(n670) );
  BUFFD0 U670 ( .I(n670), .Z(n671) );
  BUFFD0 U671 ( .I(n671), .Z(n672) );
  BUFFD0 U672 ( .I(n672), .Z(n673) );
  BUFFD0 U673 ( .I(n673), .Z(n674) );
  BUFFD0 U674 ( .I(n674), .Z(n675) );
  BUFFD0 U675 ( .I(n675), .Z(n676) );
  BUFFD0 U676 ( .I(n676), .Z(n677) );
  BUFFD0 U677 ( .I(n677), .Z(n678) );
  BUFFD0 U678 ( .I(n678), .Z(n679) );
  BUFFD0 U679 ( .I(n679), .Z(n680) );
  BUFFD0 U680 ( .I(n680), .Z(n681) );
  BUFFD0 U681 ( .I(n681), .Z(n682) );
  BUFFD0 U682 ( .I(n682), .Z(n683) );
  BUFFD0 U683 ( .I(n683), .Z(n684) );
  BUFFD0 U684 ( .I(n684), .Z(n685) );
  BUFFD0 U685 ( .I(n685), .Z(n686) );
  BUFFD0 U686 ( .I(n686), .Z(n687) );
  BUFFD0 U687 ( .I(n687), .Z(n688) );
  BUFFD0 U688 ( .I(n688), .Z(n689) );
  BUFFD0 U689 ( .I(n689), .Z(n690) );
  BUFFD0 U690 ( .I(n690), .Z(n691) );
  BUFFD0 U691 ( .I(n691), .Z(n692) );
  BUFFD0 U692 ( .I(n692), .Z(n693) );
  BUFFD0 U693 ( .I(n693), .Z(n694) );
  BUFFD0 U694 ( .I(n694), .Z(n695) );
  CKBD0 U695 ( .CLK(n695), .C(n696) );
  BUFFD0 U696 ( .I(n3732), .Z(n697) );
  BUFFD0 U697 ( .I(n697), .Z(n698) );
  BUFFD0 U698 ( .I(n698), .Z(n699) );
  BUFFD0 U699 ( .I(n699), .Z(n700) );
  BUFFD0 U700 ( .I(n700), .Z(n701) );
  BUFFD0 U701 ( .I(n701), .Z(n702) );
  BUFFD0 U702 ( .I(n702), .Z(n703) );
  BUFFD0 U703 ( .I(n703), .Z(n704) );
  BUFFD0 U704 ( .I(n704), .Z(n705) );
  BUFFD0 U705 ( .I(n705), .Z(n706) );
  BUFFD0 U706 ( .I(n706), .Z(n707) );
  BUFFD0 U707 ( .I(n707), .Z(n708) );
  BUFFD0 U708 ( .I(n708), .Z(n709) );
  BUFFD0 U709 ( .I(n709), .Z(n710) );
  BUFFD0 U710 ( .I(n710), .Z(n711) );
  BUFFD0 U711 ( .I(n711), .Z(n712) );
  BUFFD0 U712 ( .I(n712), .Z(n713) );
  BUFFD0 U713 ( .I(n713), .Z(n714) );
  BUFFD0 U714 ( .I(n714), .Z(n715) );
  BUFFD0 U715 ( .I(n715), .Z(n716) );
  BUFFD0 U716 ( .I(n716), .Z(n717) );
  BUFFD0 U717 ( .I(n717), .Z(n718) );
  BUFFD0 U718 ( .I(n718), .Z(n719) );
  BUFFD0 U719 ( .I(n719), .Z(n720) );
  BUFFD0 U720 ( .I(n720), .Z(n721) );
  BUFFD0 U721 ( .I(n721), .Z(n722) );
  BUFFD0 U722 ( .I(n722), .Z(n723) );
  BUFFD0 U723 ( .I(n723), .Z(n724) );
  BUFFD0 U724 ( .I(n724), .Z(n725) );
  BUFFD0 U725 ( .I(n725), .Z(n726) );
  BUFFD0 U726 ( .I(n726), .Z(n727) );
  BUFFD0 U727 ( .I(n727), .Z(n728) );
  BUFFD0 U728 ( .I(n728), .Z(n729) );
  BUFFD0 U729 ( .I(n729), .Z(n730) );
  BUFFD0 U730 ( .I(n730), .Z(n731) );
  BUFFD0 U731 ( .I(n731), .Z(n732) );
  BUFFD0 U732 ( .I(n732), .Z(n733) );
  BUFFD0 U733 ( .I(n733), .Z(n734) );
  BUFFD0 U734 ( .I(n734), .Z(n735) );
  BUFFD0 U735 ( .I(n735), .Z(n736) );
  BUFFD0 U736 ( .I(n736), .Z(n737) );
  BUFFD0 U737 ( .I(n737), .Z(n738) );
  BUFFD0 U738 ( .I(n738), .Z(n739) );
  BUFFD0 U739 ( .I(n739), .Z(n740) );
  BUFFD0 U740 ( .I(n740), .Z(n741) );
  BUFFD0 U741 ( .I(n741), .Z(n742) );
  BUFFD0 U742 ( .I(n742), .Z(n743) );
  BUFFD0 U743 ( .I(n743), .Z(n744) );
  BUFFD0 U744 ( .I(n744), .Z(n745) );
  BUFFD0 U745 ( .I(n745), .Z(n746) );
  BUFFD0 U746 ( .I(n746), .Z(n747) );
  BUFFD0 U747 ( .I(n747), .Z(n748) );
  BUFFD0 U748 ( .I(n748), .Z(n749) );
  BUFFD0 U749 ( .I(n749), .Z(n750) );
  BUFFD0 U750 ( .I(n750), .Z(n751) );
  CKBD0 U751 ( .CLK(n751), .C(n752) );
  CKBD0 U752 ( .CLK(n3731), .C(n753) );
  CKBD12 U753 ( .CLK(DataI[6]), .C(n3731) );
  BUFFD0 U754 ( .I(n756), .Z(n755) );
  BUFFD0 U755 ( .I(n757), .Z(n756) );
  BUFFD0 U756 ( .I(n758), .Z(n757) );
  BUFFD0 U757 ( .I(n759), .Z(n758) );
  BUFFD0 U758 ( .I(n760), .Z(n759) );
  BUFFD0 U759 ( .I(n761), .Z(n760) );
  BUFFD0 U760 ( .I(n762), .Z(n761) );
  BUFFD0 U761 ( .I(n763), .Z(n762) );
  BUFFD0 U762 ( .I(n764), .Z(n763) );
  BUFFD0 U763 ( .I(n765), .Z(n764) );
  BUFFD0 U764 ( .I(n766), .Z(n765) );
  BUFFD0 U765 ( .I(n767), .Z(n766) );
  BUFFD0 U766 ( .I(n768), .Z(n767) );
  BUFFD0 U767 ( .I(n769), .Z(n768) );
  BUFFD0 U768 ( .I(n770), .Z(n769) );
  BUFFD0 U769 ( .I(n771), .Z(n770) );
  BUFFD0 U770 ( .I(n772), .Z(n771) );
  BUFFD0 U771 ( .I(n773), .Z(n772) );
  BUFFD0 U772 ( .I(n774), .Z(n773) );
  BUFFD0 U773 ( .I(n775), .Z(n774) );
  BUFFD0 U774 ( .I(n776), .Z(n775) );
  BUFFD0 U775 ( .I(n777), .Z(n776) );
  BUFFD0 U776 ( .I(n778), .Z(n777) );
  BUFFD0 U777 ( .I(n779), .Z(n778) );
  BUFFD0 U778 ( .I(n780), .Z(n779) );
  BUFFD0 U779 ( .I(n781), .Z(n780) );
  BUFFD0 U780 ( .I(n782), .Z(n781) );
  BUFFD0 U781 ( .I(n783), .Z(n782) );
  BUFFD0 U782 ( .I(n784), .Z(n783) );
  BUFFD0 U783 ( .I(n785), .Z(n784) );
  BUFFD0 U784 ( .I(n786), .Z(n785) );
  BUFFD0 U785 ( .I(n787), .Z(n786) );
  BUFFD0 U786 ( .I(n788), .Z(n787) );
  BUFFD0 U787 ( .I(n789), .Z(n788) );
  BUFFD0 U788 ( .I(n790), .Z(n789) );
  BUFFD0 U789 ( .I(n791), .Z(n790) );
  BUFFD0 U790 ( .I(n792), .Z(n791) );
  BUFFD0 U791 ( .I(n793), .Z(n792) );
  BUFFD0 U792 ( .I(n794), .Z(n793) );
  BUFFD0 U793 ( .I(n795), .Z(n794) );
  BUFFD0 U794 ( .I(n796), .Z(n795) );
  BUFFD0 U795 ( .I(n797), .Z(n796) );
  BUFFD0 U796 ( .I(n798), .Z(n797) );
  BUFFD0 U797 ( .I(n799), .Z(n798) );
  BUFFD0 U798 ( .I(n800), .Z(n799) );
  BUFFD0 U799 ( .I(n801), .Z(n800) );
  BUFFD0 U800 ( .I(n802), .Z(n801) );
  BUFFD0 U801 ( .I(n804), .Z(n802) );
  INVD0 U802 ( .I(n803), .ZN(n804) );
  CKNXD16 U803 ( .I(n753), .ZN(n803) );
  INVD0 U804 ( .I(n805), .ZN(n806) );
  INVD16 U805 ( .I(DataI[5]), .ZN(n805) );
  BUFFD0 U806 ( .I(n809), .Z(n808) );
  BUFFD0 U807 ( .I(n810), .Z(n809) );
  BUFFD0 U808 ( .I(n811), .Z(n810) );
  BUFFD0 U809 ( .I(n812), .Z(n811) );
  BUFFD0 U810 ( .I(n813), .Z(n812) );
  BUFFD0 U811 ( .I(n814), .Z(n813) );
  BUFFD0 U812 ( .I(n815), .Z(n814) );
  BUFFD0 U813 ( .I(n816), .Z(n815) );
  BUFFD0 U814 ( .I(n817), .Z(n816) );
  BUFFD0 U815 ( .I(n818), .Z(n817) );
  BUFFD0 U816 ( .I(n819), .Z(n818) );
  BUFFD0 U817 ( .I(n820), .Z(n819) );
  BUFFD0 U818 ( .I(n821), .Z(n820) );
  BUFFD0 U819 ( .I(n822), .Z(n821) );
  BUFFD0 U820 ( .I(n823), .Z(n822) );
  BUFFD0 U821 ( .I(n824), .Z(n823) );
  BUFFD0 U822 ( .I(n825), .Z(n824) );
  BUFFD0 U823 ( .I(n826), .Z(n825) );
  BUFFD0 U824 ( .I(n827), .Z(n826) );
  BUFFD0 U825 ( .I(n828), .Z(n827) );
  BUFFD0 U826 ( .I(n829), .Z(n828) );
  BUFFD0 U827 ( .I(n830), .Z(n829) );
  BUFFD0 U828 ( .I(n831), .Z(n830) );
  BUFFD0 U829 ( .I(n832), .Z(n831) );
  BUFFD0 U830 ( .I(n833), .Z(n832) );
  BUFFD0 U831 ( .I(n834), .Z(n833) );
  BUFFD0 U832 ( .I(n835), .Z(n834) );
  BUFFD0 U833 ( .I(n836), .Z(n835) );
  BUFFD0 U834 ( .I(n837), .Z(n836) );
  BUFFD0 U835 ( .I(n838), .Z(n837) );
  BUFFD0 U836 ( .I(n839), .Z(n838) );
  BUFFD0 U837 ( .I(n840), .Z(n839) );
  BUFFD0 U838 ( .I(n841), .Z(n840) );
  BUFFD0 U839 ( .I(n842), .Z(n841) );
  BUFFD0 U840 ( .I(n843), .Z(n842) );
  BUFFD0 U841 ( .I(n844), .Z(n843) );
  BUFFD0 U842 ( .I(n845), .Z(n844) );
  BUFFD0 U843 ( .I(n846), .Z(n845) );
  BUFFD0 U844 ( .I(n847), .Z(n846) );
  BUFFD0 U845 ( .I(n848), .Z(n847) );
  BUFFD0 U846 ( .I(n849), .Z(n848) );
  BUFFD0 U847 ( .I(n850), .Z(n849) );
  BUFFD0 U848 ( .I(n851), .Z(n850) );
  BUFFD0 U849 ( .I(n852), .Z(n851) );
  BUFFD0 U850 ( .I(n853), .Z(n852) );
  BUFFD0 U851 ( .I(n854), .Z(n853) );
  BUFFD0 U852 ( .I(n855), .Z(n854) );
  BUFFD0 U853 ( .I(n856), .Z(n855) );
  BUFFD0 U854 ( .I(n858), .Z(n856) );
  INVD0 U855 ( .I(n857), .ZN(n858) );
  CKNXD16 U856 ( .I(n806), .ZN(n857) );
  BUFFD0 U857 ( .I(n914), .Z(n859) );
  BUFFD0 U858 ( .I(n859), .Z(n860) );
  BUFFD0 U859 ( .I(n860), .Z(n861) );
  BUFFD0 U860 ( .I(n861), .Z(n862) );
  BUFFD0 U861 ( .I(n862), .Z(n863) );
  BUFFD0 U862 ( .I(n863), .Z(n864) );
  BUFFD0 U863 ( .I(n864), .Z(n865) );
  BUFFD0 U864 ( .I(n865), .Z(n866) );
  BUFFD0 U865 ( .I(n866), .Z(n867) );
  BUFFD0 U866 ( .I(n867), .Z(n868) );
  BUFFD0 U867 ( .I(n868), .Z(n869) );
  BUFFD0 U868 ( .I(n869), .Z(n870) );
  BUFFD0 U869 ( .I(n870), .Z(n871) );
  BUFFD0 U870 ( .I(n871), .Z(n872) );
  BUFFD0 U871 ( .I(n872), .Z(n873) );
  BUFFD0 U872 ( .I(n873), .Z(n874) );
  BUFFD0 U873 ( .I(n874), .Z(n875) );
  BUFFD0 U874 ( .I(n875), .Z(n876) );
  BUFFD0 U875 ( .I(n876), .Z(n877) );
  BUFFD0 U876 ( .I(n877), .Z(n878) );
  BUFFD0 U877 ( .I(n878), .Z(n879) );
  BUFFD0 U878 ( .I(n879), .Z(n880) );
  BUFFD0 U879 ( .I(n880), .Z(n881) );
  BUFFD0 U880 ( .I(n881), .Z(n882) );
  BUFFD0 U881 ( .I(n882), .Z(n883) );
  BUFFD0 U882 ( .I(n883), .Z(n884) );
  BUFFD0 U883 ( .I(n884), .Z(n885) );
  BUFFD0 U884 ( .I(n885), .Z(n886) );
  BUFFD0 U885 ( .I(n886), .Z(n887) );
  BUFFD0 U886 ( .I(n887), .Z(n888) );
  BUFFD0 U887 ( .I(n888), .Z(n889) );
  BUFFD0 U888 ( .I(n889), .Z(n890) );
  BUFFD0 U889 ( .I(n890), .Z(n891) );
  BUFFD0 U890 ( .I(n891), .Z(n892) );
  BUFFD0 U891 ( .I(n892), .Z(n893) );
  BUFFD0 U892 ( .I(n893), .Z(n894) );
  BUFFD0 U893 ( .I(n894), .Z(n895) );
  BUFFD0 U894 ( .I(n895), .Z(n896) );
  BUFFD0 U895 ( .I(n896), .Z(n897) );
  BUFFD0 U896 ( .I(n897), .Z(n898) );
  BUFFD0 U897 ( .I(n898), .Z(n899) );
  BUFFD0 U898 ( .I(n899), .Z(n900) );
  BUFFD0 U899 ( .I(n900), .Z(n901) );
  BUFFD0 U900 ( .I(n901), .Z(n902) );
  BUFFD0 U901 ( .I(n902), .Z(n903) );
  BUFFD0 U902 ( .I(n903), .Z(n904) );
  BUFFD0 U903 ( .I(n904), .Z(n905) );
  BUFFD0 U904 ( .I(n905), .Z(n906) );
  BUFFD0 U905 ( .I(n906), .Z(n907) );
  BUFFD0 U906 ( .I(n907), .Z(n908) );
  BUFFD0 U907 ( .I(n908), .Z(n909) );
  BUFFD0 U908 ( .I(n909), .Z(n910) );
  BUFFD0 U909 ( .I(n910), .Z(n911) );
  BUFFD0 U910 ( .I(n911), .Z(n912) );
  BUFFD0 U911 ( .I(n912), .Z(n913) );
  BUFFD0 U912 ( .I(n3730), .Z(n914) );
  CKBD0 U913 ( .CLK(n913), .C(n915) );
  CKBD0 U914 ( .CLK(n3729), .C(n916) );
  BUFFD0 U915 ( .I(n916), .Z(n917) );
  BUFFD0 U916 ( .I(n917), .Z(n918) );
  BUFFD0 U917 ( .I(n918), .Z(n919) );
  BUFFD0 U918 ( .I(n919), .Z(n920) );
  BUFFD0 U919 ( .I(n920), .Z(n921) );
  BUFFD0 U920 ( .I(n921), .Z(n922) );
  BUFFD0 U921 ( .I(n922), .Z(n923) );
  BUFFD0 U922 ( .I(n923), .Z(n924) );
  BUFFD0 U923 ( .I(n924), .Z(n925) );
  BUFFD0 U924 ( .I(n925), .Z(n926) );
  BUFFD0 U925 ( .I(n926), .Z(n927) );
  BUFFD0 U926 ( .I(n927), .Z(n928) );
  BUFFD0 U927 ( .I(n928), .Z(n929) );
  BUFFD0 U928 ( .I(n929), .Z(n930) );
  BUFFD0 U929 ( .I(n930), .Z(n931) );
  BUFFD0 U930 ( .I(n931), .Z(n932) );
  BUFFD0 U931 ( .I(n932), .Z(n933) );
  BUFFD0 U932 ( .I(n933), .Z(n934) );
  BUFFD0 U933 ( .I(n934), .Z(n935) );
  BUFFD0 U934 ( .I(n935), .Z(n936) );
  BUFFD0 U935 ( .I(n936), .Z(n937) );
  BUFFD0 U936 ( .I(n937), .Z(n938) );
  BUFFD0 U937 ( .I(n938), .Z(n939) );
  BUFFD0 U938 ( .I(n939), .Z(n940) );
  BUFFD0 U939 ( .I(n940), .Z(n941) );
  BUFFD0 U940 ( .I(n941), .Z(n942) );
  BUFFD0 U941 ( .I(n942), .Z(n943) );
  BUFFD0 U942 ( .I(n943), .Z(n944) );
  BUFFD0 U943 ( .I(n944), .Z(n945) );
  BUFFD0 U944 ( .I(n945), .Z(n946) );
  BUFFD0 U945 ( .I(n946), .Z(n947) );
  BUFFD0 U946 ( .I(n947), .Z(n948) );
  BUFFD0 U947 ( .I(n948), .Z(n949) );
  BUFFD0 U948 ( .I(n949), .Z(n950) );
  BUFFD0 U949 ( .I(n950), .Z(n951) );
  BUFFD0 U950 ( .I(n951), .Z(n952) );
  BUFFD0 U951 ( .I(n952), .Z(n953) );
  BUFFD0 U952 ( .I(n953), .Z(n954) );
  BUFFD0 U953 ( .I(n954), .Z(n955) );
  BUFFD0 U954 ( .I(n955), .Z(n956) );
  BUFFD0 U955 ( .I(n956), .Z(n957) );
  BUFFD0 U956 ( .I(n957), .Z(n958) );
  BUFFD0 U957 ( .I(n958), .Z(n959) );
  BUFFD0 U958 ( .I(n959), .Z(n960) );
  BUFFD0 U959 ( .I(n960), .Z(n961) );
  BUFFD0 U960 ( .I(n961), .Z(n962) );
  BUFFD0 U961 ( .I(n962), .Z(n963) );
  BUFFD0 U962 ( .I(n963), .Z(n964) );
  BUFFD0 U963 ( .I(n964), .Z(n965) );
  BUFFD0 U964 ( .I(n965), .Z(n966) );
  BUFFD0 U965 ( .I(n966), .Z(n967) );
  BUFFD0 U966 ( .I(n967), .Z(n968) );
  BUFFD0 U967 ( .I(n968), .Z(n969) );
  BUFFD0 U968 ( .I(n969), .Z(n970) );
  CKBD0 U969 ( .CLK(n970), .C(n971) );
  INVD10 U970 ( .I(n3728), .ZN(n972) );
  BUFFD0 U971 ( .I(n976), .Z(n974) );
  BUFFD0 U972 ( .I(n974), .Z(n975) );
  BUFFD0 U973 ( .I(n977), .Z(n976) );
  BUFFD0 U974 ( .I(n978), .Z(n977) );
  BUFFD0 U975 ( .I(n979), .Z(n978) );
  BUFFD0 U976 ( .I(n980), .Z(n979) );
  BUFFD0 U977 ( .I(n981), .Z(n980) );
  BUFFD0 U978 ( .I(n982), .Z(n981) );
  BUFFD0 U979 ( .I(n983), .Z(n982) );
  BUFFD0 U980 ( .I(n984), .Z(n983) );
  BUFFD0 U981 ( .I(n985), .Z(n984) );
  BUFFD0 U982 ( .I(n986), .Z(n985) );
  BUFFD0 U983 ( .I(n987), .Z(n986) );
  BUFFD0 U984 ( .I(n988), .Z(n987) );
  BUFFD0 U985 ( .I(n989), .Z(n988) );
  BUFFD0 U986 ( .I(n990), .Z(n989) );
  BUFFD0 U987 ( .I(n991), .Z(n990) );
  BUFFD0 U988 ( .I(n992), .Z(n991) );
  BUFFD0 U989 ( .I(n993), .Z(n992) );
  BUFFD0 U990 ( .I(n994), .Z(n993) );
  BUFFD0 U991 ( .I(n995), .Z(n994) );
  BUFFD0 U992 ( .I(n996), .Z(n995) );
  BUFFD0 U993 ( .I(n997), .Z(n996) );
  BUFFD0 U994 ( .I(n998), .Z(n997) );
  BUFFD0 U995 ( .I(n999), .Z(n998) );
  BUFFD0 U996 ( .I(n1000), .Z(n999) );
  BUFFD0 U997 ( .I(n1001), .Z(n1000) );
  BUFFD0 U998 ( .I(n1002), .Z(n1001) );
  BUFFD0 U999 ( .I(n1003), .Z(n1002) );
  BUFFD0 U1000 ( .I(n1004), .Z(n1003) );
  BUFFD0 U1001 ( .I(n1005), .Z(n1004) );
  BUFFD0 U1002 ( .I(n1006), .Z(n1005) );
  BUFFD0 U1003 ( .I(n1007), .Z(n1006) );
  BUFFD0 U1004 ( .I(n1008), .Z(n1007) );
  BUFFD0 U1005 ( .I(n1009), .Z(n1008) );
  BUFFD0 U1006 ( .I(n1010), .Z(n1009) );
  BUFFD0 U1007 ( .I(n1011), .Z(n1010) );
  BUFFD0 U1008 ( .I(n1012), .Z(n1011) );
  BUFFD0 U1009 ( .I(n1013), .Z(n1012) );
  BUFFD0 U1010 ( .I(n1014), .Z(n1013) );
  BUFFD0 U1011 ( .I(n1015), .Z(n1014) );
  BUFFD0 U1012 ( .I(n1016), .Z(n1015) );
  BUFFD0 U1013 ( .I(n1017), .Z(n1016) );
  BUFFD0 U1014 ( .I(n1018), .Z(n1017) );
  BUFFD0 U1015 ( .I(n1019), .Z(n1018) );
  BUFFD0 U1016 ( .I(n1020), .Z(n1019) );
  BUFFD0 U1017 ( .I(n1022), .Z(n1020) );
  INVD0 U1018 ( .I(n1021), .ZN(n1022) );
  CKNXD16 U1019 ( .I(n3727), .ZN(n1021) );
  INVD10 U1020 ( .I(n3726), .ZN(n1023) );
  BUFFD0 U1021 ( .I(n1029), .Z(n1025) );
  BUFFD0 U1022 ( .I(n3617), .Z(n1026) );
  BUFFD0 U1023 ( .I(n1026), .Z(n1027) );
  BUFFD0 U1024 ( .I(n1027), .Z(n1028) );
  BUFFD0 U1025 ( .I(n1030), .Z(n1029) );
  BUFFD0 U1026 ( .I(n1031), .Z(n1030) );
  BUFFD0 U1027 ( .I(n1032), .Z(n1031) );
  BUFFD0 U1028 ( .I(n1033), .Z(n1032) );
  BUFFD0 U1029 ( .I(n1034), .Z(n1033) );
  BUFFD0 U1030 ( .I(n1035), .Z(n1034) );
  BUFFD0 U1031 ( .I(n1036), .Z(n1035) );
  BUFFD0 U1032 ( .I(n1037), .Z(n1036) );
  BUFFD0 U1033 ( .I(n1038), .Z(n1037) );
  BUFFD0 U1034 ( .I(n1039), .Z(n1038) );
  BUFFD0 U1035 ( .I(n1040), .Z(n1039) );
  BUFFD0 U1036 ( .I(n1041), .Z(n1040) );
  BUFFD0 U1037 ( .I(n1042), .Z(n1041) );
  BUFFD0 U1038 ( .I(n1043), .Z(n1042) );
  BUFFD0 U1039 ( .I(n1044), .Z(n1043) );
  BUFFD0 U1040 ( .I(n1045), .Z(n1044) );
  BUFFD0 U1041 ( .I(n1046), .Z(n1045) );
  BUFFD0 U1042 ( .I(n1047), .Z(n1046) );
  BUFFD0 U1043 ( .I(n1048), .Z(n1047) );
  BUFFD0 U1044 ( .I(n1049), .Z(n1048) );
  BUFFD0 U1045 ( .I(n1050), .Z(n1049) );
  BUFFD0 U1046 ( .I(n1051), .Z(n1050) );
  BUFFD0 U1047 ( .I(n1052), .Z(n1051) );
  BUFFD0 U1048 ( .I(n1053), .Z(n1052) );
  BUFFD0 U1049 ( .I(n1054), .Z(n1053) );
  BUFFD0 U1050 ( .I(n1055), .Z(n1054) );
  BUFFD0 U1051 ( .I(n1056), .Z(n1055) );
  BUFFD0 U1052 ( .I(n1057), .Z(n1056) );
  BUFFD0 U1053 ( .I(n1058), .Z(n1057) );
  BUFFD0 U1054 ( .I(n1059), .Z(n1058) );
  BUFFD0 U1055 ( .I(n1060), .Z(n1059) );
  BUFFD0 U1056 ( .I(n1061), .Z(n1060) );
  BUFFD0 U1057 ( .I(n1062), .Z(n1061) );
  BUFFD0 U1058 ( .I(n1063), .Z(n1062) );
  BUFFD0 U1059 ( .I(n1064), .Z(n1063) );
  BUFFD0 U1060 ( .I(n1065), .Z(n1064) );
  BUFFD0 U1061 ( .I(n1066), .Z(n1065) );
  BUFFD0 U1062 ( .I(n1067), .Z(n1066) );
  BUFFD0 U1063 ( .I(n1068), .Z(n1067) );
  BUFFD0 U1064 ( .I(n1069), .Z(n1068) );
  BUFFD0 U1065 ( .I(n1070), .Z(n1069) );
  BUFFD0 U1066 ( .I(n1071), .Z(n1070) );
  BUFFD0 U1067 ( .I(n1072), .Z(n1071) );
  BUFFD0 U1068 ( .I(n1073), .Z(n1072) );
  BUFFD0 U1069 ( .I(n1074), .Z(n1073) );
  BUFFD0 U1070 ( .I(n1075), .Z(n1074) );
  BUFFD0 U1071 ( .I(n1076), .Z(n1075) );
  BUFFD0 U1072 ( .I(n1077), .Z(n1076) );
  BUFFD0 U1073 ( .I(n1078), .Z(n1077) );
  BUFFD0 U1074 ( .I(n1079), .Z(n1078) );
  BUFFD0 U1075 ( .I(n1080), .Z(n1079) );
  BUFFD0 U1076 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1077 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1078 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1079 ( .I(n1085), .Z(n1083) );
  BUFFD0 U1080 ( .I(n1087), .Z(n1084) );
  BUFFD0 U1081 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1082 ( .I(n1028), .Z(n1086) );
  BUFFD0 U1083 ( .I(Dreadyr), .Z(n1087) );
  OR2D0 U1084 ( .A1(n3815), .A2(n1084), .Z(n3617) );
  IND2D0 U1085 ( .A1(AddrW[2]), .B1(Write), .ZN(n66) );
  BUFFD0 U1086 ( .I(N87), .Z(n1088) );
  BUFFD0 U1087 ( .I(n1088), .Z(n1089) );
  BUFFD0 U1088 ( .I(n1089), .Z(n1090) );
  BUFFD0 U1089 ( .I(n1090), .Z(n1091) );
  BUFFD0 U1090 ( .I(n1091), .Z(n1092) );
  BUFFD0 U1091 ( .I(n1092), .Z(n1093) );
  BUFFD0 U1092 ( .I(n1093), .Z(n1094) );
  BUFFD0 U1093 ( .I(n1094), .Z(n1095) );
  BUFFD0 U1094 ( .I(n1095), .Z(n1096) );
  BUFFD0 U1095 ( .I(n1096), .Z(n1097) );
  BUFFD0 U1096 ( .I(n1097), .Z(n1098) );
  BUFFD0 U1097 ( .I(n1098), .Z(n1099) );
  BUFFD0 U1098 ( .I(n1099), .Z(n1100) );
  BUFFD0 U1099 ( .I(n1100), .Z(n1101) );
  BUFFD0 U1100 ( .I(n1101), .Z(n1102) );
  BUFFD0 U1101 ( .I(n1102), .Z(n1103) );
  BUFFD0 U1102 ( .I(n1103), .Z(n1104) );
  BUFFD0 U1103 ( .I(n1104), .Z(n1105) );
  BUFFD0 U1104 ( .I(n1105), .Z(n1106) );
  BUFFD0 U1105 ( .I(n1106), .Z(n1107) );
  BUFFD0 U1106 ( .I(n1107), .Z(n1108) );
  BUFFD0 U1107 ( .I(n1108), .Z(n1109) );
  BUFFD0 U1108 ( .I(n1109), .Z(n1110) );
  BUFFD0 U1109 ( .I(n1110), .Z(n1111) );
  BUFFD0 U1110 ( .I(n1111), .Z(n1112) );
  BUFFD0 U1111 ( .I(n1112), .Z(n1113) );
  BUFFD0 U1112 ( .I(n1113), .Z(n1114) );
  BUFFD0 U1113 ( .I(n1114), .Z(n1115) );
  BUFFD0 U1114 ( .I(n1115), .Z(n1116) );
  BUFFD0 U1115 ( .I(n1116), .Z(n1117) );
  BUFFD0 U1116 ( .I(n1117), .Z(n1118) );
  BUFFD0 U1117 ( .I(n1118), .Z(n1119) );
  BUFFD0 U1118 ( .I(n1119), .Z(n1120) );
  BUFFD0 U1119 ( .I(n1120), .Z(n1121) );
  BUFFD0 U1120 ( .I(n1121), .Z(n1122) );
  BUFFD0 U1121 ( .I(n1122), .Z(n1123) );
  BUFFD0 U1122 ( .I(n1123), .Z(n1124) );
  BUFFD0 U1123 ( .I(n1124), .Z(n1125) );
  BUFFD0 U1124 ( .I(n1125), .Z(n1126) );
  BUFFD0 U1125 ( .I(n1126), .Z(n1127) );
  BUFFD0 U1126 ( .I(n1127), .Z(n1128) );
  BUFFD0 U1127 ( .I(n1128), .Z(n1129) );
  BUFFD0 U1128 ( .I(n1129), .Z(n1130) );
  BUFFD0 U1129 ( .I(n1130), .Z(n1131) );
  BUFFD0 U1130 ( .I(n1131), .Z(n1132) );
  BUFFD0 U1131 ( .I(n1132), .Z(n1133) );
  BUFFD0 U1132 ( .I(n1133), .Z(n1134) );
  BUFFD0 U1133 ( .I(n1134), .Z(n1135) );
  BUFFD0 U1134 ( .I(n1135), .Z(n1136) );
  XOR3D0 U1135 ( .A1(n3740), .A2(n1264), .A3(n76), .Z(n75) );
  CKBD0 U1136 ( .CLK(DataI[22]), .C(n3743) );
  CKBD0 U1137 ( .CLK(DataI[17]), .C(n3738) );
  CKBD0 U1138 ( .CLK(DataI[15]), .C(n3737) );
  CKBD0 U1139 ( .CLK(DataI[10]), .C(n3734) );
  CKBD0 U1140 ( .CLK(DataI[14]), .C(n3736) );
  CKBD0 U1141 ( .CLK(DataI[11]), .C(n3735) );
  XOR3D0 U1142 ( .A1(n3726), .A2(n68), .A3(n69), .Z(n67) );
  CKBD0 U1143 ( .CLK(DataI[8]), .C(n3733) );
  CKBD0 U1144 ( .CLK(DataI[7]), .C(n3732) );
  CKBD0 U1145 ( .CLK(DataI[3]), .C(n3729) );
  CKBD0 U1146 ( .CLK(n1136), .C(n1137) );
  XOR3D0 U1147 ( .A1(n3728), .A2(n3727), .A3(n67), .Z(N87) );
  CKBD0 U1148 ( .CLK(DataI[4]), .C(n3730) );
  CKBD0 U1149 ( .CLK(DataI[1]), .C(n3727) );
  BUFFD0 U1150 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1151 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1152 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1153 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1154 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1155 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1156 ( .I(n1147), .Z(n1145) );
  INVD0 U1157 ( .I(n1146), .ZN(n1147) );
  CKNXD16 U1158 ( .I(n3751), .ZN(n1146) );
  CKBD0 U1159 ( .CLK(DataI[31]), .C(n3751) );
  BUFFD0 U1160 ( .I(n1159), .Z(n1148) );
  BUFFD0 U1161 ( .I(n1148), .Z(n1149) );
  BUFFD0 U1162 ( .I(n1149), .Z(n1150) );
  BUFFD0 U1163 ( .I(n1150), .Z(n1151) );
  BUFFD0 U1164 ( .I(n1151), .Z(n1152) );
  BUFFD0 U1165 ( .I(n1152), .Z(n1153) );
  BUFFD0 U1166 ( .I(n1153), .Z(n1154) );
  BUFFD0 U1167 ( .I(n1154), .Z(n1155) );
  BUFFD0 U1168 ( .I(n1155), .Z(n1156) );
  BUFFD0 U1169 ( .I(n1156), .Z(n1157) );
  BUFFD0 U1170 ( .I(n1157), .Z(n1158) );
  BUFFD0 U1171 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1172 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1173 ( .I(n3750), .Z(n1161) );
  CKBD0 U1174 ( .CLK(n1158), .C(n1162) );
  CKBD0 U1175 ( .CLK(DataI[30]), .C(n3750) );
  BUFFD0 U1176 ( .I(n1174), .Z(n1163) );
  BUFFD0 U1177 ( .I(n1163), .Z(n1164) );
  BUFFD0 U1178 ( .I(n1164), .Z(n1165) );
  BUFFD0 U1179 ( .I(n1165), .Z(n1166) );
  BUFFD0 U1180 ( .I(n1166), .Z(n1167) );
  BUFFD0 U1181 ( .I(n1167), .Z(n1168) );
  BUFFD0 U1182 ( .I(n1168), .Z(n1169) );
  BUFFD0 U1183 ( .I(n1169), .Z(n1170) );
  BUFFD0 U1184 ( .I(n1170), .Z(n1171) );
  BUFFD0 U1185 ( .I(n1171), .Z(n1172) );
  BUFFD0 U1186 ( .I(n1172), .Z(n1173) );
  BUFFD0 U1187 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1188 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1189 ( .I(n3749), .Z(n1176) );
  CKBD0 U1190 ( .CLK(n1173), .C(n1177) );
  CKBD0 U1191 ( .CLK(DataI[29]), .C(n3749) );
  BUFFD0 U1192 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1193 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1194 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1195 ( .I(n1183), .Z(n1182) );
  BUFFD0 U1196 ( .I(n1184), .Z(n1183) );
  BUFFD0 U1197 ( .I(n1185), .Z(n1184) );
  BUFFD0 U1198 ( .I(n1187), .Z(n1185) );
  INVD0 U1199 ( .I(n1186), .ZN(n1187) );
  CKNXD16 U1200 ( .I(n3748), .ZN(n1186) );
  CKBD0 U1201 ( .CLK(DataI[28]), .C(n3748) );
  BUFFD0 U1202 ( .I(n1190), .Z(n1189) );
  BUFFD0 U1203 ( .I(n1191), .Z(n1190) );
  BUFFD0 U1204 ( .I(n1192), .Z(n1191) );
  BUFFD0 U1205 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1206 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1207 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1208 ( .I(n1197), .Z(n1195) );
  INVD0 U1209 ( .I(n1196), .ZN(n1197) );
  CKNXD16 U1210 ( .I(n3747), .ZN(n1196) );
  CKBD0 U1211 ( .CLK(DataI[27]), .C(n3747) );
  BUFFD0 U1212 ( .I(n1208), .Z(n1198) );
  BUFFD0 U1213 ( .I(n1198), .Z(n1199) );
  BUFFD0 U1214 ( .I(n1199), .Z(n1200) );
  BUFFD0 U1215 ( .I(n1200), .Z(n1201) );
  BUFFD0 U1216 ( .I(n1201), .Z(n1202) );
  BUFFD0 U1217 ( .I(n1202), .Z(n1203) );
  BUFFD0 U1218 ( .I(n1203), .Z(n1204) );
  BUFFD0 U1219 ( .I(n1204), .Z(n1205) );
  BUFFD0 U1220 ( .I(n1205), .Z(n1206) );
  BUFFD0 U1221 ( .I(n1206), .Z(n1207) );
  BUFFD0 U1222 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1223 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1224 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1225 ( .I(n3746), .Z(n1211) );
  CKBD0 U1226 ( .CLK(n1207), .C(n1212) );
  CKBD0 U1227 ( .CLK(DataI[26]), .C(n3746) );
  BUFFD0 U1228 ( .I(n1223), .Z(n1213) );
  BUFFD0 U1229 ( .I(n1213), .Z(n1214) );
  BUFFD0 U1230 ( .I(n1214), .Z(n1215) );
  BUFFD0 U1231 ( .I(n1215), .Z(n1216) );
  BUFFD0 U1232 ( .I(n1216), .Z(n1217) );
  BUFFD0 U1233 ( .I(n1217), .Z(n1218) );
  BUFFD0 U1234 ( .I(n1218), .Z(n1219) );
  BUFFD0 U1235 ( .I(n1219), .Z(n1220) );
  BUFFD0 U1236 ( .I(n1220), .Z(n1221) );
  BUFFD0 U1237 ( .I(n1221), .Z(n1222) );
  BUFFD0 U1238 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1239 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1240 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1241 ( .I(n3745), .Z(n1226) );
  CKBD0 U1242 ( .CLK(n1222), .C(n1227) );
  CKBD0 U1243 ( .CLK(DataI[25]), .C(n3745) );
  CKBD0 U1244 ( .CLK(n3744), .C(n1228) );
  CKBXD2 U1245 ( .I(DataI[24]), .Z(n3744) );
  BUFFD0 U1246 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1247 ( .I(n1233), .Z(n1231) );
  INVD0 U1248 ( .I(n1232), .ZN(n1233) );
  CKNXD16 U1249 ( .I(n1228), .ZN(n1232) );
  BUFFD0 U1250 ( .I(n3742), .Z(n1234) );
  BUFFD0 U1251 ( .I(n1234), .Z(n1235) );
  BUFFD0 U1252 ( .I(n1235), .Z(n1236) );
  BUFFD0 U1253 ( .I(n1236), .Z(n1237) );
  BUFFD0 U1254 ( .I(n1237), .Z(n1238) );
  BUFFD0 U1255 ( .I(n1238), .Z(n1239) );
  BUFFD0 U1256 ( .I(n1239), .Z(n1240) );
  BUFFD0 U1257 ( .I(n1240), .Z(n1241) );
  BUFFD0 U1258 ( .I(n1241), .Z(n1242) );
  CKBD0 U1259 ( .CLK(n1242), .C(n1243) );
  CKBD0 U1260 ( .CLK(DataI[21]), .C(n3742) );
  CKBD0 U1261 ( .CLK(n3741), .C(n1244) );
  BUFFD10 U1262 ( .I(DataI[20]), .Z(n3741) );
  BUFFD0 U1263 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1264 ( .I(n1249), .Z(n1247) );
  INVD0 U1265 ( .I(n1248), .ZN(n1249) );
  CKNXD16 U1266 ( .I(n1244), .ZN(n1248) );
  INVD16 U1267 ( .I(n3740), .ZN(n1250) );
  INVD1 U1268 ( .I(n1250), .ZN(n1251) );
  BUFFD0 U1269 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1270 ( .I(n1256), .Z(n1254) );
  INVD0 U1271 ( .I(n1255), .ZN(n1256) );
  CKNXD16 U1272 ( .I(n1251), .ZN(n1255) );
  CKBD0 U1273 ( .CLK(DataI[19]), .C(n3740) );
  BUFFD0 U1274 ( .I(n1264), .Z(n1257) );
  BUFFD0 U1275 ( .I(n1257), .Z(n1258) );
  BUFFD0 U1276 ( .I(n1258), .Z(n1259) );
  BUFFD0 U1277 ( .I(n1259), .Z(n1260) );
  BUFFD0 U1278 ( .I(n1260), .Z(n1261) );
  BUFFD0 U1279 ( .I(n1261), .Z(n1262) );
  BUFFD0 U1280 ( .I(n1262), .Z(n1263) );
  BUFFD0 U1281 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1282 ( .I(n3739), .Z(n1265) );
  CKBD0 U1283 ( .CLK(n1263), .C(n1266) );
  CKBD0 U1284 ( .CLK(DataI[18]), .C(n3739) );
  BUFFD0 U1285 ( .I(n92), .Z(n1267) );
  BUFFD0 U1286 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1287 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1288 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1289 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1290 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1291 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1292 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1293 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1294 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1295 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1296 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1297 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1298 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1299 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1300 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1301 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1302 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1303 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1304 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1305 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1306 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1307 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1308 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1309 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1310 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1311 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1312 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1313 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1314 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1315 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1316 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1317 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1318 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1319 ( .I(n1302), .Z(n1301) );
  BUFFD0 U1320 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1321 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1322 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1323 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1324 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1325 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1326 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1327 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1328 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1329 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1330 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1331 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1332 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1333 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1334 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1335 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1336 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1337 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1338 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1339 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1340 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1341 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1342 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1343 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1344 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1345 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1346 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1347 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1348 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1349 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1350 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1351 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1352 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1353 ( .I(n1336), .Z(n1335) );
  BUFFD0 U1354 ( .I(n1337), .Z(n1336) );
  BUFFD0 U1355 ( .I(N53), .Z(n1337) );
  BUFFD0 U1356 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1357 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1358 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1359 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1360 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1361 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1362 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1363 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1364 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1365 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1366 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1367 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1368 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1369 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1370 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1371 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1372 ( .I(n1355), .Z(n1354) );
  BUFFD0 U1373 ( .I(n1356), .Z(n1355) );
  BUFFD0 U1374 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1375 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1376 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1377 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1378 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1379 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1380 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1381 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1382 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1383 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1384 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1385 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1386 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1387 ( .I(n1370), .Z(n1369) );
  BUFFD0 U1388 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1389 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1390 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1391 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1392 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1393 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1394 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1395 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1396 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1397 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1398 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1399 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1400 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1401 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1402 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1403 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1404 ( .I(n1387), .Z(n1386) );
  BUFFD0 U1405 ( .I(n1388), .Z(n1387) );
  BUFFD0 U1406 ( .I(n1389), .Z(n1388) );
  BUFFD0 U1407 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1408 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1409 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1410 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1411 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1412 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1413 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1414 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1415 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1416 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1417 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1418 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1419 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1420 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1421 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1422 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1423 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1424 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1425 ( .I(N54), .Z(n1407) );
  BUFFD0 U1426 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1427 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1428 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1429 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1430 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1431 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1432 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1433 ( .I(n1416), .Z(n1415) );
  BUFFD0 U1434 ( .I(n1417), .Z(n1416) );
  BUFFD0 U1435 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1436 ( .I(n1419), .Z(n1418) );
  BUFFD0 U1437 ( .I(n1420), .Z(n1419) );
  BUFFD0 U1438 ( .I(n1421), .Z(n1420) );
  BUFFD0 U1439 ( .I(n1422), .Z(n1421) );
  BUFFD0 U1440 ( .I(n1423), .Z(n1422) );
  BUFFD0 U1441 ( .I(n1424), .Z(n1423) );
  BUFFD0 U1442 ( .I(n1425), .Z(n1424) );
  BUFFD0 U1443 ( .I(n1426), .Z(n1425) );
  BUFFD0 U1444 ( .I(n1427), .Z(n1426) );
  BUFFD0 U1445 ( .I(n1428), .Z(n1427) );
  BUFFD0 U1446 ( .I(n1429), .Z(n1428) );
  BUFFD0 U1447 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1448 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1449 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1450 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1451 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1452 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1453 ( .I(n1436), .Z(n1435) );
  BUFFD0 U1454 ( .I(n1437), .Z(n1436) );
  BUFFD0 U1455 ( .I(n1438), .Z(n1437) );
  BUFFD0 U1456 ( .I(n1439), .Z(n1438) );
  BUFFD0 U1457 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1458 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1459 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1460 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1461 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1462 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1463 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1464 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1465 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1466 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1467 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1468 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1469 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1470 ( .I(n1453), .Z(n1452) );
  BUFFD0 U1471 ( .I(n1454), .Z(n1453) );
  BUFFD0 U1472 ( .I(n1455), .Z(n1454) );
  BUFFD0 U1473 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1474 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1475 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1476 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1477 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1478 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1479 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1480 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1481 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1482 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1483 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1484 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1485 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1486 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1487 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1488 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1489 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1490 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1491 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1492 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1493 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1494 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1495 ( .I(N55), .Z(n1477) );
  BUFFD0 U1496 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1497 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1498 ( .I(n1481), .Z(n1480) );
  BUFFD0 U1499 ( .I(n1482), .Z(n1481) );
  BUFFD0 U1500 ( .I(n1483), .Z(n1482) );
  BUFFD0 U1501 ( .I(n1484), .Z(n1483) );
  BUFFD0 U1502 ( .I(n1485), .Z(n1484) );
  BUFFD0 U1503 ( .I(n1486), .Z(n1485) );
  BUFFD0 U1504 ( .I(n1487), .Z(n1486) );
  BUFFD0 U1505 ( .I(n1488), .Z(n1487) );
  BUFFD0 U1506 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1507 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1508 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1509 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1510 ( .I(n1493), .Z(n1492) );
  BUFFD0 U1511 ( .I(n1494), .Z(n1493) );
  BUFFD0 U1512 ( .I(n1495), .Z(n1494) );
  BUFFD0 U1513 ( .I(n1496), .Z(n1495) );
  BUFFD0 U1514 ( .I(n1497), .Z(n1496) );
  BUFFD0 U1515 ( .I(n1498), .Z(n1497) );
  BUFFD0 U1516 ( .I(n1499), .Z(n1498) );
  BUFFD0 U1517 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1518 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1519 ( .I(n1502), .Z(n1501) );
  BUFFD0 U1520 ( .I(n1503), .Z(n1502) );
  BUFFD0 U1521 ( .I(n1504), .Z(n1503) );
  BUFFD0 U1522 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1523 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1524 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1525 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1526 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1527 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1528 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1529 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1530 ( .I(n1513), .Z(n1512) );
  BUFFD0 U1531 ( .I(n1514), .Z(n1513) );
  BUFFD0 U1532 ( .I(n1515), .Z(n1514) );
  BUFFD0 U1533 ( .I(n1516), .Z(n1515) );
  BUFFD0 U1534 ( .I(n1517), .Z(n1516) );
  BUFFD0 U1535 ( .I(n1518), .Z(n1517) );
  BUFFD0 U1536 ( .I(n1519), .Z(n1518) );
  BUFFD0 U1537 ( .I(n1520), .Z(n1519) );
  BUFFD0 U1538 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1539 ( .I(n1522), .Z(n1521) );
  BUFFD0 U1540 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1541 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1542 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1543 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1544 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1545 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1546 ( .I(n1529), .Z(n1528) );
  BUFFD0 U1547 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1548 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1549 ( .I(n1532), .Z(n1531) );
  BUFFD0 U1550 ( .I(n1533), .Z(n1532) );
  BUFFD0 U1551 ( .I(n1534), .Z(n1533) );
  BUFFD0 U1552 ( .I(n1535), .Z(n1534) );
  BUFFD0 U1553 ( .I(n1536), .Z(n1535) );
  BUFFD0 U1554 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1555 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1556 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1557 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1558 ( .I(n1541), .Z(n1540) );
  BUFFD0 U1559 ( .I(n1542), .Z(n1541) );
  BUFFD0 U1560 ( .I(n1543), .Z(n1542) );
  BUFFD0 U1561 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1562 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1563 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1564 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1565 ( .I(N56), .Z(n1547) );
  BUFFD0 U1566 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1567 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1568 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1569 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1570 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1571 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1572 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1573 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1574 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1575 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1576 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1577 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1578 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1579 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1580 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1581 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1582 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1583 ( .I(n1566), .Z(n1565) );
  BUFFD0 U1584 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1585 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1586 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1587 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1588 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1589 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1590 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1591 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1592 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1593 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1594 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1595 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1596 ( .I(n1579), .Z(n1578) );
  BUFFD0 U1597 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1598 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1599 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1600 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1601 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1602 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1603 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1604 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1605 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1606 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1607 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1608 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1609 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1610 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1611 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1612 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1613 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1614 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1615 ( .I(n1598), .Z(n1597) );
  BUFFD0 U1616 ( .I(n1599), .Z(n1598) );
  BUFFD0 U1617 ( .I(n1600), .Z(n1599) );
  BUFFD0 U1618 ( .I(n1601), .Z(n1600) );
  BUFFD0 U1619 ( .I(n1602), .Z(n1601) );
  BUFFD0 U1620 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1621 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1622 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1623 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1624 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1625 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1626 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1627 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1628 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1629 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1630 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1631 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1632 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1633 ( .I(n1616), .Z(n1615) );
  BUFFD0 U1634 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1635 ( .I(N57), .Z(n1617) );
  BUFFD0 U1636 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1637 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1638 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1639 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1640 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1641 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1642 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1643 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1644 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1645 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1646 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1647 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1648 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1649 ( .I(n1632), .Z(n1631) );
  BUFFD0 U1650 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1651 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1652 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1653 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1654 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1655 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1656 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1657 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1658 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1659 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1660 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1661 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1662 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1663 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1664 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1665 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1666 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1667 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1668 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1669 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1670 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1671 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1672 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1673 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1674 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1675 ( .I(n1658), .Z(n1657) );
  BUFFD0 U1676 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1677 ( .I(n1660), .Z(n1659) );
  BUFFD0 U1678 ( .I(n1661), .Z(n1660) );
  BUFFD0 U1679 ( .I(n1662), .Z(n1661) );
  BUFFD0 U1680 ( .I(n1663), .Z(n1662) );
  BUFFD0 U1681 ( .I(n1664), .Z(n1663) );
  BUFFD0 U1682 ( .I(n1665), .Z(n1664) );
  BUFFD0 U1683 ( .I(n1666), .Z(n1665) );
  BUFFD0 U1684 ( .I(n1667), .Z(n1666) );
  BUFFD0 U1685 ( .I(n1668), .Z(n1667) );
  BUFFD0 U1686 ( .I(n1669), .Z(n1668) );
  BUFFD0 U1687 ( .I(n1670), .Z(n1669) );
  BUFFD0 U1688 ( .I(n1671), .Z(n1670) );
  BUFFD0 U1689 ( .I(n1672), .Z(n1671) );
  BUFFD0 U1690 ( .I(n1673), .Z(n1672) );
  BUFFD0 U1691 ( .I(n1674), .Z(n1673) );
  BUFFD0 U1692 ( .I(n1675), .Z(n1674) );
  BUFFD0 U1693 ( .I(n1676), .Z(n1675) );
  BUFFD0 U1694 ( .I(n1677), .Z(n1676) );
  BUFFD0 U1695 ( .I(n1678), .Z(n1677) );
  BUFFD0 U1696 ( .I(n1679), .Z(n1678) );
  BUFFD0 U1697 ( .I(n1680), .Z(n1679) );
  BUFFD0 U1698 ( .I(n1681), .Z(n1680) );
  BUFFD0 U1699 ( .I(n1682), .Z(n1681) );
  BUFFD0 U1700 ( .I(n1683), .Z(n1682) );
  BUFFD0 U1701 ( .I(n1684), .Z(n1683) );
  BUFFD0 U1702 ( .I(n1685), .Z(n1684) );
  BUFFD0 U1703 ( .I(n1686), .Z(n1685) );
  BUFFD0 U1704 ( .I(n1687), .Z(n1686) );
  BUFFD0 U1705 ( .I(N58), .Z(n1687) );
  BUFFD0 U1706 ( .I(n1689), .Z(n1688) );
  BUFFD0 U1707 ( .I(n1690), .Z(n1689) );
  BUFFD0 U1708 ( .I(n1691), .Z(n1690) );
  BUFFD0 U1709 ( .I(n1692), .Z(n1691) );
  BUFFD0 U1710 ( .I(n1693), .Z(n1692) );
  BUFFD0 U1711 ( .I(n1694), .Z(n1693) );
  BUFFD0 U1712 ( .I(n1695), .Z(n1694) );
  BUFFD0 U1713 ( .I(n1696), .Z(n1695) );
  BUFFD0 U1714 ( .I(n1697), .Z(n1696) );
  BUFFD0 U1715 ( .I(n1698), .Z(n1697) );
  BUFFD0 U1716 ( .I(n1699), .Z(n1698) );
  BUFFD0 U1717 ( .I(n1700), .Z(n1699) );
  BUFFD0 U1718 ( .I(n1701), .Z(n1700) );
  BUFFD0 U1719 ( .I(n1702), .Z(n1701) );
  BUFFD0 U1720 ( .I(n1703), .Z(n1702) );
  BUFFD0 U1721 ( .I(n1704), .Z(n1703) );
  BUFFD0 U1722 ( .I(n1705), .Z(n1704) );
  BUFFD0 U1723 ( .I(n1706), .Z(n1705) );
  BUFFD0 U1724 ( .I(n1707), .Z(n1706) );
  BUFFD0 U1725 ( .I(n1708), .Z(n1707) );
  BUFFD0 U1726 ( .I(n1709), .Z(n1708) );
  BUFFD0 U1727 ( .I(n1710), .Z(n1709) );
  BUFFD0 U1728 ( .I(n1711), .Z(n1710) );
  BUFFD0 U1729 ( .I(n1712), .Z(n1711) );
  BUFFD0 U1730 ( .I(n1713), .Z(n1712) );
  BUFFD0 U1731 ( .I(n1714), .Z(n1713) );
  BUFFD0 U1732 ( .I(n1715), .Z(n1714) );
  BUFFD0 U1733 ( .I(n1716), .Z(n1715) );
  BUFFD0 U1734 ( .I(n1717), .Z(n1716) );
  BUFFD0 U1735 ( .I(n1718), .Z(n1717) );
  BUFFD0 U1736 ( .I(n1719), .Z(n1718) );
  BUFFD0 U1737 ( .I(n1720), .Z(n1719) );
  BUFFD0 U1738 ( .I(n1721), .Z(n1720) );
  BUFFD0 U1739 ( .I(n1722), .Z(n1721) );
  BUFFD0 U1740 ( .I(n1723), .Z(n1722) );
  BUFFD0 U1741 ( .I(n1724), .Z(n1723) );
  BUFFD0 U1742 ( .I(n1725), .Z(n1724) );
  BUFFD0 U1743 ( .I(n1726), .Z(n1725) );
  BUFFD0 U1744 ( .I(n1727), .Z(n1726) );
  BUFFD0 U1745 ( .I(n1728), .Z(n1727) );
  BUFFD0 U1746 ( .I(n1729), .Z(n1728) );
  BUFFD0 U1747 ( .I(n1730), .Z(n1729) );
  BUFFD0 U1748 ( .I(n1731), .Z(n1730) );
  BUFFD0 U1749 ( .I(n1732), .Z(n1731) );
  BUFFD0 U1750 ( .I(n1733), .Z(n1732) );
  BUFFD0 U1751 ( .I(n1734), .Z(n1733) );
  BUFFD0 U1752 ( .I(n1735), .Z(n1734) );
  BUFFD0 U1753 ( .I(n1736), .Z(n1735) );
  BUFFD0 U1754 ( .I(n1737), .Z(n1736) );
  BUFFD0 U1755 ( .I(n1738), .Z(n1737) );
  BUFFD0 U1756 ( .I(n1739), .Z(n1738) );
  BUFFD0 U1757 ( .I(n1740), .Z(n1739) );
  BUFFD0 U1758 ( .I(n1741), .Z(n1740) );
  BUFFD0 U1759 ( .I(n1742), .Z(n1741) );
  BUFFD0 U1760 ( .I(n1743), .Z(n1742) );
  BUFFD0 U1761 ( .I(n1744), .Z(n1743) );
  BUFFD0 U1762 ( .I(n1745), .Z(n1744) );
  BUFFD0 U1763 ( .I(n1746), .Z(n1745) );
  BUFFD0 U1764 ( .I(n1747), .Z(n1746) );
  BUFFD0 U1765 ( .I(n1748), .Z(n1747) );
  BUFFD0 U1766 ( .I(n1749), .Z(n1748) );
  BUFFD0 U1767 ( .I(n1750), .Z(n1749) );
  BUFFD0 U1768 ( .I(n1751), .Z(n1750) );
  BUFFD0 U1769 ( .I(n1752), .Z(n1751) );
  BUFFD0 U1770 ( .I(n1753), .Z(n1752) );
  BUFFD0 U1771 ( .I(n1754), .Z(n1753) );
  BUFFD0 U1772 ( .I(n1755), .Z(n1754) );
  BUFFD0 U1773 ( .I(n1756), .Z(n1755) );
  BUFFD0 U1774 ( .I(n1757), .Z(n1756) );
  BUFFD0 U1775 ( .I(N59), .Z(n1757) );
  BUFFD0 U1776 ( .I(n1759), .Z(n1758) );
  BUFFD0 U1777 ( .I(n1760), .Z(n1759) );
  BUFFD0 U1778 ( .I(n1761), .Z(n1760) );
  BUFFD0 U1779 ( .I(n1762), .Z(n1761) );
  BUFFD0 U1780 ( .I(n1763), .Z(n1762) );
  BUFFD0 U1781 ( .I(n1764), .Z(n1763) );
  BUFFD0 U1782 ( .I(n1765), .Z(n1764) );
  BUFFD0 U1783 ( .I(n1766), .Z(n1765) );
  BUFFD0 U1784 ( .I(n1767), .Z(n1766) );
  BUFFD0 U1785 ( .I(n1768), .Z(n1767) );
  BUFFD0 U1786 ( .I(n1769), .Z(n1768) );
  BUFFD0 U1787 ( .I(n1770), .Z(n1769) );
  BUFFD0 U1788 ( .I(n1771), .Z(n1770) );
  BUFFD0 U1789 ( .I(n1772), .Z(n1771) );
  BUFFD0 U1790 ( .I(n1773), .Z(n1772) );
  BUFFD0 U1791 ( .I(n1774), .Z(n1773) );
  BUFFD0 U1792 ( .I(n1775), .Z(n1774) );
  BUFFD0 U1793 ( .I(n1776), .Z(n1775) );
  BUFFD0 U1794 ( .I(n1777), .Z(n1776) );
  BUFFD0 U1795 ( .I(n1778), .Z(n1777) );
  BUFFD0 U1796 ( .I(n1779), .Z(n1778) );
  BUFFD0 U1797 ( .I(n1780), .Z(n1779) );
  BUFFD0 U1798 ( .I(n1781), .Z(n1780) );
  BUFFD0 U1799 ( .I(n1782), .Z(n1781) );
  BUFFD0 U1800 ( .I(n1783), .Z(n1782) );
  BUFFD0 U1801 ( .I(n1784), .Z(n1783) );
  BUFFD0 U1802 ( .I(n1785), .Z(n1784) );
  BUFFD0 U1803 ( .I(n1786), .Z(n1785) );
  BUFFD0 U1804 ( .I(n1787), .Z(n1786) );
  BUFFD0 U1805 ( .I(n1788), .Z(n1787) );
  BUFFD0 U1806 ( .I(n1789), .Z(n1788) );
  BUFFD0 U1807 ( .I(n1790), .Z(n1789) );
  BUFFD0 U1808 ( .I(n1791), .Z(n1790) );
  BUFFD0 U1809 ( .I(n1792), .Z(n1791) );
  BUFFD0 U1810 ( .I(n1793), .Z(n1792) );
  BUFFD0 U1811 ( .I(n1794), .Z(n1793) );
  BUFFD0 U1812 ( .I(n1795), .Z(n1794) );
  BUFFD0 U1813 ( .I(n1796), .Z(n1795) );
  BUFFD0 U1814 ( .I(n1797), .Z(n1796) );
  BUFFD0 U1815 ( .I(n1798), .Z(n1797) );
  BUFFD0 U1816 ( .I(n1799), .Z(n1798) );
  BUFFD0 U1817 ( .I(n1800), .Z(n1799) );
  BUFFD0 U1818 ( .I(n1801), .Z(n1800) );
  BUFFD0 U1819 ( .I(n1802), .Z(n1801) );
  BUFFD0 U1820 ( .I(n1803), .Z(n1802) );
  BUFFD0 U1821 ( .I(n1804), .Z(n1803) );
  BUFFD0 U1822 ( .I(n1805), .Z(n1804) );
  BUFFD0 U1823 ( .I(n1806), .Z(n1805) );
  BUFFD0 U1824 ( .I(n1807), .Z(n1806) );
  BUFFD0 U1825 ( .I(n1808), .Z(n1807) );
  BUFFD0 U1826 ( .I(n1809), .Z(n1808) );
  BUFFD0 U1827 ( .I(n1810), .Z(n1809) );
  BUFFD0 U1828 ( .I(n1811), .Z(n1810) );
  BUFFD0 U1829 ( .I(n1812), .Z(n1811) );
  BUFFD0 U1830 ( .I(n1813), .Z(n1812) );
  BUFFD0 U1831 ( .I(n1814), .Z(n1813) );
  BUFFD0 U1832 ( .I(n1815), .Z(n1814) );
  BUFFD0 U1833 ( .I(n1816), .Z(n1815) );
  BUFFD0 U1834 ( .I(n1817), .Z(n1816) );
  BUFFD0 U1835 ( .I(n1818), .Z(n1817) );
  BUFFD0 U1836 ( .I(n1819), .Z(n1818) );
  BUFFD0 U1837 ( .I(n1820), .Z(n1819) );
  BUFFD0 U1838 ( .I(n1821), .Z(n1820) );
  BUFFD0 U1839 ( .I(n1822), .Z(n1821) );
  BUFFD0 U1840 ( .I(n1823), .Z(n1822) );
  BUFFD0 U1841 ( .I(n1824), .Z(n1823) );
  BUFFD0 U1842 ( .I(n1825), .Z(n1824) );
  BUFFD0 U1843 ( .I(n1826), .Z(n1825) );
  BUFFD0 U1844 ( .I(n1827), .Z(n1826) );
  BUFFD0 U1845 ( .I(N60), .Z(n1827) );
  BUFFD0 U1846 ( .I(n1829), .Z(n1828) );
  BUFFD0 U1847 ( .I(n1830), .Z(n1829) );
  BUFFD0 U1848 ( .I(n1831), .Z(n1830) );
  BUFFD0 U1849 ( .I(n1832), .Z(n1831) );
  BUFFD0 U1850 ( .I(n1833), .Z(n1832) );
  BUFFD0 U1851 ( .I(n1834), .Z(n1833) );
  BUFFD0 U1852 ( .I(n1835), .Z(n1834) );
  BUFFD0 U1853 ( .I(n1836), .Z(n1835) );
  BUFFD0 U1854 ( .I(n1837), .Z(n1836) );
  BUFFD0 U1855 ( .I(n1838), .Z(n1837) );
  BUFFD0 U1856 ( .I(n1839), .Z(n1838) );
  BUFFD0 U1857 ( .I(n1840), .Z(n1839) );
  BUFFD0 U1858 ( .I(n1841), .Z(n1840) );
  BUFFD0 U1859 ( .I(n1842), .Z(n1841) );
  BUFFD0 U1860 ( .I(n1843), .Z(n1842) );
  BUFFD0 U1861 ( .I(n1844), .Z(n1843) );
  BUFFD0 U1862 ( .I(n1845), .Z(n1844) );
  BUFFD0 U1863 ( .I(n1846), .Z(n1845) );
  BUFFD0 U1864 ( .I(n1847), .Z(n1846) );
  BUFFD0 U1865 ( .I(n1848), .Z(n1847) );
  BUFFD0 U1866 ( .I(n1849), .Z(n1848) );
  BUFFD0 U1867 ( .I(n1850), .Z(n1849) );
  BUFFD0 U1868 ( .I(n1851), .Z(n1850) );
  BUFFD0 U1869 ( .I(n1852), .Z(n1851) );
  BUFFD0 U1870 ( .I(n1853), .Z(n1852) );
  BUFFD0 U1871 ( .I(n1854), .Z(n1853) );
  BUFFD0 U1872 ( .I(n1855), .Z(n1854) );
  BUFFD0 U1873 ( .I(n1856), .Z(n1855) );
  BUFFD0 U1874 ( .I(n1857), .Z(n1856) );
  BUFFD0 U1875 ( .I(n1858), .Z(n1857) );
  BUFFD0 U1876 ( .I(n1859), .Z(n1858) );
  BUFFD0 U1877 ( .I(n1860), .Z(n1859) );
  BUFFD0 U1878 ( .I(n1861), .Z(n1860) );
  BUFFD0 U1879 ( .I(n1862), .Z(n1861) );
  BUFFD0 U1880 ( .I(n1863), .Z(n1862) );
  BUFFD0 U1881 ( .I(n1864), .Z(n1863) );
  BUFFD0 U1882 ( .I(n1865), .Z(n1864) );
  BUFFD0 U1883 ( .I(n1866), .Z(n1865) );
  BUFFD0 U1884 ( .I(n1867), .Z(n1866) );
  BUFFD0 U1885 ( .I(n1868), .Z(n1867) );
  BUFFD0 U1886 ( .I(n1869), .Z(n1868) );
  BUFFD0 U1887 ( .I(n1870), .Z(n1869) );
  BUFFD0 U1888 ( .I(n1871), .Z(n1870) );
  BUFFD0 U1889 ( .I(n1872), .Z(n1871) );
  BUFFD0 U1890 ( .I(n1873), .Z(n1872) );
  BUFFD0 U1891 ( .I(n1874), .Z(n1873) );
  BUFFD0 U1892 ( .I(n1875), .Z(n1874) );
  BUFFD0 U1893 ( .I(n1876), .Z(n1875) );
  BUFFD0 U1894 ( .I(n1877), .Z(n1876) );
  BUFFD0 U1895 ( .I(n1878), .Z(n1877) );
  BUFFD0 U1896 ( .I(n1879), .Z(n1878) );
  BUFFD0 U1897 ( .I(n1880), .Z(n1879) );
  BUFFD0 U1898 ( .I(n1881), .Z(n1880) );
  BUFFD0 U1899 ( .I(n1882), .Z(n1881) );
  BUFFD0 U1900 ( .I(n1883), .Z(n1882) );
  BUFFD0 U1901 ( .I(n1884), .Z(n1883) );
  BUFFD0 U1902 ( .I(n1885), .Z(n1884) );
  BUFFD0 U1903 ( .I(n1886), .Z(n1885) );
  BUFFD0 U1904 ( .I(n1887), .Z(n1886) );
  BUFFD0 U1905 ( .I(n1888), .Z(n1887) );
  BUFFD0 U1906 ( .I(n1889), .Z(n1888) );
  BUFFD0 U1907 ( .I(n1890), .Z(n1889) );
  BUFFD0 U1908 ( .I(n1891), .Z(n1890) );
  BUFFD0 U1909 ( .I(n1892), .Z(n1891) );
  BUFFD0 U1910 ( .I(n1893), .Z(n1892) );
  BUFFD0 U1911 ( .I(n1894), .Z(n1893) );
  BUFFD0 U1912 ( .I(n1895), .Z(n1894) );
  BUFFD0 U1913 ( .I(n1896), .Z(n1895) );
  BUFFD0 U1914 ( .I(n1897), .Z(n1896) );
  BUFFD0 U1915 ( .I(N61), .Z(n1897) );
  BUFFD0 U1916 ( .I(n1899), .Z(n1898) );
  BUFFD0 U1917 ( .I(n1900), .Z(n1899) );
  BUFFD0 U1918 ( .I(n1901), .Z(n1900) );
  BUFFD0 U1919 ( .I(n1902), .Z(n1901) );
  BUFFD0 U1920 ( .I(n1903), .Z(n1902) );
  BUFFD0 U1921 ( .I(n1904), .Z(n1903) );
  BUFFD0 U1922 ( .I(n1905), .Z(n1904) );
  BUFFD0 U1923 ( .I(n1906), .Z(n1905) );
  BUFFD0 U1924 ( .I(n1907), .Z(n1906) );
  BUFFD0 U1925 ( .I(n1908), .Z(n1907) );
  BUFFD0 U1926 ( .I(n1909), .Z(n1908) );
  BUFFD0 U1927 ( .I(n1910), .Z(n1909) );
  BUFFD0 U1928 ( .I(n1911), .Z(n1910) );
  BUFFD0 U1929 ( .I(n1912), .Z(n1911) );
  BUFFD0 U1930 ( .I(n1913), .Z(n1912) );
  BUFFD0 U1931 ( .I(n1914), .Z(n1913) );
  BUFFD0 U1932 ( .I(n1915), .Z(n1914) );
  BUFFD0 U1933 ( .I(n1916), .Z(n1915) );
  BUFFD0 U1934 ( .I(n1917), .Z(n1916) );
  BUFFD0 U1935 ( .I(n1918), .Z(n1917) );
  BUFFD0 U1936 ( .I(n1919), .Z(n1918) );
  BUFFD0 U1937 ( .I(n1920), .Z(n1919) );
  BUFFD0 U1938 ( .I(n1921), .Z(n1920) );
  BUFFD0 U1939 ( .I(n1922), .Z(n1921) );
  BUFFD0 U1940 ( .I(n1923), .Z(n1922) );
  BUFFD0 U1941 ( .I(n1924), .Z(n1923) );
  BUFFD0 U1942 ( .I(n1925), .Z(n1924) );
  BUFFD0 U1943 ( .I(n1926), .Z(n1925) );
  BUFFD0 U1944 ( .I(n1927), .Z(n1926) );
  BUFFD0 U1945 ( .I(n1928), .Z(n1927) );
  BUFFD0 U1946 ( .I(n1929), .Z(n1928) );
  BUFFD0 U1947 ( .I(n1930), .Z(n1929) );
  BUFFD0 U1948 ( .I(n1931), .Z(n1930) );
  BUFFD0 U1949 ( .I(n1932), .Z(n1931) );
  BUFFD0 U1950 ( .I(n1933), .Z(n1932) );
  BUFFD0 U1951 ( .I(n1934), .Z(n1933) );
  BUFFD0 U1952 ( .I(n1935), .Z(n1934) );
  BUFFD0 U1953 ( .I(n1936), .Z(n1935) );
  BUFFD0 U1954 ( .I(n1937), .Z(n1936) );
  BUFFD0 U1955 ( .I(n1938), .Z(n1937) );
  BUFFD0 U1956 ( .I(n1939), .Z(n1938) );
  BUFFD0 U1957 ( .I(n1940), .Z(n1939) );
  BUFFD0 U1958 ( .I(n1941), .Z(n1940) );
  BUFFD0 U1959 ( .I(n1942), .Z(n1941) );
  BUFFD0 U1960 ( .I(n1943), .Z(n1942) );
  BUFFD0 U1961 ( .I(n1944), .Z(n1943) );
  BUFFD0 U1962 ( .I(n1945), .Z(n1944) );
  BUFFD0 U1963 ( .I(n1946), .Z(n1945) );
  BUFFD0 U1964 ( .I(n1947), .Z(n1946) );
  BUFFD0 U1965 ( .I(n1948), .Z(n1947) );
  BUFFD0 U1966 ( .I(n1949), .Z(n1948) );
  BUFFD0 U1967 ( .I(n1950), .Z(n1949) );
  BUFFD0 U1968 ( .I(n1951), .Z(n1950) );
  BUFFD0 U1969 ( .I(n1952), .Z(n1951) );
  BUFFD0 U1970 ( .I(n1953), .Z(n1952) );
  BUFFD0 U1971 ( .I(n1954), .Z(n1953) );
  BUFFD0 U1972 ( .I(n1955), .Z(n1954) );
  BUFFD0 U1973 ( .I(n1956), .Z(n1955) );
  BUFFD0 U1974 ( .I(n1957), .Z(n1956) );
  BUFFD0 U1975 ( .I(n1958), .Z(n1957) );
  BUFFD0 U1976 ( .I(n1959), .Z(n1958) );
  BUFFD0 U1977 ( .I(n1960), .Z(n1959) );
  BUFFD0 U1978 ( .I(n1961), .Z(n1960) );
  BUFFD0 U1979 ( .I(n1962), .Z(n1961) );
  BUFFD0 U1980 ( .I(n1963), .Z(n1962) );
  BUFFD0 U1981 ( .I(n1964), .Z(n1963) );
  BUFFD0 U1982 ( .I(n1965), .Z(n1964) );
  BUFFD0 U1983 ( .I(n1966), .Z(n1965) );
  BUFFD0 U1984 ( .I(n1967), .Z(n1966) );
  BUFFD0 U1985 ( .I(N62), .Z(n1967) );
  BUFFD0 U1986 ( .I(n1969), .Z(n1968) );
  BUFFD0 U1987 ( .I(n1970), .Z(n1969) );
  BUFFD0 U1988 ( .I(n1971), .Z(n1970) );
  BUFFD0 U1989 ( .I(n1972), .Z(n1971) );
  BUFFD0 U1990 ( .I(n1973), .Z(n1972) );
  BUFFD0 U1991 ( .I(n1974), .Z(n1973) );
  BUFFD0 U1992 ( .I(n1975), .Z(n1974) );
  BUFFD0 U1993 ( .I(n1976), .Z(n1975) );
  BUFFD0 U1994 ( .I(n1977), .Z(n1976) );
  BUFFD0 U1995 ( .I(n1978), .Z(n1977) );
  BUFFD0 U1996 ( .I(n1979), .Z(n1978) );
  BUFFD0 U1997 ( .I(n1980), .Z(n1979) );
  BUFFD0 U1998 ( .I(n1981), .Z(n1980) );
  BUFFD0 U1999 ( .I(n1982), .Z(n1981) );
  BUFFD0 U2000 ( .I(n1983), .Z(n1982) );
  BUFFD0 U2001 ( .I(n1984), .Z(n1983) );
  BUFFD0 U2002 ( .I(n1985), .Z(n1984) );
  BUFFD0 U2003 ( .I(n1986), .Z(n1985) );
  BUFFD0 U2004 ( .I(n1987), .Z(n1986) );
  BUFFD0 U2005 ( .I(n1988), .Z(n1987) );
  BUFFD0 U2006 ( .I(n1989), .Z(n1988) );
  BUFFD0 U2007 ( .I(n1990), .Z(n1989) );
  BUFFD0 U2008 ( .I(n1991), .Z(n1990) );
  BUFFD0 U2009 ( .I(n1992), .Z(n1991) );
  BUFFD0 U2010 ( .I(n1993), .Z(n1992) );
  BUFFD0 U2011 ( .I(n1994), .Z(n1993) );
  BUFFD0 U2012 ( .I(n1995), .Z(n1994) );
  BUFFD0 U2013 ( .I(n1996), .Z(n1995) );
  BUFFD0 U2014 ( .I(n1997), .Z(n1996) );
  BUFFD0 U2015 ( .I(n1998), .Z(n1997) );
  BUFFD0 U2016 ( .I(n1999), .Z(n1998) );
  BUFFD0 U2017 ( .I(n2000), .Z(n1999) );
  BUFFD0 U2018 ( .I(n2001), .Z(n2000) );
  BUFFD0 U2019 ( .I(n2002), .Z(n2001) );
  BUFFD0 U2020 ( .I(n2003), .Z(n2002) );
  BUFFD0 U2021 ( .I(n2004), .Z(n2003) );
  BUFFD0 U2022 ( .I(n2005), .Z(n2004) );
  BUFFD0 U2023 ( .I(n2006), .Z(n2005) );
  BUFFD0 U2024 ( .I(n2007), .Z(n2006) );
  BUFFD0 U2025 ( .I(n2008), .Z(n2007) );
  BUFFD0 U2026 ( .I(n2009), .Z(n2008) );
  BUFFD0 U2027 ( .I(n2010), .Z(n2009) );
  BUFFD0 U2028 ( .I(n2011), .Z(n2010) );
  BUFFD0 U2029 ( .I(n2012), .Z(n2011) );
  BUFFD0 U2030 ( .I(n2013), .Z(n2012) );
  BUFFD0 U2031 ( .I(n2014), .Z(n2013) );
  BUFFD0 U2032 ( .I(n2015), .Z(n2014) );
  BUFFD0 U2033 ( .I(n2016), .Z(n2015) );
  BUFFD0 U2034 ( .I(n2017), .Z(n2016) );
  BUFFD0 U2035 ( .I(n2018), .Z(n2017) );
  BUFFD0 U2036 ( .I(n2019), .Z(n2018) );
  BUFFD0 U2037 ( .I(n2020), .Z(n2019) );
  BUFFD0 U2038 ( .I(n2021), .Z(n2020) );
  BUFFD0 U2039 ( .I(n2022), .Z(n2021) );
  BUFFD0 U2040 ( .I(n2023), .Z(n2022) );
  BUFFD0 U2041 ( .I(n2024), .Z(n2023) );
  BUFFD0 U2042 ( .I(n2025), .Z(n2024) );
  BUFFD0 U2043 ( .I(n2026), .Z(n2025) );
  BUFFD0 U2044 ( .I(n2027), .Z(n2026) );
  BUFFD0 U2045 ( .I(n2028), .Z(n2027) );
  BUFFD0 U2046 ( .I(n2029), .Z(n2028) );
  BUFFD0 U2047 ( .I(n2030), .Z(n2029) );
  BUFFD0 U2048 ( .I(n2031), .Z(n2030) );
  BUFFD0 U2049 ( .I(n2032), .Z(n2031) );
  BUFFD0 U2050 ( .I(n2033), .Z(n2032) );
  BUFFD0 U2051 ( .I(n2034), .Z(n2033) );
  BUFFD0 U2052 ( .I(n2035), .Z(n2034) );
  BUFFD0 U2053 ( .I(n2036), .Z(n2035) );
  BUFFD0 U2054 ( .I(n2037), .Z(n2036) );
  BUFFD0 U2055 ( .I(N63), .Z(n2037) );
  BUFFD0 U2056 ( .I(n2039), .Z(n2038) );
  BUFFD0 U2057 ( .I(n2040), .Z(n2039) );
  BUFFD0 U2058 ( .I(n2041), .Z(n2040) );
  BUFFD0 U2059 ( .I(n2042), .Z(n2041) );
  BUFFD0 U2060 ( .I(n2043), .Z(n2042) );
  BUFFD0 U2061 ( .I(n2044), .Z(n2043) );
  BUFFD0 U2062 ( .I(n2045), .Z(n2044) );
  BUFFD0 U2063 ( .I(n2046), .Z(n2045) );
  BUFFD0 U2064 ( .I(n2047), .Z(n2046) );
  BUFFD0 U2065 ( .I(n2048), .Z(n2047) );
  BUFFD0 U2066 ( .I(n2049), .Z(n2048) );
  BUFFD0 U2067 ( .I(n2050), .Z(n2049) );
  BUFFD0 U2068 ( .I(n2051), .Z(n2050) );
  BUFFD0 U2069 ( .I(n2052), .Z(n2051) );
  BUFFD0 U2070 ( .I(n2053), .Z(n2052) );
  BUFFD0 U2071 ( .I(n2054), .Z(n2053) );
  BUFFD0 U2072 ( .I(n2055), .Z(n2054) );
  BUFFD0 U2073 ( .I(n2056), .Z(n2055) );
  BUFFD0 U2074 ( .I(n2057), .Z(n2056) );
  BUFFD0 U2075 ( .I(n2058), .Z(n2057) );
  BUFFD0 U2076 ( .I(n2059), .Z(n2058) );
  BUFFD0 U2077 ( .I(n2060), .Z(n2059) );
  BUFFD0 U2078 ( .I(n2061), .Z(n2060) );
  BUFFD0 U2079 ( .I(n2062), .Z(n2061) );
  BUFFD0 U2080 ( .I(n2063), .Z(n2062) );
  BUFFD0 U2081 ( .I(n2064), .Z(n2063) );
  BUFFD0 U2082 ( .I(n2065), .Z(n2064) );
  BUFFD0 U2083 ( .I(n2066), .Z(n2065) );
  BUFFD0 U2084 ( .I(n2067), .Z(n2066) );
  BUFFD0 U2085 ( .I(n2068), .Z(n2067) );
  BUFFD0 U2086 ( .I(n2069), .Z(n2068) );
  BUFFD0 U2087 ( .I(n2070), .Z(n2069) );
  BUFFD0 U2088 ( .I(n2071), .Z(n2070) );
  BUFFD0 U2089 ( .I(n2072), .Z(n2071) );
  BUFFD0 U2090 ( .I(n2073), .Z(n2072) );
  BUFFD0 U2091 ( .I(n2074), .Z(n2073) );
  BUFFD0 U2092 ( .I(n2075), .Z(n2074) );
  BUFFD0 U2093 ( .I(n2076), .Z(n2075) );
  BUFFD0 U2094 ( .I(n2077), .Z(n2076) );
  BUFFD0 U2095 ( .I(n2078), .Z(n2077) );
  BUFFD0 U2096 ( .I(n2079), .Z(n2078) );
  BUFFD0 U2097 ( .I(n2080), .Z(n2079) );
  BUFFD0 U2098 ( .I(n2081), .Z(n2080) );
  BUFFD0 U2099 ( .I(n2082), .Z(n2081) );
  BUFFD0 U2100 ( .I(n2083), .Z(n2082) );
  BUFFD0 U2101 ( .I(n2084), .Z(n2083) );
  BUFFD0 U2102 ( .I(n2085), .Z(n2084) );
  BUFFD0 U2103 ( .I(n2086), .Z(n2085) );
  BUFFD0 U2104 ( .I(n2087), .Z(n2086) );
  BUFFD0 U2105 ( .I(n2088), .Z(n2087) );
  BUFFD0 U2106 ( .I(n2089), .Z(n2088) );
  BUFFD0 U2107 ( .I(n2090), .Z(n2089) );
  BUFFD0 U2108 ( .I(n2091), .Z(n2090) );
  BUFFD0 U2109 ( .I(n2092), .Z(n2091) );
  BUFFD0 U2110 ( .I(n2093), .Z(n2092) );
  BUFFD0 U2111 ( .I(n2094), .Z(n2093) );
  BUFFD0 U2112 ( .I(n2095), .Z(n2094) );
  BUFFD0 U2113 ( .I(n2096), .Z(n2095) );
  BUFFD0 U2114 ( .I(n2097), .Z(n2096) );
  BUFFD0 U2115 ( .I(n2098), .Z(n2097) );
  BUFFD0 U2116 ( .I(n2099), .Z(n2098) );
  BUFFD0 U2117 ( .I(n2100), .Z(n2099) );
  BUFFD0 U2118 ( .I(n2101), .Z(n2100) );
  BUFFD0 U2119 ( .I(n2102), .Z(n2101) );
  BUFFD0 U2120 ( .I(n2103), .Z(n2102) );
  BUFFD0 U2121 ( .I(n2104), .Z(n2103) );
  BUFFD0 U2122 ( .I(n2105), .Z(n2104) );
  BUFFD0 U2123 ( .I(n2106), .Z(n2105) );
  BUFFD0 U2124 ( .I(n2107), .Z(n2106) );
  BUFFD0 U2125 ( .I(N64), .Z(n2107) );
  BUFFD0 U2126 ( .I(n2109), .Z(n2108) );
  BUFFD0 U2127 ( .I(n2110), .Z(n2109) );
  BUFFD0 U2128 ( .I(n2111), .Z(n2110) );
  BUFFD0 U2129 ( .I(n2112), .Z(n2111) );
  BUFFD0 U2130 ( .I(n2113), .Z(n2112) );
  BUFFD0 U2131 ( .I(n2114), .Z(n2113) );
  BUFFD0 U2132 ( .I(n2115), .Z(n2114) );
  BUFFD0 U2133 ( .I(n2116), .Z(n2115) );
  BUFFD0 U2134 ( .I(n2117), .Z(n2116) );
  BUFFD0 U2135 ( .I(n2118), .Z(n2117) );
  BUFFD0 U2136 ( .I(n2119), .Z(n2118) );
  BUFFD0 U2137 ( .I(n2120), .Z(n2119) );
  BUFFD0 U2138 ( .I(n2121), .Z(n2120) );
  BUFFD0 U2139 ( .I(n2122), .Z(n2121) );
  BUFFD0 U2140 ( .I(n2123), .Z(n2122) );
  BUFFD0 U2141 ( .I(n2124), .Z(n2123) );
  BUFFD0 U2142 ( .I(n2125), .Z(n2124) );
  BUFFD0 U2143 ( .I(n2126), .Z(n2125) );
  BUFFD0 U2144 ( .I(n2127), .Z(n2126) );
  BUFFD0 U2145 ( .I(n2128), .Z(n2127) );
  BUFFD0 U2146 ( .I(n2129), .Z(n2128) );
  BUFFD0 U2147 ( .I(n2130), .Z(n2129) );
  BUFFD0 U2148 ( .I(n2131), .Z(n2130) );
  BUFFD0 U2149 ( .I(n2132), .Z(n2131) );
  BUFFD0 U2150 ( .I(n2133), .Z(n2132) );
  BUFFD0 U2151 ( .I(n2134), .Z(n2133) );
  BUFFD0 U2152 ( .I(n2135), .Z(n2134) );
  BUFFD0 U2153 ( .I(n2136), .Z(n2135) );
  BUFFD0 U2154 ( .I(n2137), .Z(n2136) );
  BUFFD0 U2155 ( .I(n2138), .Z(n2137) );
  BUFFD0 U2156 ( .I(n2139), .Z(n2138) );
  BUFFD0 U2157 ( .I(n2140), .Z(n2139) );
  BUFFD0 U2158 ( .I(n2141), .Z(n2140) );
  BUFFD0 U2159 ( .I(n2142), .Z(n2141) );
  BUFFD0 U2160 ( .I(n2143), .Z(n2142) );
  BUFFD0 U2161 ( .I(n2144), .Z(n2143) );
  BUFFD0 U2162 ( .I(n2145), .Z(n2144) );
  BUFFD0 U2163 ( .I(n2146), .Z(n2145) );
  BUFFD0 U2164 ( .I(n2147), .Z(n2146) );
  BUFFD0 U2165 ( .I(n2148), .Z(n2147) );
  BUFFD0 U2166 ( .I(n2149), .Z(n2148) );
  BUFFD0 U2167 ( .I(n2150), .Z(n2149) );
  BUFFD0 U2168 ( .I(n2151), .Z(n2150) );
  BUFFD0 U2169 ( .I(n2152), .Z(n2151) );
  BUFFD0 U2170 ( .I(n2153), .Z(n2152) );
  BUFFD0 U2171 ( .I(n2154), .Z(n2153) );
  BUFFD0 U2172 ( .I(n2155), .Z(n2154) );
  BUFFD0 U2173 ( .I(n2156), .Z(n2155) );
  BUFFD0 U2174 ( .I(n2157), .Z(n2156) );
  BUFFD0 U2175 ( .I(n2158), .Z(n2157) );
  BUFFD0 U2176 ( .I(n2159), .Z(n2158) );
  BUFFD0 U2177 ( .I(n2160), .Z(n2159) );
  BUFFD0 U2178 ( .I(n2161), .Z(n2160) );
  BUFFD0 U2179 ( .I(n2162), .Z(n2161) );
  BUFFD0 U2180 ( .I(n2163), .Z(n2162) );
  BUFFD0 U2181 ( .I(n2164), .Z(n2163) );
  BUFFD0 U2182 ( .I(n2165), .Z(n2164) );
  BUFFD0 U2183 ( .I(n2166), .Z(n2165) );
  BUFFD0 U2184 ( .I(n2167), .Z(n2166) );
  BUFFD0 U2185 ( .I(n2168), .Z(n2167) );
  BUFFD0 U2186 ( .I(n2169), .Z(n2168) );
  BUFFD0 U2187 ( .I(n2170), .Z(n2169) );
  BUFFD0 U2188 ( .I(n2171), .Z(n2170) );
  BUFFD0 U2189 ( .I(n2172), .Z(n2171) );
  BUFFD0 U2190 ( .I(n2173), .Z(n2172) );
  BUFFD0 U2191 ( .I(n2174), .Z(n2173) );
  BUFFD0 U2192 ( .I(n2175), .Z(n2174) );
  BUFFD0 U2193 ( .I(n2176), .Z(n2175) );
  BUFFD0 U2194 ( .I(n2177), .Z(n2176) );
  BUFFD0 U2195 ( .I(N65), .Z(n2177) );
  BUFFD0 U2196 ( .I(n2179), .Z(n2178) );
  BUFFD0 U2197 ( .I(n2180), .Z(n2179) );
  BUFFD0 U2198 ( .I(n2181), .Z(n2180) );
  BUFFD0 U2199 ( .I(n2182), .Z(n2181) );
  BUFFD0 U2200 ( .I(n2183), .Z(n2182) );
  BUFFD0 U2201 ( .I(n2184), .Z(n2183) );
  BUFFD0 U2202 ( .I(n2185), .Z(n2184) );
  BUFFD0 U2203 ( .I(n2186), .Z(n2185) );
  BUFFD0 U2204 ( .I(n2187), .Z(n2186) );
  BUFFD0 U2205 ( .I(n2188), .Z(n2187) );
  BUFFD0 U2206 ( .I(n2189), .Z(n2188) );
  BUFFD0 U2207 ( .I(n2190), .Z(n2189) );
  BUFFD0 U2208 ( .I(n2191), .Z(n2190) );
  BUFFD0 U2209 ( .I(n2192), .Z(n2191) );
  BUFFD0 U2210 ( .I(n2193), .Z(n2192) );
  BUFFD0 U2211 ( .I(n2194), .Z(n2193) );
  BUFFD0 U2212 ( .I(n2195), .Z(n2194) );
  BUFFD0 U2213 ( .I(n2196), .Z(n2195) );
  BUFFD0 U2214 ( .I(n2197), .Z(n2196) );
  BUFFD0 U2215 ( .I(n2198), .Z(n2197) );
  BUFFD0 U2216 ( .I(n2199), .Z(n2198) );
  BUFFD0 U2217 ( .I(n2200), .Z(n2199) );
  BUFFD0 U2218 ( .I(n2201), .Z(n2200) );
  BUFFD0 U2219 ( .I(n2202), .Z(n2201) );
  BUFFD0 U2220 ( .I(n2203), .Z(n2202) );
  BUFFD0 U2221 ( .I(n2204), .Z(n2203) );
  BUFFD0 U2222 ( .I(n2205), .Z(n2204) );
  BUFFD0 U2223 ( .I(n2206), .Z(n2205) );
  BUFFD0 U2224 ( .I(n2207), .Z(n2206) );
  BUFFD0 U2225 ( .I(n2208), .Z(n2207) );
  BUFFD0 U2226 ( .I(n2209), .Z(n2208) );
  BUFFD0 U2227 ( .I(n2210), .Z(n2209) );
  BUFFD0 U2228 ( .I(n2211), .Z(n2210) );
  BUFFD0 U2229 ( .I(n2212), .Z(n2211) );
  BUFFD0 U2230 ( .I(n2213), .Z(n2212) );
  BUFFD0 U2231 ( .I(n2214), .Z(n2213) );
  BUFFD0 U2232 ( .I(n2215), .Z(n2214) );
  BUFFD0 U2233 ( .I(n2216), .Z(n2215) );
  BUFFD0 U2234 ( .I(n2217), .Z(n2216) );
  BUFFD0 U2235 ( .I(n2218), .Z(n2217) );
  BUFFD0 U2236 ( .I(n2219), .Z(n2218) );
  BUFFD0 U2237 ( .I(n2220), .Z(n2219) );
  BUFFD0 U2238 ( .I(n2221), .Z(n2220) );
  BUFFD0 U2239 ( .I(n2222), .Z(n2221) );
  BUFFD0 U2240 ( .I(n2223), .Z(n2222) );
  BUFFD0 U2241 ( .I(n2224), .Z(n2223) );
  BUFFD0 U2242 ( .I(n2225), .Z(n2224) );
  BUFFD0 U2243 ( .I(n2226), .Z(n2225) );
  BUFFD0 U2244 ( .I(n2227), .Z(n2226) );
  BUFFD0 U2245 ( .I(n2228), .Z(n2227) );
  BUFFD0 U2246 ( .I(n2229), .Z(n2228) );
  BUFFD0 U2247 ( .I(n2230), .Z(n2229) );
  BUFFD0 U2248 ( .I(n2231), .Z(n2230) );
  BUFFD0 U2249 ( .I(n2232), .Z(n2231) );
  BUFFD0 U2250 ( .I(n2233), .Z(n2232) );
  BUFFD0 U2251 ( .I(n2234), .Z(n2233) );
  BUFFD0 U2252 ( .I(n2235), .Z(n2234) );
  BUFFD0 U2253 ( .I(n2236), .Z(n2235) );
  BUFFD0 U2254 ( .I(n2237), .Z(n2236) );
  BUFFD0 U2255 ( .I(n2238), .Z(n2237) );
  BUFFD0 U2256 ( .I(n2239), .Z(n2238) );
  BUFFD0 U2257 ( .I(n2240), .Z(n2239) );
  BUFFD0 U2258 ( .I(n2241), .Z(n2240) );
  BUFFD0 U2259 ( .I(n2242), .Z(n2241) );
  BUFFD0 U2260 ( .I(n2243), .Z(n2242) );
  BUFFD0 U2261 ( .I(n2244), .Z(n2243) );
  BUFFD0 U2262 ( .I(n2245), .Z(n2244) );
  BUFFD0 U2263 ( .I(n2246), .Z(n2245) );
  BUFFD0 U2264 ( .I(n2247), .Z(n2246) );
  BUFFD0 U2265 ( .I(N66), .Z(n2247) );
  BUFFD0 U2266 ( .I(n2249), .Z(n2248) );
  BUFFD0 U2267 ( .I(n2250), .Z(n2249) );
  BUFFD0 U2268 ( .I(n2251), .Z(n2250) );
  BUFFD0 U2269 ( .I(n2252), .Z(n2251) );
  BUFFD0 U2270 ( .I(n2253), .Z(n2252) );
  BUFFD0 U2271 ( .I(n2254), .Z(n2253) );
  BUFFD0 U2272 ( .I(n2255), .Z(n2254) );
  BUFFD0 U2273 ( .I(n2256), .Z(n2255) );
  BUFFD0 U2274 ( .I(n2257), .Z(n2256) );
  BUFFD0 U2275 ( .I(n2258), .Z(n2257) );
  BUFFD0 U2276 ( .I(n2259), .Z(n2258) );
  BUFFD0 U2277 ( .I(n2260), .Z(n2259) );
  BUFFD0 U2278 ( .I(n2261), .Z(n2260) );
  BUFFD0 U2279 ( .I(n2262), .Z(n2261) );
  BUFFD0 U2280 ( .I(n2263), .Z(n2262) );
  BUFFD0 U2281 ( .I(n2264), .Z(n2263) );
  BUFFD0 U2282 ( .I(n2265), .Z(n2264) );
  BUFFD0 U2283 ( .I(n2266), .Z(n2265) );
  BUFFD0 U2284 ( .I(n2267), .Z(n2266) );
  BUFFD0 U2285 ( .I(n2268), .Z(n2267) );
  BUFFD0 U2286 ( .I(n2269), .Z(n2268) );
  BUFFD0 U2287 ( .I(n2270), .Z(n2269) );
  BUFFD0 U2288 ( .I(n2271), .Z(n2270) );
  BUFFD0 U2289 ( .I(n2272), .Z(n2271) );
  BUFFD0 U2290 ( .I(n2273), .Z(n2272) );
  BUFFD0 U2291 ( .I(n2274), .Z(n2273) );
  BUFFD0 U2292 ( .I(n2275), .Z(n2274) );
  BUFFD0 U2293 ( .I(n2276), .Z(n2275) );
  BUFFD0 U2294 ( .I(n2277), .Z(n2276) );
  BUFFD0 U2295 ( .I(n2278), .Z(n2277) );
  BUFFD0 U2296 ( .I(n2279), .Z(n2278) );
  BUFFD0 U2297 ( .I(n2280), .Z(n2279) );
  BUFFD0 U2298 ( .I(n2281), .Z(n2280) );
  BUFFD0 U2299 ( .I(n2282), .Z(n2281) );
  BUFFD0 U2300 ( .I(n2283), .Z(n2282) );
  BUFFD0 U2301 ( .I(n2284), .Z(n2283) );
  BUFFD0 U2302 ( .I(n2285), .Z(n2284) );
  BUFFD0 U2303 ( .I(n2286), .Z(n2285) );
  BUFFD0 U2304 ( .I(n2287), .Z(n2286) );
  BUFFD0 U2305 ( .I(n2288), .Z(n2287) );
  BUFFD0 U2306 ( .I(n2289), .Z(n2288) );
  BUFFD0 U2307 ( .I(n2290), .Z(n2289) );
  BUFFD0 U2308 ( .I(n2291), .Z(n2290) );
  BUFFD0 U2309 ( .I(n2292), .Z(n2291) );
  BUFFD0 U2310 ( .I(n2293), .Z(n2292) );
  BUFFD0 U2311 ( .I(n2294), .Z(n2293) );
  BUFFD0 U2312 ( .I(n2295), .Z(n2294) );
  BUFFD0 U2313 ( .I(n2296), .Z(n2295) );
  BUFFD0 U2314 ( .I(n2297), .Z(n2296) );
  BUFFD0 U2315 ( .I(n2298), .Z(n2297) );
  BUFFD0 U2316 ( .I(n2299), .Z(n2298) );
  BUFFD0 U2317 ( .I(n2300), .Z(n2299) );
  BUFFD0 U2318 ( .I(n2301), .Z(n2300) );
  BUFFD0 U2319 ( .I(n2302), .Z(n2301) );
  BUFFD0 U2320 ( .I(n2303), .Z(n2302) );
  BUFFD0 U2321 ( .I(n2304), .Z(n2303) );
  BUFFD0 U2322 ( .I(n2305), .Z(n2304) );
  BUFFD0 U2323 ( .I(n2306), .Z(n2305) );
  BUFFD0 U2324 ( .I(n2307), .Z(n2306) );
  BUFFD0 U2325 ( .I(n2308), .Z(n2307) );
  BUFFD0 U2326 ( .I(n2309), .Z(n2308) );
  BUFFD0 U2327 ( .I(n2310), .Z(n2309) );
  BUFFD0 U2328 ( .I(n2311), .Z(n2310) );
  BUFFD0 U2329 ( .I(n2312), .Z(n2311) );
  BUFFD0 U2330 ( .I(n2313), .Z(n2312) );
  BUFFD0 U2331 ( .I(n2314), .Z(n2313) );
  BUFFD0 U2332 ( .I(n2315), .Z(n2314) );
  BUFFD0 U2333 ( .I(n2316), .Z(n2315) );
  BUFFD0 U2334 ( .I(n2317), .Z(n2316) );
  BUFFD0 U2335 ( .I(N67), .Z(n2317) );
  BUFFD0 U2336 ( .I(n2319), .Z(n2318) );
  BUFFD0 U2337 ( .I(n2320), .Z(n2319) );
  BUFFD0 U2338 ( .I(n2321), .Z(n2320) );
  BUFFD0 U2339 ( .I(n2322), .Z(n2321) );
  BUFFD0 U2340 ( .I(n2323), .Z(n2322) );
  BUFFD0 U2341 ( .I(n2324), .Z(n2323) );
  BUFFD0 U2342 ( .I(n2325), .Z(n2324) );
  BUFFD0 U2343 ( .I(n2326), .Z(n2325) );
  BUFFD0 U2344 ( .I(n2327), .Z(n2326) );
  BUFFD0 U2345 ( .I(n2328), .Z(n2327) );
  BUFFD0 U2346 ( .I(n2329), .Z(n2328) );
  BUFFD0 U2347 ( .I(n2330), .Z(n2329) );
  BUFFD0 U2348 ( .I(n2331), .Z(n2330) );
  BUFFD0 U2349 ( .I(n2332), .Z(n2331) );
  BUFFD0 U2350 ( .I(n2333), .Z(n2332) );
  BUFFD0 U2351 ( .I(n2334), .Z(n2333) );
  BUFFD0 U2352 ( .I(n2335), .Z(n2334) );
  BUFFD0 U2353 ( .I(n2336), .Z(n2335) );
  BUFFD0 U2354 ( .I(n2337), .Z(n2336) );
  BUFFD0 U2355 ( .I(n2338), .Z(n2337) );
  BUFFD0 U2356 ( .I(n2339), .Z(n2338) );
  BUFFD0 U2357 ( .I(n2340), .Z(n2339) );
  BUFFD0 U2358 ( .I(n2341), .Z(n2340) );
  BUFFD0 U2359 ( .I(n2342), .Z(n2341) );
  BUFFD0 U2360 ( .I(n2343), .Z(n2342) );
  BUFFD0 U2361 ( .I(n2344), .Z(n2343) );
  BUFFD0 U2362 ( .I(n2345), .Z(n2344) );
  BUFFD0 U2363 ( .I(n2346), .Z(n2345) );
  BUFFD0 U2364 ( .I(n2347), .Z(n2346) );
  BUFFD0 U2365 ( .I(n2348), .Z(n2347) );
  BUFFD0 U2366 ( .I(n2349), .Z(n2348) );
  BUFFD0 U2367 ( .I(n2350), .Z(n2349) );
  BUFFD0 U2368 ( .I(n2351), .Z(n2350) );
  BUFFD0 U2369 ( .I(n2352), .Z(n2351) );
  BUFFD0 U2370 ( .I(n2353), .Z(n2352) );
  BUFFD0 U2371 ( .I(n2354), .Z(n2353) );
  BUFFD0 U2372 ( .I(n2355), .Z(n2354) );
  BUFFD0 U2373 ( .I(n2356), .Z(n2355) );
  BUFFD0 U2374 ( .I(n2357), .Z(n2356) );
  BUFFD0 U2375 ( .I(n2358), .Z(n2357) );
  BUFFD0 U2376 ( .I(n2359), .Z(n2358) );
  BUFFD0 U2377 ( .I(n2360), .Z(n2359) );
  BUFFD0 U2378 ( .I(n2361), .Z(n2360) );
  BUFFD0 U2379 ( .I(n2362), .Z(n2361) );
  BUFFD0 U2380 ( .I(n2363), .Z(n2362) );
  BUFFD0 U2381 ( .I(n2364), .Z(n2363) );
  BUFFD0 U2382 ( .I(n2365), .Z(n2364) );
  BUFFD0 U2383 ( .I(n2366), .Z(n2365) );
  BUFFD0 U2384 ( .I(n2367), .Z(n2366) );
  BUFFD0 U2385 ( .I(n2368), .Z(n2367) );
  BUFFD0 U2386 ( .I(n2369), .Z(n2368) );
  BUFFD0 U2387 ( .I(n2370), .Z(n2369) );
  BUFFD0 U2388 ( .I(n2371), .Z(n2370) );
  BUFFD0 U2389 ( .I(n2372), .Z(n2371) );
  BUFFD0 U2390 ( .I(n2373), .Z(n2372) );
  BUFFD0 U2391 ( .I(n2374), .Z(n2373) );
  BUFFD0 U2392 ( .I(n2375), .Z(n2374) );
  BUFFD0 U2393 ( .I(n2376), .Z(n2375) );
  BUFFD0 U2394 ( .I(n2377), .Z(n2376) );
  BUFFD0 U2395 ( .I(n2378), .Z(n2377) );
  BUFFD0 U2396 ( .I(n2379), .Z(n2378) );
  BUFFD0 U2397 ( .I(n2380), .Z(n2379) );
  BUFFD0 U2398 ( .I(n2381), .Z(n2380) );
  BUFFD0 U2399 ( .I(n2382), .Z(n2381) );
  BUFFD0 U2400 ( .I(n2383), .Z(n2382) );
  BUFFD0 U2401 ( .I(n2384), .Z(n2383) );
  BUFFD0 U2402 ( .I(n2385), .Z(n2384) );
  BUFFD0 U2403 ( .I(n2386), .Z(n2385) );
  BUFFD0 U2404 ( .I(n2387), .Z(n2386) );
  BUFFD0 U2405 ( .I(N68), .Z(n2387) );
  BUFFD0 U2406 ( .I(n2389), .Z(n2388) );
  BUFFD0 U2407 ( .I(n2390), .Z(n2389) );
  BUFFD0 U2408 ( .I(n2391), .Z(n2390) );
  BUFFD0 U2409 ( .I(n2392), .Z(n2391) );
  BUFFD0 U2410 ( .I(n2393), .Z(n2392) );
  BUFFD0 U2411 ( .I(n2394), .Z(n2393) );
  BUFFD0 U2412 ( .I(n2395), .Z(n2394) );
  BUFFD0 U2413 ( .I(n2396), .Z(n2395) );
  BUFFD0 U2414 ( .I(n2397), .Z(n2396) );
  BUFFD0 U2415 ( .I(n2398), .Z(n2397) );
  BUFFD0 U2416 ( .I(n2399), .Z(n2398) );
  BUFFD0 U2417 ( .I(n2400), .Z(n2399) );
  BUFFD0 U2418 ( .I(n2401), .Z(n2400) );
  BUFFD0 U2419 ( .I(n2402), .Z(n2401) );
  BUFFD0 U2420 ( .I(n2403), .Z(n2402) );
  BUFFD0 U2421 ( .I(n2404), .Z(n2403) );
  BUFFD0 U2422 ( .I(n2405), .Z(n2404) );
  BUFFD0 U2423 ( .I(n2406), .Z(n2405) );
  BUFFD0 U2424 ( .I(n2407), .Z(n2406) );
  BUFFD0 U2425 ( .I(n2408), .Z(n2407) );
  BUFFD0 U2426 ( .I(n2409), .Z(n2408) );
  BUFFD0 U2427 ( .I(n2410), .Z(n2409) );
  BUFFD0 U2428 ( .I(n2411), .Z(n2410) );
  BUFFD0 U2429 ( .I(n2412), .Z(n2411) );
  BUFFD0 U2430 ( .I(n2413), .Z(n2412) );
  BUFFD0 U2431 ( .I(n2414), .Z(n2413) );
  BUFFD0 U2432 ( .I(n2415), .Z(n2414) );
  BUFFD0 U2433 ( .I(n2416), .Z(n2415) );
  BUFFD0 U2434 ( .I(n2417), .Z(n2416) );
  BUFFD0 U2435 ( .I(n2418), .Z(n2417) );
  BUFFD0 U2436 ( .I(n2419), .Z(n2418) );
  BUFFD0 U2437 ( .I(n2420), .Z(n2419) );
  BUFFD0 U2438 ( .I(n2421), .Z(n2420) );
  BUFFD0 U2439 ( .I(n2422), .Z(n2421) );
  BUFFD0 U2440 ( .I(n2423), .Z(n2422) );
  BUFFD0 U2441 ( .I(n2424), .Z(n2423) );
  BUFFD0 U2442 ( .I(n2425), .Z(n2424) );
  BUFFD0 U2443 ( .I(n2426), .Z(n2425) );
  BUFFD0 U2444 ( .I(n2427), .Z(n2426) );
  BUFFD0 U2445 ( .I(n2428), .Z(n2427) );
  BUFFD0 U2446 ( .I(n2429), .Z(n2428) );
  BUFFD0 U2447 ( .I(n2430), .Z(n2429) );
  BUFFD0 U2448 ( .I(n2431), .Z(n2430) );
  BUFFD0 U2449 ( .I(n2432), .Z(n2431) );
  BUFFD0 U2450 ( .I(n2433), .Z(n2432) );
  BUFFD0 U2451 ( .I(n2434), .Z(n2433) );
  BUFFD0 U2452 ( .I(n2435), .Z(n2434) );
  BUFFD0 U2453 ( .I(n2436), .Z(n2435) );
  BUFFD0 U2454 ( .I(n2437), .Z(n2436) );
  BUFFD0 U2455 ( .I(n2438), .Z(n2437) );
  BUFFD0 U2456 ( .I(n2439), .Z(n2438) );
  BUFFD0 U2457 ( .I(n2440), .Z(n2439) );
  BUFFD0 U2458 ( .I(n2441), .Z(n2440) );
  BUFFD0 U2459 ( .I(n2442), .Z(n2441) );
  BUFFD0 U2460 ( .I(n2443), .Z(n2442) );
  BUFFD0 U2461 ( .I(n2444), .Z(n2443) );
  BUFFD0 U2462 ( .I(n2445), .Z(n2444) );
  BUFFD0 U2463 ( .I(n2446), .Z(n2445) );
  BUFFD0 U2464 ( .I(n2447), .Z(n2446) );
  BUFFD0 U2465 ( .I(n2448), .Z(n2447) );
  BUFFD0 U2466 ( .I(n2449), .Z(n2448) );
  BUFFD0 U2467 ( .I(n2450), .Z(n2449) );
  BUFFD0 U2468 ( .I(n2451), .Z(n2450) );
  BUFFD0 U2469 ( .I(n2452), .Z(n2451) );
  BUFFD0 U2470 ( .I(n2453), .Z(n2452) );
  BUFFD0 U2471 ( .I(n2454), .Z(n2453) );
  BUFFD0 U2472 ( .I(n2455), .Z(n2454) );
  BUFFD0 U2473 ( .I(n2456), .Z(n2455) );
  BUFFD0 U2474 ( .I(n2457), .Z(n2456) );
  BUFFD0 U2475 ( .I(N69), .Z(n2457) );
  BUFFD0 U2476 ( .I(n2459), .Z(n2458) );
  BUFFD0 U2477 ( .I(n2460), .Z(n2459) );
  BUFFD0 U2478 ( .I(n2461), .Z(n2460) );
  BUFFD0 U2479 ( .I(n2462), .Z(n2461) );
  BUFFD0 U2480 ( .I(n2463), .Z(n2462) );
  BUFFD0 U2481 ( .I(n2464), .Z(n2463) );
  BUFFD0 U2482 ( .I(n2465), .Z(n2464) );
  BUFFD0 U2483 ( .I(n2466), .Z(n2465) );
  BUFFD0 U2484 ( .I(n2467), .Z(n2466) );
  BUFFD0 U2485 ( .I(n2468), .Z(n2467) );
  BUFFD0 U2486 ( .I(n2469), .Z(n2468) );
  BUFFD0 U2487 ( .I(n2470), .Z(n2469) );
  BUFFD0 U2488 ( .I(n2471), .Z(n2470) );
  BUFFD0 U2489 ( .I(n2472), .Z(n2471) );
  BUFFD0 U2490 ( .I(n2473), .Z(n2472) );
  BUFFD0 U2491 ( .I(n2474), .Z(n2473) );
  BUFFD0 U2492 ( .I(n2475), .Z(n2474) );
  BUFFD0 U2493 ( .I(n2476), .Z(n2475) );
  BUFFD0 U2494 ( .I(n2477), .Z(n2476) );
  BUFFD0 U2495 ( .I(n2478), .Z(n2477) );
  BUFFD0 U2496 ( .I(n2479), .Z(n2478) );
  BUFFD0 U2497 ( .I(n2480), .Z(n2479) );
  BUFFD0 U2498 ( .I(n2481), .Z(n2480) );
  BUFFD0 U2499 ( .I(n2482), .Z(n2481) );
  BUFFD0 U2500 ( .I(n2483), .Z(n2482) );
  BUFFD0 U2501 ( .I(n2484), .Z(n2483) );
  BUFFD0 U2502 ( .I(n2485), .Z(n2484) );
  BUFFD0 U2503 ( .I(n2486), .Z(n2485) );
  BUFFD0 U2504 ( .I(n2487), .Z(n2486) );
  BUFFD0 U2505 ( .I(n2488), .Z(n2487) );
  BUFFD0 U2506 ( .I(n2489), .Z(n2488) );
  BUFFD0 U2507 ( .I(n2490), .Z(n2489) );
  BUFFD0 U2508 ( .I(n2491), .Z(n2490) );
  BUFFD0 U2509 ( .I(n2492), .Z(n2491) );
  BUFFD0 U2510 ( .I(n2493), .Z(n2492) );
  BUFFD0 U2511 ( .I(n2494), .Z(n2493) );
  BUFFD0 U2512 ( .I(n2495), .Z(n2494) );
  BUFFD0 U2513 ( .I(n2496), .Z(n2495) );
  BUFFD0 U2514 ( .I(n2497), .Z(n2496) );
  BUFFD0 U2515 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2516 ( .I(n2499), .Z(n2498) );
  BUFFD0 U2517 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2518 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2519 ( .I(n2502), .Z(n2501) );
  BUFFD0 U2520 ( .I(n2503), .Z(n2502) );
  BUFFD0 U2521 ( .I(n2504), .Z(n2503) );
  BUFFD0 U2522 ( .I(n2505), .Z(n2504) );
  BUFFD0 U2523 ( .I(n2506), .Z(n2505) );
  BUFFD0 U2524 ( .I(n2507), .Z(n2506) );
  BUFFD0 U2525 ( .I(n2508), .Z(n2507) );
  BUFFD0 U2526 ( .I(n2509), .Z(n2508) );
  BUFFD0 U2527 ( .I(n2510), .Z(n2509) );
  BUFFD0 U2528 ( .I(n2511), .Z(n2510) );
  BUFFD0 U2529 ( .I(n2512), .Z(n2511) );
  BUFFD0 U2530 ( .I(n2513), .Z(n2512) );
  BUFFD0 U2531 ( .I(n2514), .Z(n2513) );
  BUFFD0 U2532 ( .I(n2515), .Z(n2514) );
  BUFFD0 U2533 ( .I(n2516), .Z(n2515) );
  BUFFD0 U2534 ( .I(n2517), .Z(n2516) );
  BUFFD0 U2535 ( .I(n2518), .Z(n2517) );
  BUFFD0 U2536 ( .I(n2519), .Z(n2518) );
  BUFFD0 U2537 ( .I(n2520), .Z(n2519) );
  BUFFD0 U2538 ( .I(n2521), .Z(n2520) );
  BUFFD0 U2539 ( .I(n2522), .Z(n2521) );
  BUFFD0 U2540 ( .I(n2523), .Z(n2522) );
  BUFFD0 U2541 ( .I(n2524), .Z(n2523) );
  BUFFD0 U2542 ( .I(n2525), .Z(n2524) );
  BUFFD0 U2543 ( .I(n2526), .Z(n2525) );
  BUFFD0 U2544 ( .I(n2527), .Z(n2526) );
  BUFFD0 U2545 ( .I(N70), .Z(n2527) );
  BUFFD0 U2546 ( .I(n2529), .Z(n2528) );
  BUFFD0 U2547 ( .I(n2530), .Z(n2529) );
  BUFFD0 U2548 ( .I(n2531), .Z(n2530) );
  BUFFD0 U2549 ( .I(n2532), .Z(n2531) );
  BUFFD0 U2550 ( .I(n2533), .Z(n2532) );
  BUFFD0 U2551 ( .I(n2534), .Z(n2533) );
  BUFFD0 U2552 ( .I(n2535), .Z(n2534) );
  BUFFD0 U2553 ( .I(n2536), .Z(n2535) );
  BUFFD0 U2554 ( .I(n2537), .Z(n2536) );
  BUFFD0 U2555 ( .I(n2538), .Z(n2537) );
  BUFFD0 U2556 ( .I(n2539), .Z(n2538) );
  BUFFD0 U2557 ( .I(n2540), .Z(n2539) );
  BUFFD0 U2558 ( .I(n2541), .Z(n2540) );
  BUFFD0 U2559 ( .I(n2542), .Z(n2541) );
  BUFFD0 U2560 ( .I(n2543), .Z(n2542) );
  BUFFD0 U2561 ( .I(n2544), .Z(n2543) );
  BUFFD0 U2562 ( .I(n2545), .Z(n2544) );
  BUFFD0 U2563 ( .I(n2546), .Z(n2545) );
  BUFFD0 U2564 ( .I(n2547), .Z(n2546) );
  BUFFD0 U2565 ( .I(n2548), .Z(n2547) );
  BUFFD0 U2566 ( .I(n2549), .Z(n2548) );
  BUFFD0 U2567 ( .I(n2550), .Z(n2549) );
  BUFFD0 U2568 ( .I(n2551), .Z(n2550) );
  BUFFD0 U2569 ( .I(n2552), .Z(n2551) );
  BUFFD0 U2570 ( .I(n2553), .Z(n2552) );
  BUFFD0 U2571 ( .I(n2554), .Z(n2553) );
  BUFFD0 U2572 ( .I(n2555), .Z(n2554) );
  BUFFD0 U2573 ( .I(n2556), .Z(n2555) );
  BUFFD0 U2574 ( .I(n2557), .Z(n2556) );
  BUFFD0 U2575 ( .I(n2558), .Z(n2557) );
  BUFFD0 U2576 ( .I(n2559), .Z(n2558) );
  BUFFD0 U2577 ( .I(n2560), .Z(n2559) );
  BUFFD0 U2578 ( .I(n2561), .Z(n2560) );
  BUFFD0 U2579 ( .I(n2562), .Z(n2561) );
  BUFFD0 U2580 ( .I(n2563), .Z(n2562) );
  BUFFD0 U2581 ( .I(n2564), .Z(n2563) );
  BUFFD0 U2582 ( .I(n2565), .Z(n2564) );
  BUFFD0 U2583 ( .I(n2566), .Z(n2565) );
  BUFFD0 U2584 ( .I(n2567), .Z(n2566) );
  BUFFD0 U2585 ( .I(n2568), .Z(n2567) );
  BUFFD0 U2586 ( .I(n2569), .Z(n2568) );
  BUFFD0 U2587 ( .I(n2570), .Z(n2569) );
  BUFFD0 U2588 ( .I(n2571), .Z(n2570) );
  BUFFD0 U2589 ( .I(n2572), .Z(n2571) );
  BUFFD0 U2590 ( .I(n2573), .Z(n2572) );
  BUFFD0 U2591 ( .I(n2574), .Z(n2573) );
  BUFFD0 U2592 ( .I(n2575), .Z(n2574) );
  BUFFD0 U2593 ( .I(n2576), .Z(n2575) );
  BUFFD0 U2594 ( .I(n2577), .Z(n2576) );
  BUFFD0 U2595 ( .I(n2578), .Z(n2577) );
  BUFFD0 U2596 ( .I(n2579), .Z(n2578) );
  BUFFD0 U2597 ( .I(n2580), .Z(n2579) );
  BUFFD0 U2598 ( .I(n2581), .Z(n2580) );
  BUFFD0 U2599 ( .I(n2582), .Z(n2581) );
  BUFFD0 U2600 ( .I(n2583), .Z(n2582) );
  BUFFD0 U2601 ( .I(n2584), .Z(n2583) );
  BUFFD0 U2602 ( .I(n2585), .Z(n2584) );
  BUFFD0 U2603 ( .I(n2586), .Z(n2585) );
  BUFFD0 U2604 ( .I(n2587), .Z(n2586) );
  BUFFD0 U2605 ( .I(n2588), .Z(n2587) );
  BUFFD0 U2606 ( .I(n2589), .Z(n2588) );
  BUFFD0 U2607 ( .I(n2590), .Z(n2589) );
  BUFFD0 U2608 ( .I(n2591), .Z(n2590) );
  BUFFD0 U2609 ( .I(n2592), .Z(n2591) );
  BUFFD0 U2610 ( .I(n2593), .Z(n2592) );
  BUFFD0 U2611 ( .I(n2594), .Z(n2593) );
  BUFFD0 U2612 ( .I(n2595), .Z(n2594) );
  BUFFD0 U2613 ( .I(n2596), .Z(n2595) );
  BUFFD0 U2614 ( .I(n2597), .Z(n2596) );
  BUFFD0 U2615 ( .I(N71), .Z(n2597) );
  BUFFD0 U2616 ( .I(n2599), .Z(n2598) );
  BUFFD0 U2617 ( .I(n2600), .Z(n2599) );
  BUFFD0 U2618 ( .I(n2601), .Z(n2600) );
  BUFFD0 U2619 ( .I(n2602), .Z(n2601) );
  BUFFD0 U2620 ( .I(n2603), .Z(n2602) );
  BUFFD0 U2621 ( .I(n2604), .Z(n2603) );
  BUFFD0 U2622 ( .I(n2605), .Z(n2604) );
  BUFFD0 U2623 ( .I(n2606), .Z(n2605) );
  BUFFD0 U2624 ( .I(n2607), .Z(n2606) );
  BUFFD0 U2625 ( .I(n2608), .Z(n2607) );
  BUFFD0 U2626 ( .I(n2609), .Z(n2608) );
  BUFFD0 U2627 ( .I(n2610), .Z(n2609) );
  BUFFD0 U2628 ( .I(n2611), .Z(n2610) );
  BUFFD0 U2629 ( .I(n2612), .Z(n2611) );
  BUFFD0 U2630 ( .I(n2613), .Z(n2612) );
  BUFFD0 U2631 ( .I(n2614), .Z(n2613) );
  BUFFD0 U2632 ( .I(n2615), .Z(n2614) );
  BUFFD0 U2633 ( .I(n2616), .Z(n2615) );
  BUFFD0 U2634 ( .I(n2617), .Z(n2616) );
  BUFFD0 U2635 ( .I(n2618), .Z(n2617) );
  BUFFD0 U2636 ( .I(n2619), .Z(n2618) );
  BUFFD0 U2637 ( .I(n2620), .Z(n2619) );
  BUFFD0 U2638 ( .I(n2621), .Z(n2620) );
  BUFFD0 U2639 ( .I(n2622), .Z(n2621) );
  BUFFD0 U2640 ( .I(n2623), .Z(n2622) );
  BUFFD0 U2641 ( .I(n2624), .Z(n2623) );
  BUFFD0 U2642 ( .I(n2625), .Z(n2624) );
  BUFFD0 U2643 ( .I(n2626), .Z(n2625) );
  BUFFD0 U2644 ( .I(n2627), .Z(n2626) );
  BUFFD0 U2645 ( .I(n2628), .Z(n2627) );
  BUFFD0 U2646 ( .I(n2629), .Z(n2628) );
  BUFFD0 U2647 ( .I(n2630), .Z(n2629) );
  BUFFD0 U2648 ( .I(n2631), .Z(n2630) );
  BUFFD0 U2649 ( .I(n2632), .Z(n2631) );
  BUFFD0 U2650 ( .I(n2633), .Z(n2632) );
  BUFFD0 U2651 ( .I(n2634), .Z(n2633) );
  BUFFD0 U2652 ( .I(n2635), .Z(n2634) );
  BUFFD0 U2653 ( .I(n2636), .Z(n2635) );
  BUFFD0 U2654 ( .I(n2637), .Z(n2636) );
  BUFFD0 U2655 ( .I(n2638), .Z(n2637) );
  BUFFD0 U2656 ( .I(n2639), .Z(n2638) );
  BUFFD0 U2657 ( .I(n2640), .Z(n2639) );
  BUFFD0 U2658 ( .I(n2641), .Z(n2640) );
  BUFFD0 U2659 ( .I(n2642), .Z(n2641) );
  BUFFD0 U2660 ( .I(n2643), .Z(n2642) );
  BUFFD0 U2661 ( .I(n2644), .Z(n2643) );
  BUFFD0 U2662 ( .I(n2645), .Z(n2644) );
  BUFFD0 U2663 ( .I(n2646), .Z(n2645) );
  BUFFD0 U2664 ( .I(n2647), .Z(n2646) );
  BUFFD0 U2665 ( .I(n2648), .Z(n2647) );
  BUFFD0 U2666 ( .I(n2649), .Z(n2648) );
  BUFFD0 U2667 ( .I(n2650), .Z(n2649) );
  BUFFD0 U2668 ( .I(n2651), .Z(n2650) );
  BUFFD0 U2669 ( .I(n2652), .Z(n2651) );
  BUFFD0 U2670 ( .I(n2653), .Z(n2652) );
  BUFFD0 U2671 ( .I(n2654), .Z(n2653) );
  BUFFD0 U2672 ( .I(n2655), .Z(n2654) );
  BUFFD0 U2673 ( .I(n2656), .Z(n2655) );
  BUFFD0 U2674 ( .I(n2657), .Z(n2656) );
  BUFFD0 U2675 ( .I(n2658), .Z(n2657) );
  BUFFD0 U2676 ( .I(n2659), .Z(n2658) );
  BUFFD0 U2677 ( .I(n2660), .Z(n2659) );
  BUFFD0 U2678 ( .I(n2661), .Z(n2660) );
  BUFFD0 U2679 ( .I(n2662), .Z(n2661) );
  BUFFD0 U2680 ( .I(n2663), .Z(n2662) );
  BUFFD0 U2681 ( .I(n2664), .Z(n2663) );
  BUFFD0 U2682 ( .I(n2665), .Z(n2664) );
  BUFFD0 U2683 ( .I(n2666), .Z(n2665) );
  BUFFD0 U2684 ( .I(n2667), .Z(n2666) );
  BUFFD0 U2685 ( .I(N72), .Z(n2667) );
  BUFFD0 U2686 ( .I(n2669), .Z(n2668) );
  BUFFD0 U2687 ( .I(n2670), .Z(n2669) );
  BUFFD0 U2688 ( .I(n2671), .Z(n2670) );
  BUFFD0 U2689 ( .I(n2672), .Z(n2671) );
  BUFFD0 U2690 ( .I(n2673), .Z(n2672) );
  BUFFD0 U2691 ( .I(n2674), .Z(n2673) );
  BUFFD0 U2692 ( .I(n2675), .Z(n2674) );
  BUFFD0 U2693 ( .I(n2676), .Z(n2675) );
  BUFFD0 U2694 ( .I(n2677), .Z(n2676) );
  BUFFD0 U2695 ( .I(n2678), .Z(n2677) );
  BUFFD0 U2696 ( .I(n2679), .Z(n2678) );
  BUFFD0 U2697 ( .I(n2680), .Z(n2679) );
  BUFFD0 U2698 ( .I(n2681), .Z(n2680) );
  BUFFD0 U2699 ( .I(n2682), .Z(n2681) );
  BUFFD0 U2700 ( .I(n2683), .Z(n2682) );
  BUFFD0 U2701 ( .I(n2684), .Z(n2683) );
  BUFFD0 U2702 ( .I(n2685), .Z(n2684) );
  BUFFD0 U2703 ( .I(n2686), .Z(n2685) );
  BUFFD0 U2704 ( .I(n2687), .Z(n2686) );
  BUFFD0 U2705 ( .I(n2688), .Z(n2687) );
  BUFFD0 U2706 ( .I(n2689), .Z(n2688) );
  BUFFD0 U2707 ( .I(n2690), .Z(n2689) );
  BUFFD0 U2708 ( .I(n2691), .Z(n2690) );
  BUFFD0 U2709 ( .I(n2692), .Z(n2691) );
  BUFFD0 U2710 ( .I(n2693), .Z(n2692) );
  BUFFD0 U2711 ( .I(n2694), .Z(n2693) );
  BUFFD0 U2712 ( .I(n2695), .Z(n2694) );
  BUFFD0 U2713 ( .I(n2696), .Z(n2695) );
  BUFFD0 U2714 ( .I(n2697), .Z(n2696) );
  BUFFD0 U2715 ( .I(n2698), .Z(n2697) );
  BUFFD0 U2716 ( .I(n2699), .Z(n2698) );
  BUFFD0 U2717 ( .I(n2700), .Z(n2699) );
  BUFFD0 U2718 ( .I(n2701), .Z(n2700) );
  BUFFD0 U2719 ( .I(n2702), .Z(n2701) );
  BUFFD0 U2720 ( .I(n2703), .Z(n2702) );
  BUFFD0 U2721 ( .I(n2704), .Z(n2703) );
  BUFFD0 U2722 ( .I(n2705), .Z(n2704) );
  BUFFD0 U2723 ( .I(n2706), .Z(n2705) );
  BUFFD0 U2724 ( .I(n2707), .Z(n2706) );
  BUFFD0 U2725 ( .I(n2708), .Z(n2707) );
  BUFFD0 U2726 ( .I(n2709), .Z(n2708) );
  BUFFD0 U2727 ( .I(n2710), .Z(n2709) );
  BUFFD0 U2728 ( .I(n2711), .Z(n2710) );
  BUFFD0 U2729 ( .I(n2712), .Z(n2711) );
  BUFFD0 U2730 ( .I(n2713), .Z(n2712) );
  BUFFD0 U2731 ( .I(n2714), .Z(n2713) );
  BUFFD0 U2732 ( .I(n2715), .Z(n2714) );
  BUFFD0 U2733 ( .I(n2716), .Z(n2715) );
  BUFFD0 U2734 ( .I(n2717), .Z(n2716) );
  BUFFD0 U2735 ( .I(n2718), .Z(n2717) );
  BUFFD0 U2736 ( .I(n2719), .Z(n2718) );
  BUFFD0 U2737 ( .I(n2720), .Z(n2719) );
  BUFFD0 U2738 ( .I(n2721), .Z(n2720) );
  BUFFD0 U2739 ( .I(n2722), .Z(n2721) );
  BUFFD0 U2740 ( .I(n2723), .Z(n2722) );
  BUFFD0 U2741 ( .I(n2724), .Z(n2723) );
  BUFFD0 U2742 ( .I(n2725), .Z(n2724) );
  BUFFD0 U2743 ( .I(n2726), .Z(n2725) );
  BUFFD0 U2744 ( .I(n2727), .Z(n2726) );
  BUFFD0 U2745 ( .I(n2728), .Z(n2727) );
  BUFFD0 U2746 ( .I(n2729), .Z(n2728) );
  BUFFD0 U2747 ( .I(n2730), .Z(n2729) );
  BUFFD0 U2748 ( .I(n2731), .Z(n2730) );
  BUFFD0 U2749 ( .I(n2732), .Z(n2731) );
  BUFFD0 U2750 ( .I(n2733), .Z(n2732) );
  BUFFD0 U2751 ( .I(n2734), .Z(n2733) );
  BUFFD0 U2752 ( .I(n2735), .Z(n2734) );
  BUFFD0 U2753 ( .I(n2736), .Z(n2735) );
  BUFFD0 U2754 ( .I(n2737), .Z(n2736) );
  BUFFD0 U2755 ( .I(N73), .Z(n2737) );
  BUFFD0 U2756 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2757 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2758 ( .I(n2741), .Z(n2740) );
  BUFFD0 U2759 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2760 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2761 ( .I(n2744), .Z(n2743) );
  BUFFD0 U2762 ( .I(n2745), .Z(n2744) );
  BUFFD0 U2763 ( .I(n2746), .Z(n2745) );
  BUFFD0 U2764 ( .I(n2747), .Z(n2746) );
  BUFFD0 U2765 ( .I(n2748), .Z(n2747) );
  BUFFD0 U2766 ( .I(n2749), .Z(n2748) );
  BUFFD0 U2767 ( .I(n2750), .Z(n2749) );
  BUFFD0 U2768 ( .I(n2751), .Z(n2750) );
  BUFFD0 U2769 ( .I(n2752), .Z(n2751) );
  BUFFD0 U2770 ( .I(n2753), .Z(n2752) );
  BUFFD0 U2771 ( .I(n2754), .Z(n2753) );
  BUFFD0 U2772 ( .I(n2755), .Z(n2754) );
  BUFFD0 U2773 ( .I(n2756), .Z(n2755) );
  BUFFD0 U2774 ( .I(n2757), .Z(n2756) );
  BUFFD0 U2775 ( .I(n2758), .Z(n2757) );
  BUFFD0 U2776 ( .I(n2759), .Z(n2758) );
  BUFFD0 U2777 ( .I(n2760), .Z(n2759) );
  BUFFD0 U2778 ( .I(n2761), .Z(n2760) );
  BUFFD0 U2779 ( .I(n2762), .Z(n2761) );
  BUFFD0 U2780 ( .I(n2763), .Z(n2762) );
  BUFFD0 U2781 ( .I(n2764), .Z(n2763) );
  BUFFD0 U2782 ( .I(n2765), .Z(n2764) );
  BUFFD0 U2783 ( .I(n2766), .Z(n2765) );
  BUFFD0 U2784 ( .I(n2767), .Z(n2766) );
  BUFFD0 U2785 ( .I(n2768), .Z(n2767) );
  BUFFD0 U2786 ( .I(n2769), .Z(n2768) );
  BUFFD0 U2787 ( .I(n2770), .Z(n2769) );
  BUFFD0 U2788 ( .I(n2771), .Z(n2770) );
  BUFFD0 U2789 ( .I(n2772), .Z(n2771) );
  BUFFD0 U2790 ( .I(n2773), .Z(n2772) );
  BUFFD0 U2791 ( .I(n2774), .Z(n2773) );
  BUFFD0 U2792 ( .I(n2775), .Z(n2774) );
  BUFFD0 U2793 ( .I(n2776), .Z(n2775) );
  BUFFD0 U2794 ( .I(n2777), .Z(n2776) );
  BUFFD0 U2795 ( .I(n2778), .Z(n2777) );
  BUFFD0 U2796 ( .I(n2779), .Z(n2778) );
  BUFFD0 U2797 ( .I(n2780), .Z(n2779) );
  BUFFD0 U2798 ( .I(n2781), .Z(n2780) );
  BUFFD0 U2799 ( .I(n2782), .Z(n2781) );
  BUFFD0 U2800 ( .I(n2783), .Z(n2782) );
  BUFFD0 U2801 ( .I(n2784), .Z(n2783) );
  BUFFD0 U2802 ( .I(n2785), .Z(n2784) );
  BUFFD0 U2803 ( .I(n2786), .Z(n2785) );
  BUFFD0 U2804 ( .I(n2787), .Z(n2786) );
  BUFFD0 U2805 ( .I(n2788), .Z(n2787) );
  BUFFD0 U2806 ( .I(n2789), .Z(n2788) );
  BUFFD0 U2807 ( .I(n2790), .Z(n2789) );
  BUFFD0 U2808 ( .I(n2791), .Z(n2790) );
  BUFFD0 U2809 ( .I(n2792), .Z(n2791) );
  BUFFD0 U2810 ( .I(n2793), .Z(n2792) );
  BUFFD0 U2811 ( .I(n2794), .Z(n2793) );
  BUFFD0 U2812 ( .I(n2795), .Z(n2794) );
  BUFFD0 U2813 ( .I(n2796), .Z(n2795) );
  BUFFD0 U2814 ( .I(n2797), .Z(n2796) );
  BUFFD0 U2815 ( .I(n2798), .Z(n2797) );
  BUFFD0 U2816 ( .I(n2799), .Z(n2798) );
  BUFFD0 U2817 ( .I(n2800), .Z(n2799) );
  BUFFD0 U2818 ( .I(n2801), .Z(n2800) );
  BUFFD0 U2819 ( .I(n2802), .Z(n2801) );
  BUFFD0 U2820 ( .I(n2803), .Z(n2802) );
  BUFFD0 U2821 ( .I(n2804), .Z(n2803) );
  BUFFD0 U2822 ( .I(n2805), .Z(n2804) );
  BUFFD0 U2823 ( .I(n2806), .Z(n2805) );
  BUFFD0 U2824 ( .I(n2807), .Z(n2806) );
  BUFFD0 U2825 ( .I(N74), .Z(n2807) );
  BUFFD0 U2826 ( .I(n2809), .Z(n2808) );
  BUFFD0 U2827 ( .I(n2810), .Z(n2809) );
  BUFFD0 U2828 ( .I(n2811), .Z(n2810) );
  BUFFD0 U2829 ( .I(n2812), .Z(n2811) );
  BUFFD0 U2830 ( .I(n2813), .Z(n2812) );
  BUFFD0 U2831 ( .I(n2814), .Z(n2813) );
  BUFFD0 U2832 ( .I(n2815), .Z(n2814) );
  BUFFD0 U2833 ( .I(n2816), .Z(n2815) );
  BUFFD0 U2834 ( .I(n2817), .Z(n2816) );
  BUFFD0 U2835 ( .I(n2818), .Z(n2817) );
  BUFFD0 U2836 ( .I(n2819), .Z(n2818) );
  BUFFD0 U2837 ( .I(n2820), .Z(n2819) );
  BUFFD0 U2838 ( .I(n2821), .Z(n2820) );
  BUFFD0 U2839 ( .I(n2822), .Z(n2821) );
  BUFFD0 U2840 ( .I(n2823), .Z(n2822) );
  BUFFD0 U2841 ( .I(n2824), .Z(n2823) );
  BUFFD0 U2842 ( .I(n2825), .Z(n2824) );
  BUFFD0 U2843 ( .I(n2826), .Z(n2825) );
  BUFFD0 U2844 ( .I(n2827), .Z(n2826) );
  BUFFD0 U2845 ( .I(n2828), .Z(n2827) );
  BUFFD0 U2846 ( .I(n2829), .Z(n2828) );
  BUFFD0 U2847 ( .I(n2830), .Z(n2829) );
  BUFFD0 U2848 ( .I(n2831), .Z(n2830) );
  BUFFD0 U2849 ( .I(n2832), .Z(n2831) );
  BUFFD0 U2850 ( .I(n2833), .Z(n2832) );
  BUFFD0 U2851 ( .I(n2834), .Z(n2833) );
  BUFFD0 U2852 ( .I(n2835), .Z(n2834) );
  BUFFD0 U2853 ( .I(n2836), .Z(n2835) );
  BUFFD0 U2854 ( .I(n2837), .Z(n2836) );
  BUFFD0 U2855 ( .I(n2838), .Z(n2837) );
  BUFFD0 U2856 ( .I(n2839), .Z(n2838) );
  BUFFD0 U2857 ( .I(n2840), .Z(n2839) );
  BUFFD0 U2858 ( .I(n2841), .Z(n2840) );
  BUFFD0 U2859 ( .I(n2842), .Z(n2841) );
  BUFFD0 U2860 ( .I(n2843), .Z(n2842) );
  BUFFD0 U2861 ( .I(n2844), .Z(n2843) );
  BUFFD0 U2862 ( .I(n2845), .Z(n2844) );
  BUFFD0 U2863 ( .I(n2846), .Z(n2845) );
  BUFFD0 U2864 ( .I(n2847), .Z(n2846) );
  BUFFD0 U2865 ( .I(n2848), .Z(n2847) );
  BUFFD0 U2866 ( .I(n2849), .Z(n2848) );
  BUFFD0 U2867 ( .I(n2850), .Z(n2849) );
  BUFFD0 U2868 ( .I(n2851), .Z(n2850) );
  BUFFD0 U2869 ( .I(n2852), .Z(n2851) );
  BUFFD0 U2870 ( .I(n2853), .Z(n2852) );
  BUFFD0 U2871 ( .I(n2854), .Z(n2853) );
  BUFFD0 U2872 ( .I(n2855), .Z(n2854) );
  BUFFD0 U2873 ( .I(n2856), .Z(n2855) );
  BUFFD0 U2874 ( .I(n2857), .Z(n2856) );
  BUFFD0 U2875 ( .I(n2858), .Z(n2857) );
  BUFFD0 U2876 ( .I(n2859), .Z(n2858) );
  BUFFD0 U2877 ( .I(n2860), .Z(n2859) );
  BUFFD0 U2878 ( .I(n2861), .Z(n2860) );
  BUFFD0 U2879 ( .I(n2862), .Z(n2861) );
  BUFFD0 U2880 ( .I(n2863), .Z(n2862) );
  BUFFD0 U2881 ( .I(n2864), .Z(n2863) );
  BUFFD0 U2882 ( .I(n2865), .Z(n2864) );
  BUFFD0 U2883 ( .I(n2866), .Z(n2865) );
  BUFFD0 U2884 ( .I(n2867), .Z(n2866) );
  BUFFD0 U2885 ( .I(n2868), .Z(n2867) );
  BUFFD0 U2886 ( .I(n2869), .Z(n2868) );
  BUFFD0 U2887 ( .I(n2870), .Z(n2869) );
  BUFFD0 U2888 ( .I(n2871), .Z(n2870) );
  BUFFD0 U2889 ( .I(n2872), .Z(n2871) );
  BUFFD0 U2890 ( .I(n2873), .Z(n2872) );
  BUFFD0 U2891 ( .I(n2874), .Z(n2873) );
  BUFFD0 U2892 ( .I(n2875), .Z(n2874) );
  BUFFD0 U2893 ( .I(n2876), .Z(n2875) );
  BUFFD0 U2894 ( .I(n2877), .Z(n2876) );
  BUFFD0 U2895 ( .I(N75), .Z(n2877) );
  BUFFD0 U2896 ( .I(n2879), .Z(n2878) );
  BUFFD0 U2897 ( .I(n2880), .Z(n2879) );
  BUFFD0 U2898 ( .I(n2883), .Z(n2880) );
  BUFFD0 U2899 ( .I(n3501), .Z(n2881) );
  BUFFD0 U2900 ( .I(n2881), .Z(n2882) );
  BUFFD0 U2901 ( .I(n2884), .Z(n2883) );
  BUFFD0 U2902 ( .I(n2885), .Z(n2884) );
  BUFFD0 U2903 ( .I(n2886), .Z(n2885) );
  BUFFD0 U2904 ( .I(n2887), .Z(n2886) );
  BUFFD0 U2905 ( .I(n2888), .Z(n2887) );
  BUFFD0 U2906 ( .I(n2889), .Z(n2888) );
  BUFFD0 U2907 ( .I(n2890), .Z(n2889) );
  BUFFD0 U2908 ( .I(n2891), .Z(n2890) );
  BUFFD0 U2909 ( .I(n2892), .Z(n2891) );
  BUFFD0 U2910 ( .I(n2893), .Z(n2892) );
  BUFFD0 U2911 ( .I(n2894), .Z(n2893) );
  BUFFD0 U2912 ( .I(n2895), .Z(n2894) );
  BUFFD0 U2913 ( .I(n2896), .Z(n2895) );
  BUFFD0 U2914 ( .I(n2897), .Z(n2896) );
  BUFFD0 U2915 ( .I(n2898), .Z(n2897) );
  BUFFD0 U2916 ( .I(n2899), .Z(n2898) );
  BUFFD0 U2917 ( .I(n2900), .Z(n2899) );
  BUFFD0 U2918 ( .I(n2901), .Z(n2900) );
  BUFFD0 U2919 ( .I(n2902), .Z(n2901) );
  BUFFD0 U2920 ( .I(n2903), .Z(n2902) );
  BUFFD0 U2921 ( .I(n2904), .Z(n2903) );
  BUFFD0 U2922 ( .I(n2905), .Z(n2904) );
  BUFFD0 U2923 ( .I(n2906), .Z(n2905) );
  BUFFD0 U2924 ( .I(n2907), .Z(n2906) );
  BUFFD0 U2925 ( .I(n2908), .Z(n2907) );
  BUFFD0 U2926 ( .I(n2909), .Z(n2908) );
  BUFFD0 U2927 ( .I(n2910), .Z(n2909) );
  BUFFD0 U2928 ( .I(n2911), .Z(n2910) );
  BUFFD0 U2929 ( .I(n2912), .Z(n2911) );
  BUFFD0 U2930 ( .I(n2913), .Z(n2912) );
  BUFFD0 U2931 ( .I(n2914), .Z(n2913) );
  BUFFD0 U2932 ( .I(n2915), .Z(n2914) );
  BUFFD0 U2933 ( .I(n2916), .Z(n2915) );
  BUFFD0 U2934 ( .I(n2917), .Z(n2916) );
  BUFFD0 U2935 ( .I(n2918), .Z(n2917) );
  BUFFD0 U2936 ( .I(n2919), .Z(n2918) );
  BUFFD0 U2937 ( .I(n2920), .Z(n2919) );
  BUFFD0 U2938 ( .I(n2921), .Z(n2920) );
  BUFFD0 U2939 ( .I(n2922), .Z(n2921) );
  BUFFD0 U2940 ( .I(n2923), .Z(n2922) );
  BUFFD0 U2941 ( .I(n2924), .Z(n2923) );
  BUFFD0 U2942 ( .I(n2925), .Z(n2924) );
  BUFFD0 U2943 ( .I(n2926), .Z(n2925) );
  BUFFD0 U2944 ( .I(n2927), .Z(n2926) );
  BUFFD0 U2945 ( .I(n2928), .Z(n2927) );
  BUFFD0 U2946 ( .I(n2929), .Z(n2928) );
  BUFFD0 U2947 ( .I(n2930), .Z(n2929) );
  BUFFD0 U2948 ( .I(n2931), .Z(n2930) );
  BUFFD0 U2949 ( .I(n2932), .Z(n2931) );
  BUFFD0 U2950 ( .I(n2933), .Z(n2932) );
  BUFFD0 U2951 ( .I(n2934), .Z(n2933) );
  BUFFD0 U2952 ( .I(n2935), .Z(n2934) );
  BUFFD0 U2953 ( .I(n2936), .Z(n2935) );
  BUFFD0 U2954 ( .I(n2937), .Z(n2936) );
  BUFFD0 U2955 ( .I(n2938), .Z(n2937) );
  BUFFD0 U2956 ( .I(n2939), .Z(n2938) );
  BUFFD0 U2957 ( .I(n2940), .Z(n2939) );
  BUFFD0 U2958 ( .I(n2941), .Z(n2940) );
  BUFFD0 U2959 ( .I(n2942), .Z(n2941) );
  BUFFD0 U2960 ( .I(n2943), .Z(n2942) );
  BUFFD0 U2961 ( .I(n2945), .Z(n2943) );
  BUFFD0 U2962 ( .I(N76), .Z(n2944) );
  BUFFD0 U2963 ( .I(n2946), .Z(n2945) );
  BUFFD0 U2964 ( .I(n2882), .Z(n2946) );
  BUFFD0 U2965 ( .I(n2948), .Z(n2947) );
  BUFFD0 U2966 ( .I(n2949), .Z(n2948) );
  BUFFD0 U2967 ( .I(n2950), .Z(n2949) );
  BUFFD0 U2968 ( .I(n2951), .Z(n2950) );
  BUFFD0 U2969 ( .I(n2952), .Z(n2951) );
  BUFFD0 U2970 ( .I(n2953), .Z(n2952) );
  BUFFD0 U2971 ( .I(n2954), .Z(n2953) );
  BUFFD0 U2972 ( .I(n2955), .Z(n2954) );
  BUFFD0 U2973 ( .I(n2956), .Z(n2955) );
  BUFFD0 U2974 ( .I(n2957), .Z(n2956) );
  BUFFD0 U2975 ( .I(n2958), .Z(n2957) );
  BUFFD0 U2976 ( .I(n2959), .Z(n2958) );
  BUFFD0 U2977 ( .I(n2960), .Z(n2959) );
  BUFFD0 U2978 ( .I(n2961), .Z(n2960) );
  BUFFD0 U2979 ( .I(n2962), .Z(n2961) );
  BUFFD0 U2980 ( .I(n2963), .Z(n2962) );
  BUFFD0 U2981 ( .I(n2964), .Z(n2963) );
  BUFFD0 U2982 ( .I(n2965), .Z(n2964) );
  BUFFD0 U2983 ( .I(n2966), .Z(n2965) );
  BUFFD0 U2984 ( .I(n2967), .Z(n2966) );
  BUFFD0 U2985 ( .I(n2968), .Z(n2967) );
  BUFFD0 U2986 ( .I(n2969), .Z(n2968) );
  BUFFD0 U2987 ( .I(n2970), .Z(n2969) );
  BUFFD0 U2988 ( .I(n2971), .Z(n2970) );
  BUFFD0 U2989 ( .I(n2972), .Z(n2971) );
  BUFFD0 U2990 ( .I(n2973), .Z(n2972) );
  BUFFD0 U2991 ( .I(n2974), .Z(n2973) );
  BUFFD0 U2992 ( .I(n2975), .Z(n2974) );
  BUFFD0 U2993 ( .I(n2976), .Z(n2975) );
  BUFFD0 U2994 ( .I(n2977), .Z(n2976) );
  BUFFD0 U2995 ( .I(n2978), .Z(n2977) );
  BUFFD0 U2996 ( .I(n2979), .Z(n2978) );
  BUFFD0 U2997 ( .I(n2980), .Z(n2979) );
  BUFFD0 U2998 ( .I(n2981), .Z(n2980) );
  BUFFD0 U2999 ( .I(n2982), .Z(n2981) );
  BUFFD0 U3000 ( .I(n2983), .Z(n2982) );
  BUFFD0 U3001 ( .I(n2984), .Z(n2983) );
  BUFFD0 U3002 ( .I(n2985), .Z(n2984) );
  BUFFD0 U3003 ( .I(n2986), .Z(n2985) );
  BUFFD0 U3004 ( .I(n2987), .Z(n2986) );
  BUFFD0 U3005 ( .I(n2988), .Z(n2987) );
  BUFFD0 U3006 ( .I(n2989), .Z(n2988) );
  BUFFD0 U3007 ( .I(n2990), .Z(n2989) );
  BUFFD0 U3008 ( .I(n2991), .Z(n2990) );
  BUFFD0 U3009 ( .I(n2992), .Z(n2991) );
  BUFFD0 U3010 ( .I(n2993), .Z(n2992) );
  BUFFD0 U3011 ( .I(n2994), .Z(n2993) );
  BUFFD0 U3012 ( .I(n2995), .Z(n2994) );
  BUFFD0 U3013 ( .I(n2996), .Z(n2995) );
  BUFFD0 U3014 ( .I(n2997), .Z(n2996) );
  BUFFD0 U3015 ( .I(n2998), .Z(n2997) );
  BUFFD0 U3016 ( .I(n2999), .Z(n2998) );
  BUFFD0 U3017 ( .I(n3000), .Z(n2999) );
  BUFFD0 U3018 ( .I(n3001), .Z(n3000) );
  BUFFD0 U3019 ( .I(n3002), .Z(n3001) );
  BUFFD0 U3020 ( .I(n3003), .Z(n3002) );
  BUFFD0 U3021 ( .I(n3004), .Z(n3003) );
  BUFFD0 U3022 ( .I(n3005), .Z(n3004) );
  BUFFD0 U3023 ( .I(n3006), .Z(n3005) );
  BUFFD0 U3024 ( .I(n3007), .Z(n3006) );
  BUFFD0 U3025 ( .I(n3008), .Z(n3007) );
  BUFFD0 U3026 ( .I(n3009), .Z(n3008) );
  BUFFD0 U3027 ( .I(n3010), .Z(n3009) );
  BUFFD0 U3028 ( .I(n3011), .Z(n3010) );
  BUFFD0 U3029 ( .I(n3012), .Z(n3011) );
  BUFFD0 U3030 ( .I(n3013), .Z(n3012) );
  BUFFD0 U3031 ( .I(n3014), .Z(n3013) );
  BUFFD0 U3032 ( .I(n3015), .Z(n3014) );
  BUFFD0 U3033 ( .I(n3016), .Z(n3015) );
  BUFFD0 U3034 ( .I(N77), .Z(n3016) );
  BUFFD0 U3035 ( .I(n3018), .Z(n3017) );
  BUFFD0 U3036 ( .I(n3019), .Z(n3018) );
  BUFFD0 U3037 ( .I(n3020), .Z(n3019) );
  BUFFD0 U3038 ( .I(n3021), .Z(n3020) );
  BUFFD0 U3039 ( .I(n3022), .Z(n3021) );
  BUFFD0 U3040 ( .I(n3023), .Z(n3022) );
  BUFFD0 U3041 ( .I(n3024), .Z(n3023) );
  BUFFD0 U3042 ( .I(n3025), .Z(n3024) );
  BUFFD0 U3043 ( .I(n3026), .Z(n3025) );
  BUFFD0 U3044 ( .I(n3027), .Z(n3026) );
  BUFFD0 U3045 ( .I(n3028), .Z(n3027) );
  BUFFD0 U3046 ( .I(n3029), .Z(n3028) );
  BUFFD0 U3047 ( .I(n3030), .Z(n3029) );
  BUFFD0 U3048 ( .I(n3031), .Z(n3030) );
  BUFFD0 U3049 ( .I(n3032), .Z(n3031) );
  BUFFD0 U3050 ( .I(n3033), .Z(n3032) );
  BUFFD0 U3051 ( .I(n3034), .Z(n3033) );
  BUFFD0 U3052 ( .I(n3035), .Z(n3034) );
  BUFFD0 U3053 ( .I(n3036), .Z(n3035) );
  BUFFD0 U3054 ( .I(n3037), .Z(n3036) );
  BUFFD0 U3055 ( .I(n3038), .Z(n3037) );
  BUFFD0 U3056 ( .I(n3039), .Z(n3038) );
  BUFFD0 U3057 ( .I(n3040), .Z(n3039) );
  BUFFD0 U3058 ( .I(n3041), .Z(n3040) );
  BUFFD0 U3059 ( .I(n3042), .Z(n3041) );
  BUFFD0 U3060 ( .I(n3043), .Z(n3042) );
  BUFFD0 U3061 ( .I(n3044), .Z(n3043) );
  BUFFD0 U3062 ( .I(n3045), .Z(n3044) );
  BUFFD0 U3063 ( .I(n3046), .Z(n3045) );
  BUFFD0 U3064 ( .I(n3047), .Z(n3046) );
  BUFFD0 U3065 ( .I(n3048), .Z(n3047) );
  BUFFD0 U3066 ( .I(n3049), .Z(n3048) );
  BUFFD0 U3067 ( .I(n3050), .Z(n3049) );
  BUFFD0 U3068 ( .I(n3051), .Z(n3050) );
  BUFFD0 U3069 ( .I(n3052), .Z(n3051) );
  BUFFD0 U3070 ( .I(n3053), .Z(n3052) );
  BUFFD0 U3071 ( .I(n3054), .Z(n3053) );
  BUFFD0 U3072 ( .I(n3055), .Z(n3054) );
  BUFFD0 U3073 ( .I(n3056), .Z(n3055) );
  BUFFD0 U3074 ( .I(n3057), .Z(n3056) );
  BUFFD0 U3075 ( .I(n3058), .Z(n3057) );
  BUFFD0 U3076 ( .I(n3059), .Z(n3058) );
  BUFFD0 U3077 ( .I(n3060), .Z(n3059) );
  BUFFD0 U3078 ( .I(n3061), .Z(n3060) );
  BUFFD0 U3079 ( .I(n3062), .Z(n3061) );
  BUFFD0 U3080 ( .I(n3063), .Z(n3062) );
  BUFFD0 U3081 ( .I(n3064), .Z(n3063) );
  BUFFD0 U3082 ( .I(n3065), .Z(n3064) );
  BUFFD0 U3083 ( .I(n3066), .Z(n3065) );
  BUFFD0 U3084 ( .I(n3067), .Z(n3066) );
  BUFFD0 U3085 ( .I(n3068), .Z(n3067) );
  BUFFD0 U3086 ( .I(n3069), .Z(n3068) );
  BUFFD0 U3087 ( .I(n3070), .Z(n3069) );
  BUFFD0 U3088 ( .I(n3071), .Z(n3070) );
  BUFFD0 U3089 ( .I(n3072), .Z(n3071) );
  BUFFD0 U3090 ( .I(n3073), .Z(n3072) );
  BUFFD0 U3091 ( .I(n3074), .Z(n3073) );
  BUFFD0 U3092 ( .I(n3075), .Z(n3074) );
  BUFFD0 U3093 ( .I(n3076), .Z(n3075) );
  BUFFD0 U3094 ( .I(n3077), .Z(n3076) );
  BUFFD0 U3095 ( .I(n3078), .Z(n3077) );
  BUFFD0 U3096 ( .I(n3079), .Z(n3078) );
  BUFFD0 U3097 ( .I(n3080), .Z(n3079) );
  BUFFD0 U3098 ( .I(n3081), .Z(n3080) );
  BUFFD0 U3099 ( .I(n3082), .Z(n3081) );
  BUFFD0 U3100 ( .I(n3083), .Z(n3082) );
  BUFFD0 U3101 ( .I(n3084), .Z(n3083) );
  BUFFD0 U3102 ( .I(n3085), .Z(n3084) );
  BUFFD0 U3103 ( .I(n3086), .Z(n3085) );
  BUFFD0 U3104 ( .I(N78), .Z(n3086) );
  BUFFD0 U3105 ( .I(n3088), .Z(n3087) );
  BUFFD0 U3106 ( .I(n3089), .Z(n3088) );
  BUFFD0 U3107 ( .I(n3090), .Z(n3089) );
  BUFFD0 U3108 ( .I(n3091), .Z(n3090) );
  BUFFD0 U3109 ( .I(n3092), .Z(n3091) );
  BUFFD0 U3110 ( .I(n3093), .Z(n3092) );
  BUFFD0 U3111 ( .I(n3094), .Z(n3093) );
  BUFFD0 U3112 ( .I(n3095), .Z(n3094) );
  BUFFD0 U3113 ( .I(n3096), .Z(n3095) );
  BUFFD0 U3114 ( .I(n3097), .Z(n3096) );
  BUFFD0 U3115 ( .I(n3098), .Z(n3097) );
  BUFFD0 U3116 ( .I(n3099), .Z(n3098) );
  BUFFD0 U3117 ( .I(n3100), .Z(n3099) );
  BUFFD0 U3118 ( .I(n3101), .Z(n3100) );
  BUFFD0 U3119 ( .I(n3102), .Z(n3101) );
  BUFFD0 U3120 ( .I(n3103), .Z(n3102) );
  BUFFD0 U3121 ( .I(n3104), .Z(n3103) );
  BUFFD0 U3122 ( .I(n3105), .Z(n3104) );
  BUFFD0 U3123 ( .I(n3106), .Z(n3105) );
  BUFFD0 U3124 ( .I(n3107), .Z(n3106) );
  BUFFD0 U3125 ( .I(n3108), .Z(n3107) );
  BUFFD0 U3126 ( .I(n3109), .Z(n3108) );
  BUFFD0 U3127 ( .I(n3110), .Z(n3109) );
  BUFFD0 U3128 ( .I(n3111), .Z(n3110) );
  BUFFD0 U3129 ( .I(n3112), .Z(n3111) );
  BUFFD0 U3130 ( .I(n3113), .Z(n3112) );
  BUFFD0 U3131 ( .I(n3114), .Z(n3113) );
  BUFFD0 U3132 ( .I(n3115), .Z(n3114) );
  BUFFD0 U3133 ( .I(n3116), .Z(n3115) );
  BUFFD0 U3134 ( .I(n3117), .Z(n3116) );
  BUFFD0 U3135 ( .I(n3118), .Z(n3117) );
  BUFFD0 U3136 ( .I(n3119), .Z(n3118) );
  BUFFD0 U3137 ( .I(n3120), .Z(n3119) );
  BUFFD0 U3138 ( .I(n3121), .Z(n3120) );
  BUFFD0 U3139 ( .I(n3122), .Z(n3121) );
  BUFFD0 U3140 ( .I(n3123), .Z(n3122) );
  BUFFD0 U3141 ( .I(n3124), .Z(n3123) );
  BUFFD0 U3142 ( .I(n3125), .Z(n3124) );
  BUFFD0 U3143 ( .I(n3126), .Z(n3125) );
  BUFFD0 U3144 ( .I(n3127), .Z(n3126) );
  BUFFD0 U3145 ( .I(n3128), .Z(n3127) );
  BUFFD0 U3146 ( .I(n3129), .Z(n3128) );
  BUFFD0 U3147 ( .I(n3130), .Z(n3129) );
  BUFFD0 U3148 ( .I(n3131), .Z(n3130) );
  BUFFD0 U3149 ( .I(n3132), .Z(n3131) );
  BUFFD0 U3150 ( .I(n3133), .Z(n3132) );
  BUFFD0 U3151 ( .I(n3134), .Z(n3133) );
  BUFFD0 U3152 ( .I(n3135), .Z(n3134) );
  BUFFD0 U3153 ( .I(n3136), .Z(n3135) );
  BUFFD0 U3154 ( .I(n3137), .Z(n3136) );
  BUFFD0 U3155 ( .I(n3138), .Z(n3137) );
  BUFFD0 U3156 ( .I(n3139), .Z(n3138) );
  BUFFD0 U3157 ( .I(n3140), .Z(n3139) );
  BUFFD0 U3158 ( .I(n3141), .Z(n3140) );
  BUFFD0 U3159 ( .I(n3142), .Z(n3141) );
  BUFFD0 U3160 ( .I(n3143), .Z(n3142) );
  BUFFD0 U3161 ( .I(n3144), .Z(n3143) );
  BUFFD0 U3162 ( .I(n3145), .Z(n3144) );
  BUFFD0 U3163 ( .I(n3146), .Z(n3145) );
  BUFFD0 U3164 ( .I(n3147), .Z(n3146) );
  BUFFD0 U3165 ( .I(n3148), .Z(n3147) );
  BUFFD0 U3166 ( .I(n3149), .Z(n3148) );
  BUFFD0 U3167 ( .I(n3150), .Z(n3149) );
  BUFFD0 U3168 ( .I(n3151), .Z(n3150) );
  BUFFD0 U3169 ( .I(n3152), .Z(n3151) );
  BUFFD0 U3170 ( .I(n3153), .Z(n3152) );
  BUFFD0 U3171 ( .I(n3154), .Z(n3153) );
  BUFFD0 U3172 ( .I(n3155), .Z(n3154) );
  BUFFD0 U3173 ( .I(n3156), .Z(n3155) );
  BUFFD0 U3174 ( .I(N79), .Z(n3156) );
  BUFFD0 U3175 ( .I(n3158), .Z(n3157) );
  BUFFD0 U3176 ( .I(n3159), .Z(n3158) );
  BUFFD0 U3177 ( .I(n3160), .Z(n3159) );
  BUFFD0 U3178 ( .I(n3161), .Z(n3160) );
  BUFFD0 U3179 ( .I(n3162), .Z(n3161) );
  BUFFD0 U3180 ( .I(n3163), .Z(n3162) );
  BUFFD0 U3181 ( .I(n3164), .Z(n3163) );
  BUFFD0 U3182 ( .I(n3165), .Z(n3164) );
  BUFFD0 U3183 ( .I(n3166), .Z(n3165) );
  BUFFD0 U3184 ( .I(n3167), .Z(n3166) );
  BUFFD0 U3185 ( .I(n3168), .Z(n3167) );
  BUFFD0 U3186 ( .I(n3169), .Z(n3168) );
  BUFFD0 U3187 ( .I(n3170), .Z(n3169) );
  BUFFD0 U3188 ( .I(n3171), .Z(n3170) );
  BUFFD0 U3189 ( .I(n3172), .Z(n3171) );
  BUFFD0 U3190 ( .I(n3173), .Z(n3172) );
  BUFFD0 U3191 ( .I(n3174), .Z(n3173) );
  BUFFD0 U3192 ( .I(n3175), .Z(n3174) );
  BUFFD0 U3193 ( .I(n3176), .Z(n3175) );
  BUFFD0 U3194 ( .I(n3177), .Z(n3176) );
  BUFFD0 U3195 ( .I(n3178), .Z(n3177) );
  BUFFD0 U3196 ( .I(n3179), .Z(n3178) );
  BUFFD0 U3197 ( .I(n3180), .Z(n3179) );
  BUFFD0 U3198 ( .I(n3181), .Z(n3180) );
  BUFFD0 U3199 ( .I(n3182), .Z(n3181) );
  BUFFD0 U3200 ( .I(n3183), .Z(n3182) );
  BUFFD0 U3201 ( .I(n3184), .Z(n3183) );
  BUFFD0 U3202 ( .I(n3185), .Z(n3184) );
  BUFFD0 U3203 ( .I(n3186), .Z(n3185) );
  BUFFD0 U3204 ( .I(n3187), .Z(n3186) );
  BUFFD0 U3205 ( .I(n3188), .Z(n3187) );
  BUFFD0 U3206 ( .I(n3189), .Z(n3188) );
  BUFFD0 U3207 ( .I(n3190), .Z(n3189) );
  BUFFD0 U3208 ( .I(n3191), .Z(n3190) );
  BUFFD0 U3209 ( .I(n3192), .Z(n3191) );
  BUFFD0 U3210 ( .I(n3193), .Z(n3192) );
  BUFFD0 U3211 ( .I(n3194), .Z(n3193) );
  BUFFD0 U3212 ( .I(n3195), .Z(n3194) );
  BUFFD0 U3213 ( .I(n3196), .Z(n3195) );
  BUFFD0 U3214 ( .I(n3197), .Z(n3196) );
  BUFFD0 U3215 ( .I(n3198), .Z(n3197) );
  BUFFD0 U3216 ( .I(n3199), .Z(n3198) );
  BUFFD0 U3217 ( .I(n3200), .Z(n3199) );
  BUFFD0 U3218 ( .I(n3201), .Z(n3200) );
  BUFFD0 U3219 ( .I(n3202), .Z(n3201) );
  BUFFD0 U3220 ( .I(n3203), .Z(n3202) );
  BUFFD0 U3221 ( .I(n3204), .Z(n3203) );
  BUFFD0 U3222 ( .I(n3205), .Z(n3204) );
  BUFFD0 U3223 ( .I(n3206), .Z(n3205) );
  BUFFD0 U3224 ( .I(n3207), .Z(n3206) );
  BUFFD0 U3225 ( .I(n3208), .Z(n3207) );
  BUFFD0 U3226 ( .I(n3209), .Z(n3208) );
  BUFFD0 U3227 ( .I(n3210), .Z(n3209) );
  BUFFD0 U3228 ( .I(n3211), .Z(n3210) );
  BUFFD0 U3229 ( .I(n3212), .Z(n3211) );
  BUFFD0 U3230 ( .I(n3213), .Z(n3212) );
  BUFFD0 U3231 ( .I(n3214), .Z(n3213) );
  BUFFD0 U3232 ( .I(n3215), .Z(n3214) );
  BUFFD0 U3233 ( .I(n3216), .Z(n3215) );
  BUFFD0 U3234 ( .I(n3217), .Z(n3216) );
  BUFFD0 U3235 ( .I(n3218), .Z(n3217) );
  BUFFD0 U3236 ( .I(n3219), .Z(n3218) );
  BUFFD0 U3237 ( .I(n3220), .Z(n3219) );
  BUFFD0 U3238 ( .I(n3221), .Z(n3220) );
  BUFFD0 U3239 ( .I(n3222), .Z(n3221) );
  BUFFD0 U3240 ( .I(n3223), .Z(n3222) );
  BUFFD0 U3241 ( .I(n3224), .Z(n3223) );
  BUFFD0 U3242 ( .I(n3225), .Z(n3224) );
  BUFFD0 U3243 ( .I(N80), .Z(n3225) );
  CKBD0 U3244 ( .CLK(n3227), .C(n3291) );
  BUFFD0 U3245 ( .I(n3230), .Z(n3226) );
  BUFFD0 U3246 ( .I(N81), .Z(n3227) );
  BUFFD0 U3247 ( .I(n3502), .Z(n3228) );
  BUFFD0 U3248 ( .I(n3228), .Z(n3229) );
  BUFFD0 U3249 ( .I(n3231), .Z(n3230) );
  BUFFD0 U3250 ( .I(n3232), .Z(n3231) );
  BUFFD0 U3251 ( .I(n3233), .Z(n3232) );
  BUFFD0 U3252 ( .I(n3234), .Z(n3233) );
  BUFFD0 U3253 ( .I(n3235), .Z(n3234) );
  BUFFD0 U3254 ( .I(n3236), .Z(n3235) );
  BUFFD0 U3255 ( .I(n3237), .Z(n3236) );
  BUFFD0 U3256 ( .I(n3238), .Z(n3237) );
  BUFFD0 U3257 ( .I(n3239), .Z(n3238) );
  BUFFD0 U3258 ( .I(n3240), .Z(n3239) );
  BUFFD0 U3259 ( .I(n3241), .Z(n3240) );
  BUFFD0 U3260 ( .I(n3242), .Z(n3241) );
  BUFFD0 U3261 ( .I(n3243), .Z(n3242) );
  BUFFD0 U3262 ( .I(n3244), .Z(n3243) );
  BUFFD0 U3263 ( .I(n3245), .Z(n3244) );
  BUFFD0 U3264 ( .I(n3246), .Z(n3245) );
  BUFFD0 U3265 ( .I(n3247), .Z(n3246) );
  BUFFD0 U3266 ( .I(n3248), .Z(n3247) );
  BUFFD0 U3267 ( .I(n3249), .Z(n3248) );
  BUFFD0 U3268 ( .I(n3250), .Z(n3249) );
  BUFFD0 U3269 ( .I(n3251), .Z(n3250) );
  BUFFD0 U3270 ( .I(n3252), .Z(n3251) );
  BUFFD0 U3271 ( .I(n3253), .Z(n3252) );
  BUFFD0 U3272 ( .I(n3254), .Z(n3253) );
  BUFFD0 U3273 ( .I(n3255), .Z(n3254) );
  BUFFD0 U3274 ( .I(n3256), .Z(n3255) );
  BUFFD0 U3275 ( .I(n3257), .Z(n3256) );
  BUFFD0 U3276 ( .I(n3258), .Z(n3257) );
  BUFFD0 U3277 ( .I(n3259), .Z(n3258) );
  BUFFD0 U3278 ( .I(n3260), .Z(n3259) );
  BUFFD0 U3279 ( .I(n3261), .Z(n3260) );
  BUFFD0 U3280 ( .I(n3262), .Z(n3261) );
  BUFFD0 U3281 ( .I(n3263), .Z(n3262) );
  BUFFD0 U3282 ( .I(n3264), .Z(n3263) );
  BUFFD0 U3283 ( .I(n3265), .Z(n3264) );
  BUFFD0 U3284 ( .I(n3266), .Z(n3265) );
  BUFFD0 U3285 ( .I(n3267), .Z(n3266) );
  BUFFD0 U3286 ( .I(n3268), .Z(n3267) );
  BUFFD0 U3287 ( .I(n3269), .Z(n3268) );
  BUFFD0 U3288 ( .I(n3270), .Z(n3269) );
  BUFFD0 U3289 ( .I(n3271), .Z(n3270) );
  BUFFD0 U3290 ( .I(n3272), .Z(n3271) );
  BUFFD0 U3291 ( .I(n3273), .Z(n3272) );
  BUFFD0 U3292 ( .I(n3274), .Z(n3273) );
  BUFFD0 U3293 ( .I(n3275), .Z(n3274) );
  BUFFD0 U3294 ( .I(n3276), .Z(n3275) );
  BUFFD0 U3295 ( .I(n3277), .Z(n3276) );
  BUFFD0 U3296 ( .I(n3278), .Z(n3277) );
  BUFFD0 U3297 ( .I(n3279), .Z(n3278) );
  BUFFD0 U3298 ( .I(n3280), .Z(n3279) );
  BUFFD0 U3299 ( .I(n3281), .Z(n3280) );
  BUFFD0 U3300 ( .I(n3282), .Z(n3281) );
  BUFFD0 U3301 ( .I(n3283), .Z(n3282) );
  BUFFD0 U3302 ( .I(n3284), .Z(n3283) );
  BUFFD0 U3303 ( .I(n3285), .Z(n3284) );
  BUFFD0 U3304 ( .I(n3286), .Z(n3285) );
  BUFFD0 U3305 ( .I(n3287), .Z(n3286) );
  BUFFD0 U3306 ( .I(n3288), .Z(n3287) );
  BUFFD0 U3307 ( .I(n3289), .Z(n3288) );
  BUFFD0 U3308 ( .I(n3290), .Z(n3289) );
  BUFFD0 U3309 ( .I(n3292), .Z(n3290) );
  BUFFD0 U3310 ( .I(n3293), .Z(n3292) );
  BUFFD0 U3311 ( .I(n3229), .Z(n3293) );
  BUFFD0 U3312 ( .I(n3295), .Z(n3294) );
  BUFFD0 U3313 ( .I(n3296), .Z(n3295) );
  BUFFD0 U3314 ( .I(n3297), .Z(n3296) );
  BUFFD0 U3315 ( .I(n3298), .Z(n3297) );
  BUFFD0 U3316 ( .I(n3299), .Z(n3298) );
  BUFFD0 U3317 ( .I(n3300), .Z(n3299) );
  BUFFD0 U3318 ( .I(n3301), .Z(n3300) );
  BUFFD0 U3319 ( .I(n3302), .Z(n3301) );
  BUFFD0 U3320 ( .I(n3303), .Z(n3302) );
  BUFFD0 U3321 ( .I(n3304), .Z(n3303) );
  BUFFD0 U3322 ( .I(n3305), .Z(n3304) );
  BUFFD0 U3323 ( .I(n3306), .Z(n3305) );
  BUFFD0 U3324 ( .I(n3307), .Z(n3306) );
  BUFFD0 U3325 ( .I(n3308), .Z(n3307) );
  BUFFD0 U3326 ( .I(n3309), .Z(n3308) );
  BUFFD0 U3327 ( .I(n3310), .Z(n3309) );
  BUFFD0 U3328 ( .I(n3311), .Z(n3310) );
  BUFFD0 U3329 ( .I(n3312), .Z(n3311) );
  BUFFD0 U3330 ( .I(n3313), .Z(n3312) );
  BUFFD0 U3331 ( .I(n3314), .Z(n3313) );
  BUFFD0 U3332 ( .I(n3315), .Z(n3314) );
  BUFFD0 U3333 ( .I(n3316), .Z(n3315) );
  BUFFD0 U3334 ( .I(n3317), .Z(n3316) );
  BUFFD0 U3335 ( .I(n3318), .Z(n3317) );
  BUFFD0 U3336 ( .I(n3319), .Z(n3318) );
  BUFFD0 U3337 ( .I(n3320), .Z(n3319) );
  BUFFD0 U3338 ( .I(n3321), .Z(n3320) );
  BUFFD0 U3339 ( .I(n3322), .Z(n3321) );
  BUFFD0 U3340 ( .I(n3323), .Z(n3322) );
  BUFFD0 U3341 ( .I(n3324), .Z(n3323) );
  BUFFD0 U3342 ( .I(n3325), .Z(n3324) );
  BUFFD0 U3343 ( .I(n3326), .Z(n3325) );
  BUFFD0 U3344 ( .I(n3327), .Z(n3326) );
  BUFFD0 U3345 ( .I(n3328), .Z(n3327) );
  BUFFD0 U3346 ( .I(n3329), .Z(n3328) );
  BUFFD0 U3347 ( .I(n3330), .Z(n3329) );
  BUFFD0 U3348 ( .I(n3331), .Z(n3330) );
  BUFFD0 U3349 ( .I(n3332), .Z(n3331) );
  BUFFD0 U3350 ( .I(n3333), .Z(n3332) );
  BUFFD0 U3351 ( .I(n3334), .Z(n3333) );
  BUFFD0 U3352 ( .I(n3335), .Z(n3334) );
  BUFFD0 U3353 ( .I(n3336), .Z(n3335) );
  BUFFD0 U3354 ( .I(n3337), .Z(n3336) );
  BUFFD0 U3355 ( .I(n3338), .Z(n3337) );
  BUFFD0 U3356 ( .I(n3339), .Z(n3338) );
  BUFFD0 U3357 ( .I(n3340), .Z(n3339) );
  BUFFD0 U3358 ( .I(n3341), .Z(n3340) );
  BUFFD0 U3359 ( .I(n3342), .Z(n3341) );
  BUFFD0 U3360 ( .I(n3343), .Z(n3342) );
  BUFFD0 U3361 ( .I(n3344), .Z(n3343) );
  BUFFD0 U3362 ( .I(n3345), .Z(n3344) );
  BUFFD0 U3363 ( .I(n3346), .Z(n3345) );
  BUFFD0 U3364 ( .I(n3347), .Z(n3346) );
  BUFFD0 U3365 ( .I(n3348), .Z(n3347) );
  BUFFD0 U3366 ( .I(n3349), .Z(n3348) );
  BUFFD0 U3367 ( .I(n3350), .Z(n3349) );
  BUFFD0 U3368 ( .I(n3351), .Z(n3350) );
  BUFFD0 U3369 ( .I(n3352), .Z(n3351) );
  BUFFD0 U3370 ( .I(n3353), .Z(n3352) );
  BUFFD0 U3371 ( .I(n3354), .Z(n3353) );
  BUFFD0 U3372 ( .I(n3355), .Z(n3354) );
  BUFFD0 U3373 ( .I(n3356), .Z(n3355) );
  BUFFD0 U3374 ( .I(n3357), .Z(n3356) );
  BUFFD0 U3375 ( .I(n3358), .Z(n3357) );
  BUFFD0 U3376 ( .I(n3359), .Z(n3358) );
  BUFFD0 U3377 ( .I(n3360), .Z(n3359) );
  BUFFD0 U3378 ( .I(n3361), .Z(n3360) );
  BUFFD0 U3379 ( .I(n3362), .Z(n3361) );
  BUFFD0 U3380 ( .I(N82), .Z(n3362) );
  BUFFD0 U3381 ( .I(n3364), .Z(n3363) );
  BUFFD0 U3382 ( .I(n3365), .Z(n3364) );
  BUFFD0 U3383 ( .I(n3366), .Z(n3365) );
  BUFFD0 U3384 ( .I(n3367), .Z(n3366) );
  BUFFD0 U3385 ( .I(n3368), .Z(n3367) );
  BUFFD0 U3386 ( .I(n3369), .Z(n3368) );
  BUFFD0 U3387 ( .I(n3370), .Z(n3369) );
  BUFFD0 U3388 ( .I(n3371), .Z(n3370) );
  BUFFD0 U3389 ( .I(n3372), .Z(n3371) );
  BUFFD0 U3390 ( .I(n3373), .Z(n3372) );
  BUFFD0 U3391 ( .I(n3374), .Z(n3373) );
  BUFFD0 U3392 ( .I(n3375), .Z(n3374) );
  BUFFD0 U3393 ( .I(n3376), .Z(n3375) );
  BUFFD0 U3394 ( .I(n3377), .Z(n3376) );
  BUFFD0 U3395 ( .I(n3378), .Z(n3377) );
  BUFFD0 U3396 ( .I(n3379), .Z(n3378) );
  BUFFD0 U3397 ( .I(n3380), .Z(n3379) );
  BUFFD0 U3398 ( .I(n3381), .Z(n3380) );
  BUFFD0 U3399 ( .I(n3382), .Z(n3381) );
  BUFFD0 U3400 ( .I(n3383), .Z(n3382) );
  BUFFD0 U3401 ( .I(n3384), .Z(n3383) );
  BUFFD0 U3402 ( .I(n3385), .Z(n3384) );
  BUFFD0 U3403 ( .I(n3386), .Z(n3385) );
  BUFFD0 U3404 ( .I(n3387), .Z(n3386) );
  BUFFD0 U3405 ( .I(n3388), .Z(n3387) );
  BUFFD0 U3406 ( .I(n3389), .Z(n3388) );
  BUFFD0 U3407 ( .I(n3390), .Z(n3389) );
  BUFFD0 U3408 ( .I(n3391), .Z(n3390) );
  BUFFD0 U3409 ( .I(n3392), .Z(n3391) );
  BUFFD0 U3410 ( .I(n3393), .Z(n3392) );
  BUFFD0 U3411 ( .I(n3394), .Z(n3393) );
  BUFFD0 U3412 ( .I(n3395), .Z(n3394) );
  BUFFD0 U3413 ( .I(n3396), .Z(n3395) );
  BUFFD0 U3414 ( .I(n3397), .Z(n3396) );
  BUFFD0 U3415 ( .I(n3398), .Z(n3397) );
  BUFFD0 U3416 ( .I(n3399), .Z(n3398) );
  BUFFD0 U3417 ( .I(n3400), .Z(n3399) );
  BUFFD0 U3418 ( .I(n3401), .Z(n3400) );
  BUFFD0 U3419 ( .I(n3402), .Z(n3401) );
  BUFFD0 U3420 ( .I(n3403), .Z(n3402) );
  BUFFD0 U3421 ( .I(n3404), .Z(n3403) );
  BUFFD0 U3422 ( .I(n3405), .Z(n3404) );
  BUFFD0 U3423 ( .I(n3406), .Z(n3405) );
  BUFFD0 U3424 ( .I(n3407), .Z(n3406) );
  BUFFD0 U3425 ( .I(n3408), .Z(n3407) );
  BUFFD0 U3426 ( .I(n3409), .Z(n3408) );
  BUFFD0 U3427 ( .I(n3410), .Z(n3409) );
  BUFFD0 U3428 ( .I(n3411), .Z(n3410) );
  BUFFD0 U3429 ( .I(n3412), .Z(n3411) );
  BUFFD0 U3430 ( .I(n3413), .Z(n3412) );
  BUFFD0 U3431 ( .I(n3414), .Z(n3413) );
  BUFFD0 U3432 ( .I(n3415), .Z(n3414) );
  BUFFD0 U3433 ( .I(n3416), .Z(n3415) );
  BUFFD0 U3434 ( .I(n3417), .Z(n3416) );
  BUFFD0 U3435 ( .I(n3418), .Z(n3417) );
  BUFFD0 U3436 ( .I(n3419), .Z(n3418) );
  BUFFD0 U3437 ( .I(n3420), .Z(n3419) );
  BUFFD0 U3438 ( .I(n3421), .Z(n3420) );
  BUFFD0 U3439 ( .I(n3422), .Z(n3421) );
  BUFFD0 U3440 ( .I(n3423), .Z(n3422) );
  BUFFD0 U3441 ( .I(n3424), .Z(n3423) );
  BUFFD0 U3442 ( .I(n3425), .Z(n3424) );
  BUFFD0 U3443 ( .I(n3426), .Z(n3425) );
  BUFFD0 U3444 ( .I(n3427), .Z(n3426) );
  BUFFD0 U3445 ( .I(n3428), .Z(n3427) );
  BUFFD0 U3446 ( .I(n3429), .Z(n3428) );
  BUFFD0 U3447 ( .I(n3430), .Z(n3429) );
  BUFFD0 U3448 ( .I(n3431), .Z(n3430) );
  BUFFD0 U3449 ( .I(N83), .Z(n3431) );
  BUFFD0 U3450 ( .I(n3433), .Z(n3432) );
  BUFFD0 U3451 ( .I(n3434), .Z(n3433) );
  BUFFD0 U3452 ( .I(n3435), .Z(n3434) );
  BUFFD0 U3453 ( .I(n3436), .Z(n3435) );
  BUFFD0 U3454 ( .I(n3437), .Z(n3436) );
  BUFFD0 U3455 ( .I(n3438), .Z(n3437) );
  BUFFD0 U3456 ( .I(n3439), .Z(n3438) );
  BUFFD0 U3457 ( .I(n3440), .Z(n3439) );
  BUFFD0 U3458 ( .I(n3441), .Z(n3440) );
  BUFFD0 U3459 ( .I(n3442), .Z(n3441) );
  BUFFD0 U3460 ( .I(n3443), .Z(n3442) );
  BUFFD0 U3461 ( .I(n3444), .Z(n3443) );
  BUFFD0 U3462 ( .I(n3445), .Z(n3444) );
  BUFFD0 U3463 ( .I(n3446), .Z(n3445) );
  BUFFD0 U3464 ( .I(n3447), .Z(n3446) );
  BUFFD0 U3465 ( .I(n3448), .Z(n3447) );
  BUFFD0 U3466 ( .I(n3449), .Z(n3448) );
  BUFFD0 U3467 ( .I(n3450), .Z(n3449) );
  BUFFD0 U3468 ( .I(n3451), .Z(n3450) );
  BUFFD0 U3469 ( .I(n3452), .Z(n3451) );
  BUFFD0 U3470 ( .I(n3453), .Z(n3452) );
  BUFFD0 U3471 ( .I(n3454), .Z(n3453) );
  BUFFD0 U3472 ( .I(n3455), .Z(n3454) );
  BUFFD0 U3473 ( .I(n3456), .Z(n3455) );
  BUFFD0 U3474 ( .I(n3457), .Z(n3456) );
  BUFFD0 U3475 ( .I(n3458), .Z(n3457) );
  BUFFD0 U3476 ( .I(n3459), .Z(n3458) );
  BUFFD0 U3477 ( .I(n3460), .Z(n3459) );
  BUFFD0 U3478 ( .I(n3461), .Z(n3460) );
  BUFFD0 U3479 ( .I(n3462), .Z(n3461) );
  BUFFD0 U3480 ( .I(n3463), .Z(n3462) );
  BUFFD0 U3481 ( .I(n3464), .Z(n3463) );
  BUFFD0 U3482 ( .I(n3465), .Z(n3464) );
  BUFFD0 U3483 ( .I(n3466), .Z(n3465) );
  BUFFD0 U3484 ( .I(n3467), .Z(n3466) );
  BUFFD0 U3485 ( .I(n3468), .Z(n3467) );
  BUFFD0 U3486 ( .I(n3469), .Z(n3468) );
  BUFFD0 U3487 ( .I(n3470), .Z(n3469) );
  BUFFD0 U3488 ( .I(n3471), .Z(n3470) );
  BUFFD0 U3489 ( .I(n3472), .Z(n3471) );
  BUFFD0 U3490 ( .I(n3473), .Z(n3472) );
  BUFFD0 U3491 ( .I(n3474), .Z(n3473) );
  BUFFD0 U3492 ( .I(n3475), .Z(n3474) );
  BUFFD0 U3493 ( .I(n3476), .Z(n3475) );
  BUFFD0 U3494 ( .I(n3477), .Z(n3476) );
  BUFFD0 U3495 ( .I(n3478), .Z(n3477) );
  BUFFD0 U3496 ( .I(n3479), .Z(n3478) );
  BUFFD0 U3497 ( .I(n3480), .Z(n3479) );
  BUFFD0 U3498 ( .I(n3481), .Z(n3480) );
  BUFFD0 U3499 ( .I(n3482), .Z(n3481) );
  BUFFD0 U3500 ( .I(n3483), .Z(n3482) );
  BUFFD0 U3501 ( .I(n3484), .Z(n3483) );
  BUFFD0 U3502 ( .I(n3485), .Z(n3484) );
  BUFFD0 U3503 ( .I(n3486), .Z(n3485) );
  BUFFD0 U3504 ( .I(n3487), .Z(n3486) );
  BUFFD0 U3505 ( .I(n3488), .Z(n3487) );
  BUFFD0 U3506 ( .I(n3489), .Z(n3488) );
  BUFFD0 U3507 ( .I(n3490), .Z(n3489) );
  BUFFD0 U3508 ( .I(n3491), .Z(n3490) );
  BUFFD0 U3509 ( .I(n3492), .Z(n3491) );
  BUFFD0 U3510 ( .I(n3493), .Z(n3492) );
  BUFFD0 U3511 ( .I(n3494), .Z(n3493) );
  BUFFD0 U3512 ( .I(n3495), .Z(n3494) );
  BUFFD0 U3513 ( .I(n3496), .Z(n3495) );
  BUFFD0 U3514 ( .I(n3497), .Z(n3496) );
  BUFFD0 U3515 ( .I(n3498), .Z(n3497) );
  BUFFD0 U3516 ( .I(n3499), .Z(n3498) );
  BUFFD0 U3517 ( .I(n3500), .Z(n3499) );
  BUFFD0 U3518 ( .I(N84), .Z(n3500) );
  BUFFD0 U3519 ( .I(n2944), .Z(n3501) );
  BUFFD0 U3520 ( .I(n3291), .Z(n3502) );
  BUFFD0 U3521 ( .I(n3504), .Z(n3503) );
  BUFFD0 U3522 ( .I(n3505), .Z(n3504) );
  BUFFD0 U3523 ( .I(n3506), .Z(n3505) );
  BUFFD0 U3524 ( .I(n3507), .Z(n3506) );
  BUFFD0 U3525 ( .I(n3508), .Z(n3507) );
  BUFFD0 U3526 ( .I(n3509), .Z(n3508) );
  BUFFD0 U3527 ( .I(n3510), .Z(n3509) );
  BUFFD0 U3528 ( .I(n3511), .Z(n3510) );
  BUFFD0 U3529 ( .I(n3512), .Z(n3511) );
  BUFFD0 U3530 ( .I(n3513), .Z(n3512) );
  BUFFD0 U3531 ( .I(n3514), .Z(n3513) );
  BUFFD0 U3532 ( .I(n3515), .Z(n3514) );
  BUFFD0 U3533 ( .I(n3516), .Z(n3515) );
  BUFFD0 U3534 ( .I(n3517), .Z(n3516) );
  BUFFD0 U3535 ( .I(n3518), .Z(n3517) );
  BUFFD0 U3536 ( .I(n3519), .Z(n3518) );
  BUFFD0 U3537 ( .I(n3520), .Z(n3519) );
  BUFFD0 U3538 ( .I(n3521), .Z(n3520) );
  BUFFD0 U3539 ( .I(n3522), .Z(n3521) );
  BUFFD0 U3540 ( .I(n3523), .Z(n3522) );
  BUFFD0 U3541 ( .I(n3524), .Z(n3523) );
  BUFFD0 U3542 ( .I(n3525), .Z(n3524) );
  BUFFD0 U3543 ( .I(n3526), .Z(n3525) );
  BUFFD0 U3544 ( .I(n3527), .Z(n3526) );
  BUFFD0 U3545 ( .I(n3528), .Z(n3527) );
  BUFFD0 U3546 ( .I(n3529), .Z(n3528) );
  BUFFD0 U3547 ( .I(n3530), .Z(n3529) );
  BUFFD0 U3548 ( .I(n3531), .Z(n3530) );
  BUFFD0 U3549 ( .I(n3532), .Z(n3531) );
  BUFFD0 U3550 ( .I(n3533), .Z(n3532) );
  BUFFD0 U3551 ( .I(n3534), .Z(n3533) );
  BUFFD0 U3552 ( .I(n3535), .Z(n3534) );
  BUFFD0 U3553 ( .I(n3536), .Z(n3535) );
  BUFFD0 U3554 ( .I(n3537), .Z(n3536) );
  BUFFD0 U3555 ( .I(n3538), .Z(n3537) );
  BUFFD0 U3556 ( .I(n3539), .Z(n3538) );
  BUFFD0 U3557 ( .I(n3540), .Z(n3539) );
  BUFFD0 U3558 ( .I(n3541), .Z(n3540) );
  BUFFD0 U3559 ( .I(n3542), .Z(n3541) );
  BUFFD0 U3560 ( .I(n3543), .Z(n3542) );
  BUFFD0 U3561 ( .I(n3544), .Z(n3543) );
  BUFFD0 U3562 ( .I(n3545), .Z(n3544) );
  BUFFD0 U3563 ( .I(n3546), .Z(n3545) );
  BUFFD0 U3564 ( .I(n3547), .Z(n3546) );
  BUFFD0 U3565 ( .I(n3548), .Z(n3547) );
  BUFFD0 U3566 ( .I(n3549), .Z(n3548) );
  BUFFD0 U3567 ( .I(n3550), .Z(n3549) );
  BUFFD0 U3568 ( .I(n3551), .Z(n3550) );
  BUFFD0 U3569 ( .I(n3552), .Z(n3551) );
  BUFFD0 U3570 ( .I(n3553), .Z(n3552) );
  BUFFD0 U3571 ( .I(n3554), .Z(n3553) );
  BUFFD0 U3572 ( .I(n3555), .Z(n3554) );
  BUFFD0 U3573 ( .I(n3556), .Z(n3555) );
  BUFFD0 U3574 ( .I(n3557), .Z(n3556) );
  BUFFD0 U3575 ( .I(n3558), .Z(n3557) );
  BUFFD0 U3576 ( .I(n3559), .Z(n3558) );
  BUFFD0 U3577 ( .I(n3560), .Z(n3559) );
  BUFFD0 U3578 ( .I(n3561), .Z(n3560) );
  BUFFD0 U3579 ( .I(n3562), .Z(n3561) );
  BUFFD0 U3580 ( .I(n3563), .Z(n3562) );
  BUFFD0 U3581 ( .I(n3564), .Z(n3563) );
  BUFFD0 U3582 ( .I(n3565), .Z(n3564) );
  BUFFD0 U3583 ( .I(n3566), .Z(n3565) );
  BUFFD0 U3584 ( .I(n3567), .Z(n3566) );
  BUFFD0 U3585 ( .I(n3568), .Z(n3567) );
  BUFFD0 U3586 ( .I(N85), .Z(n3568) );
  BUFFD0 U3587 ( .I(n3570), .Z(n3569) );
  BUFFD0 U3588 ( .I(n3571), .Z(n3570) );
  BUFFD0 U3589 ( .I(n3572), .Z(n3571) );
  BUFFD0 U3590 ( .I(n3573), .Z(n3572) );
  BUFFD0 U3591 ( .I(n3574), .Z(n3573) );
  BUFFD0 U3592 ( .I(n3575), .Z(n3574) );
  BUFFD0 U3593 ( .I(n3576), .Z(n3575) );
  BUFFD0 U3594 ( .I(n3577), .Z(n3576) );
  BUFFD0 U3595 ( .I(n3578), .Z(n3577) );
  BUFFD0 U3596 ( .I(n3579), .Z(n3578) );
  BUFFD0 U3597 ( .I(n3580), .Z(n3579) );
  BUFFD0 U3598 ( .I(n3581), .Z(n3580) );
  BUFFD0 U3599 ( .I(n3582), .Z(n3581) );
  BUFFD0 U3600 ( .I(n3583), .Z(n3582) );
  BUFFD0 U3601 ( .I(n3584), .Z(n3583) );
  BUFFD0 U3602 ( .I(n3585), .Z(n3584) );
  BUFFD0 U3603 ( .I(n3586), .Z(n3585) );
  BUFFD0 U3604 ( .I(n3587), .Z(n3586) );
  BUFFD0 U3605 ( .I(n3588), .Z(n3587) );
  BUFFD0 U3606 ( .I(n3589), .Z(n3588) );
  BUFFD0 U3607 ( .I(n3590), .Z(n3589) );
  BUFFD0 U3608 ( .I(n3591), .Z(n3590) );
  BUFFD0 U3609 ( .I(n3592), .Z(n3591) );
  BUFFD0 U3610 ( .I(n3593), .Z(n3592) );
  BUFFD0 U3611 ( .I(n3594), .Z(n3593) );
  BUFFD0 U3612 ( .I(n3595), .Z(n3594) );
  BUFFD0 U3613 ( .I(n3596), .Z(n3595) );
  BUFFD0 U3614 ( .I(n3597), .Z(n3596) );
  BUFFD0 U3615 ( .I(n3598), .Z(n3597) );
  BUFFD0 U3616 ( .I(n3599), .Z(n3598) );
  BUFFD0 U3617 ( .I(n3600), .Z(n3599) );
  BUFFD0 U3618 ( .I(n3601), .Z(n3600) );
  BUFFD0 U3619 ( .I(n3602), .Z(n3601) );
  BUFFD0 U3620 ( .I(n3603), .Z(n3602) );
  BUFFD0 U3621 ( .I(n3604), .Z(n3603) );
  BUFFD0 U3622 ( .I(n3605), .Z(n3604) );
  BUFFD0 U3623 ( .I(n3606), .Z(n3605) );
  BUFFD0 U3624 ( .I(n3607), .Z(n3606) );
  BUFFD0 U3625 ( .I(n3608), .Z(n3607) );
  BUFFD0 U3626 ( .I(n3609), .Z(n3608) );
  BUFFD0 U3627 ( .I(n3610), .Z(n3609) );
  BUFFD0 U3628 ( .I(n3611), .Z(n3610) );
  BUFFD0 U3629 ( .I(n3612), .Z(n3611) );
  BUFFD0 U3630 ( .I(n3613), .Z(n3612) );
  BUFFD0 U3631 ( .I(n3614), .Z(n3613) );
  BUFFD0 U3632 ( .I(n3615), .Z(n3614) );
  BUFFD0 U3633 ( .I(n3616), .Z(n3615) );
  BUFFD0 U3634 ( .I(n3817), .Z(n3616) );
  CKAN2D0 U3635 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U3636 ( .I(N50), .ZN(n3717) );
  BUFFD1 U3637 ( .I(n3848), .Z(n3826) );
  BUFFD1 U3638 ( .I(n3848), .Z(n3827) );
  BUFFD1 U3639 ( .I(n3845), .Z(n3828) );
  BUFFD1 U3640 ( .I(n3845), .Z(n3829) );
  BUFFD1 U3641 ( .I(n3845), .Z(n3830) );
  BUFFD1 U3642 ( .I(n3850), .Z(n3831) );
  BUFFD1 U3643 ( .I(n3848), .Z(n3832) );
  BUFFD1 U3644 ( .I(n3848), .Z(n3833) );
  BUFFD1 U3645 ( .I(n3848), .Z(n3834) );
  BUFFD1 U3646 ( .I(n3850), .Z(n3835) );
  BUFFD1 U3647 ( .I(n3847), .Z(n3836) );
  BUFFD1 U3648 ( .I(n3847), .Z(n3837) );
  BUFFD1 U3649 ( .I(n3847), .Z(n3838) );
  BUFFD1 U3650 ( .I(n3847), .Z(n3839) );
  BUFFD1 U3651 ( .I(n3846), .Z(n3840) );
  BUFFD1 U3652 ( .I(n3846), .Z(n3841) );
  BUFFD1 U3653 ( .I(n3845), .Z(n3842) );
  BUFFD1 U3654 ( .I(n3845), .Z(n3843) );
  BUFFD1 U3655 ( .I(n3848), .Z(n3844) );
  BUFFD1 U3656 ( .I(n3850), .Z(n3820) );
  BUFFD1 U3657 ( .I(n3850), .Z(n3821) );
  BUFFD1 U3658 ( .I(n3849), .Z(n3822) );
  BUFFD1 U3659 ( .I(n3849), .Z(n3823) );
  BUFFD1 U3660 ( .I(n3850), .Z(n3824) );
  BUFFD1 U3661 ( .I(n3849), .Z(n3825) );
  BUFFD1 U3662 ( .I(n3853), .Z(n3848) );
  BUFFD1 U3663 ( .I(n3852), .Z(n3847) );
  BUFFD1 U3664 ( .I(n3852), .Z(n3846) );
  BUFFD1 U3665 ( .I(n3852), .Z(n3845) );
  BUFFD1 U3666 ( .I(n3851), .Z(n3849) );
  BUFFD1 U3667 ( .I(n3851), .Z(n3850) );
  BUFFD1 U3668 ( .I(n3854), .Z(n3852) );
  BUFFD1 U3669 ( .I(n3854), .Z(n3853) );
  BUFFD1 U3670 ( .I(n3854), .Z(n3851) );
  INVD1 U3671 ( .I(Reset), .ZN(n3854) );
  BUFFD1 U3672 ( .I(n3809), .Z(n3797) );
  BUFFD1 U3673 ( .I(n3804), .Z(n3796) );
  BUFFD1 U3674 ( .I(n3804), .Z(n3795) );
  BUFFD1 U3675 ( .I(n3805), .Z(n3794) );
  BUFFD1 U3676 ( .I(n3805), .Z(n3793) );
  BUFFD1 U3677 ( .I(n3806), .Z(n3792) );
  BUFFD1 U3678 ( .I(n3806), .Z(n3791) );
  BUFFD1 U3679 ( .I(n3807), .Z(n3790) );
  BUFFD1 U3680 ( .I(n3807), .Z(n3789) );
  BUFFD1 U3681 ( .I(n3808), .Z(n3788) );
  BUFFD1 U3682 ( .I(n3808), .Z(n3787) );
  BUFFD1 U3683 ( .I(n3809), .Z(n3786) );
  BUFFD1 U3684 ( .I(n3809), .Z(n3785) );
  BUFFD1 U3685 ( .I(n3810), .Z(n3784) );
  BUFFD1 U3686 ( .I(n3810), .Z(n3783) );
  BUFFD1 U3687 ( .I(n3811), .Z(n3782) );
  BUFFD1 U3688 ( .I(n3811), .Z(n3781) );
  BUFFD1 U3689 ( .I(n3812), .Z(n3780) );
  BUFFD1 U3690 ( .I(n3812), .Z(n3779) );
  INVD1 U3691 ( .I(n3765), .ZN(n3766) );
  INVD1 U3692 ( .I(n6), .ZN(n3762) );
  INVD1 U3693 ( .I(n3756), .ZN(n3754) );
  INVD1 U3694 ( .I(n6), .ZN(n3763) );
  INVD1 U3695 ( .I(n3756), .ZN(n3755) );
  INVD1 U3696 ( .I(n7), .ZN(n3753) );
  BUFFD1 U3697 ( .I(n3802), .Z(n3800) );
  BUFFD1 U3698 ( .I(n3803), .Z(n3799) );
  BUFFD1 U3699 ( .I(n3803), .Z(n3798) );
  BUFFD1 U3700 ( .I(n3774), .Z(n3804) );
  BUFFD1 U3701 ( .I(n3774), .Z(n3805) );
  BUFFD1 U3702 ( .I(n3774), .Z(n3806) );
  BUFFD1 U3703 ( .I(n3775), .Z(n3807) );
  BUFFD1 U3704 ( .I(n3775), .Z(n3808) );
  BUFFD1 U3705 ( .I(n3775), .Z(n3809) );
  BUFFD1 U3706 ( .I(n3776), .Z(n3810) );
  BUFFD1 U3707 ( .I(n3776), .Z(n3811) );
  BUFFD1 U3708 ( .I(n3776), .Z(n3812) );
  BUFFD1 U3709 ( .I(n3802), .Z(n3801) );
  INVD1 U3710 ( .I(N326), .ZN(n3756) );
  INVD1 U3711 ( .I(n3772), .ZN(n3771) );
  INVD1 U3712 ( .I(n3772), .ZN(n3770) );
  INVD1 U3713 ( .I(n4), .ZN(n3767) );
  INVD1 U3714 ( .I(n3), .ZN(n3761) );
  INVD1 U3715 ( .I(n3), .ZN(n3760) );
  INVD1 U3716 ( .I(n3759), .ZN(n3757) );
  INVD1 U3717 ( .I(n4), .ZN(n3768) );
  INVD1 U3718 ( .I(n3759), .ZN(n3758) );
  BUFFD1 U3719 ( .I(n3773), .Z(n3802) );
  BUFFD1 U3720 ( .I(n3773), .Z(n3803) );
  BUFFD1 U3721 ( .I(n3812), .Z(n3774) );
  BUFFD1 U3722 ( .I(n3777), .Z(n3775) );
  BUFFD1 U3723 ( .I(n3777), .Z(n3776) );
  INVD1 U3724 ( .I(n5), .ZN(n3814) );
  INVD1 U3725 ( .I(n5), .ZN(n3813) );
  XOR3D1 U3726 ( .A1(n77), .A2(n3738), .A3(n78), .Z(n76) );
  XOR3D1 U3727 ( .A1(n71), .A2(n3729), .A3(n72), .Z(n70) );
  XOR3D1 U3728 ( .A1(DataI[12]), .A2(n3735), .A3(n73), .Z(n72) );
  XOR3D1 U3729 ( .A1(n74), .A2(n3734), .A3(n75), .Z(n73) );
  XOR3D1 U3730 ( .A1(DataI[5]), .A2(n914), .A3(n70), .Z(n69) );
  XOR3D1 U3731 ( .A1(N69), .A2(N68), .A3(n85), .Z(n83) );
  XOR3D1 U3732 ( .A1(N67), .A2(n86), .A3(n87), .Z(n85) );
  BUFFD1 U3733 ( .I(n3722), .Z(n3725) );
  BUFFD1 U3734 ( .I(n3818), .Z(n3722) );
  XOR3D1 U3735 ( .A1(N62), .A2(N61), .A3(n88), .Z(n87) );
  XOR3D1 U3736 ( .A1(n89), .A2(N60), .A3(n90), .Z(n88) );
  XOR3D1 U3737 ( .A1(n3502), .A2(n3501), .A3(n79), .Z(N85) );
  XOR3D1 U3738 ( .A1(N75), .A2(n80), .A3(n81), .Z(n79) );
  XOR3D1 U3739 ( .A1(N79), .A2(N78), .A3(n82), .Z(n81) );
  BUFFD1 U3740 ( .I(n3818), .Z(n3723) );
  BUFFD1 U3741 ( .I(n3819), .Z(n3721) );
  BUFFD1 U3742 ( .I(n3818), .Z(n3724) );
  BUFFD1 U3743 ( .I(n3819), .Z(n3720) );
  INVD1 U3744 ( .I(n3717), .ZN(n3718) );
  INVD1 U3745 ( .I(n3717), .ZN(n3719) );
  INVD1 U3746 ( .I(AddrW[0]), .ZN(n93) );
  INVD1 U3747 ( .I(n3769), .ZN(n3772) );
  INVD1 U3748 ( .I(N293), .ZN(n3759) );
  INVD1 U3749 ( .I(N194), .ZN(n3765) );
  NR3D0 U3750 ( .A1(n91), .A2(AddrW[0]), .A3(n10), .ZN(N194) );
  NR3D0 U3751 ( .A1(n91), .A2(AddrW[0]), .A3(n1267), .ZN(N326) );
  INVD1 U3752 ( .I(n7), .ZN(n3752) );
  INVD1 U3753 ( .I(n2), .ZN(n3815) );
  INVD1 U3754 ( .I(n2), .ZN(n3816) );
  BUFFD1 U3755 ( .I(ClockW), .Z(n3777) );
  BUFFD1 U3756 ( .I(n3778), .Z(n3773) );
  BUFFD1 U3757 ( .I(ClockW), .Z(n3778) );
  MUX4ND0 U3758 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n3725), .S1(N49), .ZN(
        n3623) );
  MUX4ND0 U3759 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n3725), .S1(N49), .ZN(
        n3626) );
  MUX4ND0 U3760 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n3725), .S1(n3720), .ZN(
        n3641) );
  MUX4ND0 U3761 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n3818), .S1(n3720), .ZN(
        n3656) );
  MUX4ND0 U3762 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(N48), .S1(n3720), .ZN(
        n3659) );
  MUX4ND0 U3763 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n3722), .S1(n3720), .ZN(
        n3677) );
  MUX4ND0 U3764 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n3723), .S1(n3721), .ZN(
        n3680) );
  MUX4ND0 U3765 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n3723), .S1(n3720), .ZN(
        n3698) );
  MUX4ND0 U3766 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n3725), .S1(n3720), .ZN(
        n3701) );
  MUX4ND0 U3767 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n3725), .S1(n3720), .ZN(
        n3710) );
  MUX4ND0 U3768 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n3725), .S1(n3720), .ZN(
        n3713) );
  MUX4ND0 U3769 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n3818), .S1(n3720), .ZN(
        n3638) );
  MUX4ND0 U3770 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n3818), .S1(N49), .ZN(
        n3644) );
  MUX4ND0 U3771 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n3818), .S1(n3720), .ZN(
        n3668) );
  MUX4ND0 U3772 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(N48), .S1(n3721), .ZN(
        n3689) );
  MUX4ND0 U3773 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n3725), .S1(n3720), .ZN(
        n3692) );
  MUX4ND0 U3774 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n3725), .S1(N49), .ZN(
        n3620) );
  MUX4ND0 U3775 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(N48), .S1(N49), .ZN(n3632)
         );
  MUX4ND0 U3776 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n3818), .S1(n3819), .ZN(
        n3650) );
  MUX4ND0 U3777 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(N48), .S1(n3720), .ZN(
        n3653) );
  MUX4ND0 U3778 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n3818), .S1(n3720), .ZN(
        n3662) );
  MUX4ND0 U3779 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(N48), .S1(n3720), .ZN(
        n3674) );
  MUX4ND0 U3780 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n3818), .S1(N49), .ZN(
        n3683) );
  MUX4ND0 U3781 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n3723), .S1(n3720), .ZN(
        n3695) );
  MUX4ND0 U3782 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n3725), .S1(n3720), .ZN(
        n3704) );
  MUX4ND0 U3783 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n3725), .S1(n3721), .ZN(
        n3707) );
  MUX4ND0 U3784 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n3725), .S1(N49), .ZN(
        n3629) );
  MUX4ND0 U3785 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(N48), .S1(N49), .ZN(n3635)
         );
  MUX4ND0 U3786 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n3818), .S1(n3819), .ZN(
        n3647) );
  MUX4ND0 U3787 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n3818), .S1(n3720), .ZN(
        n3665) );
  MUX4ND0 U3788 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(N48), .S1(n3720), .ZN(
        n3671) );
  MUX4ND0 U3789 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n3722), .S1(n3819), .ZN(
        n3686) );
  MUX4ND0 U3790 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n3725), .S1(n3720), .ZN(
        n3716) );
  BUFFD1 U3791 ( .I(N48), .Z(n3818) );
  BUFFD1 U3792 ( .I(N49), .Z(n3819) );
  INVD1 U3793 ( .I(AddrW[1]), .ZN(n91) );
  ND2D1 U3794 ( .A1(AddrW[2]), .A2(Write), .ZN(n92) );
  NR3D0 U3795 ( .A1(n93), .A2(AddrW[1]), .A3(n1267), .ZN(N293) );
  INVD1 U3796 ( .I(Read), .ZN(n3817) );
  CKAN2D0 U3797 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  MUX3ND0 U3798 ( .I0(n3618), .I1(n3619), .I2(n3620), .S0(n3721), .S1(n3718), 
        .ZN(N84) );
  MUX3ND0 U3799 ( .I0(n3621), .I1(n3622), .I2(n3623), .S0(n3721), .S1(n3718), 
        .ZN(N83) );
  MUX3ND0 U3800 ( .I0(n3624), .I1(n3625), .I2(n3626), .S0(n3721), .S1(n3718), 
        .ZN(N82) );
  MUX3ND0 U3801 ( .I0(n3627), .I1(n3628), .I2(n3629), .S0(n3721), .S1(n3718), 
        .ZN(N81) );
  MUX3ND0 U3802 ( .I0(n3630), .I1(n3631), .I2(n3632), .S0(n3721), .S1(n3718), 
        .ZN(N80) );
  MUX3ND0 U3803 ( .I0(n3633), .I1(n3634), .I2(n3635), .S0(n3721), .S1(n3718), 
        .ZN(N79) );
  MUX3ND0 U3804 ( .I0(n3636), .I1(n3637), .I2(n3638), .S0(n3721), .S1(n3718), 
        .ZN(N78) );
  MUX3ND0 U3805 ( .I0(n3639), .I1(n3640), .I2(n3641), .S0(n3721), .S1(n3718), 
        .ZN(N77) );
  MUX3ND0 U3806 ( .I0(n3642), .I1(n3643), .I2(n3644), .S0(n3721), .S1(n3718), 
        .ZN(N76) );
  MUX3ND0 U3807 ( .I0(n3645), .I1(n3646), .I2(n3647), .S0(n3721), .S1(n3718), 
        .ZN(N75) );
  MUX3ND0 U3808 ( .I0(n3648), .I1(n3649), .I2(n3650), .S0(n3721), .S1(n3718), 
        .ZN(N74) );
  MUX3ND0 U3809 ( .I0(n3651), .I1(n3652), .I2(n3653), .S0(n3721), .S1(n3718), 
        .ZN(N73) );
  MUX3ND0 U3810 ( .I0(n3654), .I1(n3655), .I2(n3656), .S0(n3721), .S1(n3718), 
        .ZN(N72) );
  MUX3ND0 U3811 ( .I0(n3657), .I1(n3658), .I2(n3659), .S0(n3819), .S1(n3718), 
        .ZN(N71) );
  MUX3ND0 U3812 ( .I0(n3660), .I1(n3661), .I2(n3662), .S0(n3819), .S1(n3718), 
        .ZN(N70) );
  MUX3ND0 U3813 ( .I0(n3663), .I1(n3664), .I2(n3665), .S0(n3819), .S1(n3718), 
        .ZN(N69) );
  MUX3ND0 U3814 ( .I0(n3666), .I1(n3667), .I2(n3668), .S0(n3819), .S1(n3718), 
        .ZN(N68) );
  MUX3ND0 U3815 ( .I0(n3669), .I1(n3670), .I2(n3671), .S0(n3819), .S1(n3718), 
        .ZN(N67) );
  MUX3ND0 U3816 ( .I0(n3672), .I1(n3673), .I2(n3674), .S0(n3819), .S1(n3718), 
        .ZN(N66) );
  MUX3ND0 U3817 ( .I0(n3675), .I1(n3676), .I2(n3677), .S0(n3819), .S1(n3718), 
        .ZN(N65) );
  MUX3ND0 U3818 ( .I0(n3678), .I1(n3679), .I2(n3680), .S0(n3819), .S1(n3719), 
        .ZN(N64) );
  MUX3ND0 U3819 ( .I0(n3681), .I1(n3682), .I2(n3683), .S0(n3819), .S1(n3719), 
        .ZN(N63) );
  MUX3ND0 U3820 ( .I0(n3684), .I1(n3685), .I2(n3686), .S0(n3819), .S1(n3719), 
        .ZN(N62) );
  MUX3ND0 U3821 ( .I0(n3687), .I1(n3688), .I2(n3689), .S0(n3819), .S1(n3719), 
        .ZN(N61) );
  MUX3ND0 U3822 ( .I0(n3690), .I1(n3691), .I2(n3692), .S0(n3819), .S1(n3719), 
        .ZN(N60) );
  MUX3ND0 U3823 ( .I0(n3693), .I1(n3694), .I2(n3695), .S0(n3721), .S1(n3719), 
        .ZN(N59) );
  MUX3ND0 U3824 ( .I0(n3696), .I1(n3697), .I2(n3698), .S0(n3721), .S1(n3719), 
        .ZN(N58) );
  MUX3ND0 U3825 ( .I0(n3699), .I1(n3700), .I2(n3701), .S0(n3721), .S1(n3719), 
        .ZN(N57) );
  MUX3ND0 U3826 ( .I0(n3702), .I1(n3703), .I2(n3704), .S0(n3819), .S1(n3719), 
        .ZN(N56) );
  MUX3ND0 U3827 ( .I0(n3705), .I1(n3706), .I2(n3707), .S0(N49), .S1(n3719), 
        .ZN(N55) );
  MUX3ND0 U3828 ( .I0(n3708), .I1(n3709), .I2(n3710), .S0(N49), .S1(n3719), 
        .ZN(N54) );
  MUX3ND0 U3829 ( .I0(n3711), .I1(n3712), .I2(n3713), .S0(N49), .S1(n3719), 
        .ZN(N53) );
  MUX3ND0 U3830 ( .I0(n3714), .I1(n3715), .I2(n3716), .S0(N49), .S1(n3719), 
        .ZN(N52) );
  MUX2ND0 U3831 ( .I0(\Storage[2][0] ), .I1(\Storage[3][0] ), .S(n3722), .ZN(
        n3619) );
  MUX2ND0 U3832 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .S(n3723), .ZN(
        n3618) );
  MUX2ND0 U3833 ( .I0(\Storage[2][1] ), .I1(\Storage[3][1] ), .S(N48), .ZN(
        n3622) );
  MUX2ND0 U3834 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .S(n3723), .ZN(
        n3621) );
  MUX2ND0 U3835 ( .I0(\Storage[2][2] ), .I1(\Storage[3][2] ), .S(n3818), .ZN(
        n3625) );
  MUX2ND0 U3836 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .S(n3723), .ZN(
        n3624) );
  MUX2ND0 U3837 ( .I0(\Storage[2][3] ), .I1(\Storage[3][3] ), .S(n3722), .ZN(
        n3628) );
  MUX2ND0 U3838 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .S(n3723), .ZN(
        n3627) );
  MUX2ND0 U3839 ( .I0(\Storage[2][4] ), .I1(\Storage[3][4] ), .S(n3722), .ZN(
        n3631) );
  MUX2ND0 U3840 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .S(n3818), .ZN(
        n3630) );
  MUX2ND0 U3841 ( .I0(\Storage[2][5] ), .I1(\Storage[3][5] ), .S(n3722), .ZN(
        n3634) );
  MUX2ND0 U3842 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .S(n3722), .ZN(
        n3633) );
  MUX2ND0 U3843 ( .I0(\Storage[2][6] ), .I1(\Storage[3][6] ), .S(n3818), .ZN(
        n3637) );
  MUX2ND0 U3844 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .S(n3722), .ZN(
        n3636) );
  MUX2ND0 U3845 ( .I0(\Storage[2][7] ), .I1(\Storage[3][7] ), .S(n3723), .ZN(
        n3640) );
  MUX2ND0 U3846 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .S(n3723), .ZN(
        n3639) );
  MUX2ND0 U3847 ( .I0(\Storage[2][8] ), .I1(\Storage[3][8] ), .S(n3722), .ZN(
        n3643) );
  MUX2ND0 U3848 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .S(n3722), .ZN(
        n3642) );
  MUX2ND0 U3849 ( .I0(\Storage[2][9] ), .I1(\Storage[3][9] ), .S(n3722), .ZN(
        n3646) );
  MUX2ND0 U3850 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .S(n3722), .ZN(
        n3645) );
  MUX2ND0 U3851 ( .I0(\Storage[2][10] ), .I1(\Storage[3][10] ), .S(n3723), 
        .ZN(n3649) );
  MUX2ND0 U3852 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .S(n3723), 
        .ZN(n3648) );
  MUX2ND0 U3853 ( .I0(\Storage[2][11] ), .I1(\Storage[3][11] ), .S(n3723), 
        .ZN(n3652) );
  MUX2ND0 U3854 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .S(n3723), 
        .ZN(n3651) );
  MUX2ND0 U3855 ( .I0(\Storage[2][12] ), .I1(\Storage[3][12] ), .S(n3723), 
        .ZN(n3655) );
  MUX2ND0 U3856 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .S(n3724), 
        .ZN(n3654) );
  MUX2ND0 U3857 ( .I0(\Storage[2][13] ), .I1(\Storage[3][13] ), .S(n3724), 
        .ZN(n3658) );
  MUX2ND0 U3858 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .S(n3724), 
        .ZN(n3657) );
  MUX2ND0 U3859 ( .I0(\Storage[2][14] ), .I1(\Storage[3][14] ), .S(n3724), 
        .ZN(n3661) );
  MUX2ND0 U3860 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .S(n3724), 
        .ZN(n3660) );
  MUX2ND0 U3861 ( .I0(\Storage[2][15] ), .I1(\Storage[3][15] ), .S(n3818), 
        .ZN(n3664) );
  MUX2ND0 U3862 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .S(n3722), 
        .ZN(n3663) );
  MUX2ND0 U3863 ( .I0(\Storage[2][16] ), .I1(\Storage[3][16] ), .S(n3723), 
        .ZN(n3667) );
  MUX2ND0 U3864 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .S(N48), .ZN(
        n3666) );
  MUX2ND0 U3865 ( .I0(\Storage[2][17] ), .I1(\Storage[3][17] ), .S(n3724), 
        .ZN(n3670) );
  MUX2ND0 U3866 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .S(n3724), 
        .ZN(n3669) );
  MUX2ND0 U3867 ( .I0(\Storage[2][18] ), .I1(\Storage[3][18] ), .S(n3724), 
        .ZN(n3673) );
  MUX2ND0 U3868 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .S(n3724), 
        .ZN(n3672) );
  MUX2ND0 U3869 ( .I0(\Storage[2][19] ), .I1(\Storage[3][19] ), .S(n3724), 
        .ZN(n3676) );
  MUX2ND0 U3870 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .S(n3724), 
        .ZN(n3675) );
  MUX2ND0 U3871 ( .I0(\Storage[2][20] ), .I1(\Storage[3][20] ), .S(n3724), 
        .ZN(n3679) );
  MUX2ND0 U3872 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .S(n3724), 
        .ZN(n3678) );
  MUX2ND0 U3873 ( .I0(\Storage[2][21] ), .I1(\Storage[3][21] ), .S(n3724), 
        .ZN(n3682) );
  MUX2ND0 U3874 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .S(N48), .ZN(
        n3681) );
  MUX2ND0 U3875 ( .I0(\Storage[2][22] ), .I1(\Storage[3][22] ), .S(N48), .ZN(
        n3685) );
  MUX2ND0 U3876 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .S(N48), .ZN(
        n3684) );
  MUX2ND0 U3877 ( .I0(\Storage[2][23] ), .I1(\Storage[3][23] ), .S(N48), .ZN(
        n3688) );
  MUX2ND0 U3878 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .S(N48), .ZN(
        n3687) );
  MUX2ND0 U3879 ( .I0(\Storage[2][24] ), .I1(\Storage[3][24] ), .S(n3818), 
        .ZN(n3691) );
  MUX2ND0 U3880 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .S(n3818), 
        .ZN(n3690) );
  MUX2ND0 U3881 ( .I0(\Storage[2][25] ), .I1(\Storage[3][25] ), .S(n3724), 
        .ZN(n3694) );
  MUX2ND0 U3882 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .S(n3724), 
        .ZN(n3693) );
  MUX2ND0 U3883 ( .I0(\Storage[2][26] ), .I1(\Storage[3][26] ), .S(n3724), 
        .ZN(n3697) );
  MUX2ND0 U3884 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .S(n3724), 
        .ZN(n3696) );
  MUX2ND0 U3885 ( .I0(\Storage[2][27] ), .I1(\Storage[3][27] ), .S(n3722), 
        .ZN(n3700) );
  MUX2ND0 U3886 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .S(n3722), 
        .ZN(n3699) );
  MUX2ND0 U3887 ( .I0(\Storage[2][28] ), .I1(\Storage[3][28] ), .S(n3724), 
        .ZN(n3703) );
  MUX2ND0 U3888 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .S(n3722), 
        .ZN(n3702) );
  MUX2ND0 U3889 ( .I0(\Storage[2][29] ), .I1(\Storage[3][29] ), .S(n3818), 
        .ZN(n3706) );
  MUX2ND0 U3890 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .S(n3723), 
        .ZN(n3705) );
  MUX2ND0 U3891 ( .I0(\Storage[2][30] ), .I1(\Storage[3][30] ), .S(n3723), 
        .ZN(n3709) );
  MUX2ND0 U3892 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .S(n3723), 
        .ZN(n3708) );
  MUX2ND0 U3893 ( .I0(\Storage[2][31] ), .I1(\Storage[3][31] ), .S(n3818), 
        .ZN(n3712) );
  MUX2ND0 U3894 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .S(n3723), 
        .ZN(n3711) );
  MUX2ND0 U3895 ( .I0(\Storage[2][32] ), .I1(\Storage[3][32] ), .S(n3723), 
        .ZN(n3715) );
  MUX2ND0 U3896 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .S(n3724), 
        .ZN(n3714) );
endmodule


module PLLTop_0 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_0 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_0 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_0 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module FIFOStateM_AWid4_0 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [3:0] ReadAddr;
  output [3:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n1034, n1035, n1036, StateClockRaw, StateClock, N47, N48, N49, N50,
         N51, N67, N68, N69, N70, N71, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n66, n67, n68, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n83, n84, n85, n86, n87, n90,
         n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n141, n143, n144, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n69, n82, n88, n89, n93, n133, n134, n135, n136,
         n137, n138, n139, n140, n142, n145, n146, n161, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1032, n1033;
  wire   [2:0] NextState;
  wire   [3:0] OldReadAr;
  wire   [3:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n137), .CPN(StateClock), .Q(FullFIFO) );
  DFND1 EmptyFIFOr_reg ( .D(n6), .CPN(StateClock), .Q(n1034), .QN(n132) );
  OA21D1 U11 ( .A1(n172), .A2(n170), .B(n35), .Z(n44) );
  IAO21D1 U31 ( .A1(n73), .A2(n74), .B(n55), .ZN(n72) );
  OA21D1 U34 ( .A1(ReadAddr[2]), .A2(n76), .B(n75), .Z(n81) );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n202), .CPN(StateClock), .CDN(n1032), .Q(
        OldReadAr[3]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n237), .CPN(StateClock), .CDN(n1033), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n272), .CPN(StateClock), .CDN(n1032), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n306), .CPN(StateClock), .CDN(n1032), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n316), .CPN(StateClock), .CDN(n1033), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n326), .CPN(StateClock), .CDN(n1033), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n335), .CPN(StateClock), .CDN(n1032), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n344), .CPN(StateClock), .CDN(n1033), .Q(
        OldReadAr[1]) );
  DFNCND1 \NextState_reg[0]  ( .D(n383), .CPN(StateClock), .CDN(n1032), .Q(
        NextState[0]), .QN(n144) );
  DFNCND1 \NextState_reg[1]  ( .D(n419), .CPN(StateClock), .CDN(n1032), .Q(
        NextState[1]), .QN(n143) );
  DFNCND1 \NextState_reg[2]  ( .D(n455), .CPN(StateClock), .CDN(n1032), .Q(
        NextState[2]), .QN(n141) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n1032), 
        .QN(n170) );
  DFNCND1 WriteCmdr_reg ( .D(n620), .CPN(StateClock), .CDN(n1032), .Q(n1036)
         );
  DFNCND1 ReadCmdr_reg ( .D(n636), .CPN(StateClock), .CDN(n1032), .Q(n1035) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n1032), 
        .Q(n5), .QN(n171) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n1032), 
        .Q(n52), .QN(n172) );
  EDFCND1 \WriteAr_reg[1]  ( .D(n709), .E(n3), .CP(StateClock), .CDN(n1033), 
        .Q(WriteAddr[1]), .QN(n46) );
  EDFCND1 \ReadAr_reg[3]  ( .D(n744), .E(n1), .CP(StateClock), .CDN(n1033), 
        .Q(ReadAddr[3]), .QN(n163) );
  EDFCND1 \ReadAr_reg[2]  ( .D(n774), .E(n1), .CP(StateClock), .CDN(n1033), 
        .Q(ReadAddr[2]), .QN(n164) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n807), .E(n1), .CP(StateClock), .CDN(n1033), 
        .Q(ReadAddr[1]), .QN(n165) );
  EDFCND1 \ReadAr_reg[0]  ( .D(n837), .E(n1), .CP(StateClock), .CDN(n1033), 
        .Q(ReadAddr[0]), .QN(n166) );
  EDFCND1 \WriteAr_reg[3]  ( .D(n890), .E(n3), .CP(StateClock), .CDN(n1033), 
        .Q(WriteAddr[3]), .QN(n167) );
  EDFCND1 \WriteAr_reg[2]  ( .D(n925), .E(n3), .CP(StateClock), .CDN(n1033), 
        .Q(WriteAddr[2]), .QN(n168) );
  EDFCND1 \WriteAr_reg[0]  ( .D(n960), .E(n3), .CP(StateClock), .CDN(n1033), 
        .Q(WriteAddr[0]), .QN(n169) );
  BUFFD0 U3 ( .I(n867), .Z(n1) );
  BUFFD0 U4 ( .I(n1020), .Z(n2) );
  BUFFD0 U5 ( .I(n995), .Z(n3) );
  AN3D1 U6 ( .A1(n42), .A2(n1020), .A3(n56), .Z(n4) );
  INVD1 U7 ( .I(n4), .ZN(N71) );
  CKND2D0 U8 ( .A1(n868), .A2(n118), .ZN(N50) );
  BUFFD0 U9 ( .I(n9), .Z(n6) );
  BUFFD0 U10 ( .I(n8), .Z(n7) );
  BUFFD0 U12 ( .I(n132), .Z(n8) );
  BUFFD0 U13 ( .I(n10), .Z(n9) );
  BUFFD0 U14 ( .I(n11), .Z(n10) );
  BUFFD0 U15 ( .I(n12), .Z(n11) );
  BUFFD0 U16 ( .I(n13), .Z(n12) );
  BUFFD0 U17 ( .I(n14), .Z(n13) );
  BUFFD0 U18 ( .I(n15), .Z(n14) );
  BUFFD0 U19 ( .I(n16), .Z(n15) );
  BUFFD0 U20 ( .I(n17), .Z(n16) );
  BUFFD0 U21 ( .I(n18), .Z(n17) );
  BUFFD0 U22 ( .I(n19), .Z(n18) );
  BUFFD0 U23 ( .I(n20), .Z(n19) );
  BUFFD0 U24 ( .I(n21), .Z(n20) );
  BUFFD0 U25 ( .I(n22), .Z(n21) );
  BUFFD0 U26 ( .I(n23), .Z(n22) );
  BUFFD0 U27 ( .I(n24), .Z(n23) );
  BUFFD0 U28 ( .I(n25), .Z(n24) );
  BUFFD0 U29 ( .I(n26), .Z(n25) );
  BUFFD0 U30 ( .I(n27), .Z(n26) );
  BUFFD0 U32 ( .I(n28), .Z(n27) );
  BUFFD0 U33 ( .I(n29), .Z(n28) );
  BUFFD0 U35 ( .I(n30), .Z(n29) );
  BUFFD0 U36 ( .I(n31), .Z(n30) );
  BUFFD0 U37 ( .I(n32), .Z(n31) );
  BUFFD0 U38 ( .I(n33), .Z(n32) );
  BUFFD0 U39 ( .I(n34), .Z(n33) );
  BUFFD0 U40 ( .I(n69), .Z(n34) );
  BUFFD0 U41 ( .I(n82), .Z(n69) );
  BUFFD0 U42 ( .I(n88), .Z(n82) );
  BUFFD0 U43 ( .I(n89), .Z(n88) );
  BUFFD0 U44 ( .I(n93), .Z(n89) );
  BUFFD0 U45 ( .I(n133), .Z(n93) );
  BUFFD0 U46 ( .I(n134), .Z(n133) );
  BUFFD0 U47 ( .I(n135), .Z(n134) );
  BUFFD0 U48 ( .I(n136), .Z(n135) );
  BUFFD0 U49 ( .I(n147), .Z(n136) );
  BUFFD0 U50 ( .I(n139), .Z(n137) );
  OAI21D0 U51 ( .A1(n44), .A2(Reset), .B(FullFIFO), .ZN(n43) );
  BUFFD0 U52 ( .I(n43), .Z(n138) );
  BUFFD0 U53 ( .I(n140), .Z(n139) );
  BUFFD0 U54 ( .I(n142), .Z(n140) );
  BUFFD0 U55 ( .I(n145), .Z(n142) );
  BUFFD0 U56 ( .I(n146), .Z(n145) );
  BUFFD0 U57 ( .I(n161), .Z(n146) );
  BUFFD0 U58 ( .I(n173), .Z(n161) );
  BUFFD0 U59 ( .I(n174), .Z(n173) );
  BUFFD0 U60 ( .I(n175), .Z(n174) );
  BUFFD0 U61 ( .I(n176), .Z(n175) );
  BUFFD0 U62 ( .I(n177), .Z(n176) );
  BUFFD0 U63 ( .I(n178), .Z(n177) );
  BUFFD0 U64 ( .I(n179), .Z(n178) );
  BUFFD0 U65 ( .I(n180), .Z(n179) );
  BUFFD0 U66 ( .I(n181), .Z(n180) );
  BUFFD0 U67 ( .I(n182), .Z(n181) );
  BUFFD0 U68 ( .I(n183), .Z(n182) );
  BUFFD0 U69 ( .I(n184), .Z(n183) );
  BUFFD0 U70 ( .I(n185), .Z(n184) );
  BUFFD0 U71 ( .I(n186), .Z(n185) );
  BUFFD0 U72 ( .I(n187), .Z(n186) );
  BUFFD0 U73 ( .I(n188), .Z(n187) );
  BUFFD0 U74 ( .I(n189), .Z(n188) );
  BUFFD0 U75 ( .I(n190), .Z(n189) );
  BUFFD0 U76 ( .I(n191), .Z(n190) );
  BUFFD0 U77 ( .I(n192), .Z(n191) );
  BUFFD0 U78 ( .I(n193), .Z(n192) );
  BUFFD0 U79 ( .I(n194), .Z(n193) );
  BUFFD0 U80 ( .I(n195), .Z(n194) );
  BUFFD0 U81 ( .I(n196), .Z(n195) );
  BUFFD0 U82 ( .I(n197), .Z(n196) );
  BUFFD0 U83 ( .I(n198), .Z(n197) );
  BUFFD0 U84 ( .I(n199), .Z(n198) );
  BUFFD0 U85 ( .I(n200), .Z(n199) );
  BUFFD0 U86 ( .I(n201), .Z(n200) );
  BUFFD0 U87 ( .I(n151), .Z(n201) );
  BUFFD0 U88 ( .I(n204), .Z(n202) );
  BUFFD0 U89 ( .I(n150), .Z(n203) );
  BUFFD0 U90 ( .I(n205), .Z(n204) );
  BUFFD0 U91 ( .I(n206), .Z(n205) );
  BUFFD0 U92 ( .I(n207), .Z(n206) );
  BUFFD0 U93 ( .I(n208), .Z(n207) );
  BUFFD0 U94 ( .I(n209), .Z(n208) );
  BUFFD0 U95 ( .I(n210), .Z(n209) );
  BUFFD0 U96 ( .I(n211), .Z(n210) );
  BUFFD0 U97 ( .I(n212), .Z(n211) );
  BUFFD0 U98 ( .I(n213), .Z(n212) );
  BUFFD0 U99 ( .I(n214), .Z(n213) );
  BUFFD0 U100 ( .I(n215), .Z(n214) );
  BUFFD0 U101 ( .I(n216), .Z(n215) );
  BUFFD0 U102 ( .I(n217), .Z(n216) );
  BUFFD0 U103 ( .I(n218), .Z(n217) );
  BUFFD0 U104 ( .I(n219), .Z(n218) );
  BUFFD0 U105 ( .I(n220), .Z(n219) );
  BUFFD0 U106 ( .I(n221), .Z(n220) );
  BUFFD0 U107 ( .I(n222), .Z(n221) );
  BUFFD0 U108 ( .I(n223), .Z(n222) );
  BUFFD0 U109 ( .I(n224), .Z(n223) );
  BUFFD0 U110 ( .I(n225), .Z(n224) );
  BUFFD0 U111 ( .I(n226), .Z(n225) );
  BUFFD0 U112 ( .I(n227), .Z(n226) );
  BUFFD0 U113 ( .I(n228), .Z(n227) );
  BUFFD0 U114 ( .I(n229), .Z(n228) );
  BUFFD0 U115 ( .I(n230), .Z(n229) );
  BUFFD0 U116 ( .I(n231), .Z(n230) );
  BUFFD0 U117 ( .I(n232), .Z(n231) );
  BUFFD0 U118 ( .I(n233), .Z(n232) );
  BUFFD0 U119 ( .I(n234), .Z(n233) );
  BUFFD0 U120 ( .I(n235), .Z(n234) );
  BUFFD0 U121 ( .I(n236), .Z(n235) );
  BUFFD0 U122 ( .I(n203), .Z(n236) );
  BUFFD0 U123 ( .I(n239), .Z(n237) );
  BUFFD0 U124 ( .I(n148), .Z(n238) );
  BUFFD0 U125 ( .I(n240), .Z(n239) );
  BUFFD0 U126 ( .I(n241), .Z(n240) );
  BUFFD0 U127 ( .I(n242), .Z(n241) );
  BUFFD0 U128 ( .I(n243), .Z(n242) );
  BUFFD0 U129 ( .I(n244), .Z(n243) );
  BUFFD0 U130 ( .I(n245), .Z(n244) );
  BUFFD0 U131 ( .I(n246), .Z(n245) );
  BUFFD0 U132 ( .I(n247), .Z(n246) );
  BUFFD0 U133 ( .I(n248), .Z(n247) );
  BUFFD0 U134 ( .I(n249), .Z(n248) );
  BUFFD0 U135 ( .I(n250), .Z(n249) );
  BUFFD0 U136 ( .I(n251), .Z(n250) );
  BUFFD0 U137 ( .I(n252), .Z(n251) );
  BUFFD0 U138 ( .I(n253), .Z(n252) );
  BUFFD0 U139 ( .I(n254), .Z(n253) );
  BUFFD0 U140 ( .I(n255), .Z(n254) );
  BUFFD0 U141 ( .I(n256), .Z(n255) );
  BUFFD0 U142 ( .I(n257), .Z(n256) );
  BUFFD0 U143 ( .I(n258), .Z(n257) );
  BUFFD0 U144 ( .I(n259), .Z(n258) );
  BUFFD0 U145 ( .I(n260), .Z(n259) );
  BUFFD0 U146 ( .I(n261), .Z(n260) );
  BUFFD0 U147 ( .I(n262), .Z(n261) );
  BUFFD0 U148 ( .I(n263), .Z(n262) );
  BUFFD0 U149 ( .I(n264), .Z(n263) );
  BUFFD0 U150 ( .I(n265), .Z(n264) );
  BUFFD0 U151 ( .I(n266), .Z(n265) );
  BUFFD0 U152 ( .I(n267), .Z(n266) );
  BUFFD0 U153 ( .I(n268), .Z(n267) );
  BUFFD0 U154 ( .I(n269), .Z(n268) );
  BUFFD0 U155 ( .I(n270), .Z(n269) );
  BUFFD0 U156 ( .I(n271), .Z(n270) );
  BUFFD0 U157 ( .I(n238), .Z(n271) );
  MOAI22D0 U158 ( .A1(n166), .A2(n40), .B1(n40), .B2(n279), .ZN(n162) );
  BUFFD0 U159 ( .I(n274), .Z(n272) );
  BUFFD0 U160 ( .I(n162), .Z(n273) );
  BUFFD0 U161 ( .I(n275), .Z(n274) );
  BUFFD0 U162 ( .I(n276), .Z(n275) );
  BUFFD0 U163 ( .I(n277), .Z(n276) );
  BUFFD0 U164 ( .I(n278), .Z(n277) );
  BUFFD0 U165 ( .I(n304), .Z(n278) );
  BUFFD0 U166 ( .I(n280), .Z(n279) );
  BUFFD0 U167 ( .I(n281), .Z(n280) );
  BUFFD0 U168 ( .I(n282), .Z(n281) );
  BUFFD0 U169 ( .I(n283), .Z(n282) );
  BUFFD0 U170 ( .I(n284), .Z(n283) );
  BUFFD0 U171 ( .I(n285), .Z(n284) );
  BUFFD0 U172 ( .I(n286), .Z(n285) );
  BUFFD0 U173 ( .I(n287), .Z(n286) );
  BUFFD0 U174 ( .I(n288), .Z(n287) );
  BUFFD0 U175 ( .I(n289), .Z(n288) );
  BUFFD0 U176 ( .I(n290), .Z(n289) );
  BUFFD0 U177 ( .I(n291), .Z(n290) );
  BUFFD0 U178 ( .I(n292), .Z(n291) );
  BUFFD0 U179 ( .I(n293), .Z(n292) );
  BUFFD0 U180 ( .I(n294), .Z(n293) );
  BUFFD0 U181 ( .I(n295), .Z(n294) );
  BUFFD0 U182 ( .I(n296), .Z(n295) );
  BUFFD0 U183 ( .I(n297), .Z(n296) );
  BUFFD0 U184 ( .I(n298), .Z(n297) );
  BUFFD0 U185 ( .I(n299), .Z(n298) );
  BUFFD0 U186 ( .I(n300), .Z(n299) );
  BUFFD0 U187 ( .I(n301), .Z(n300) );
  BUFFD0 U188 ( .I(n302), .Z(n301) );
  BUFFD0 U189 ( .I(n668), .Z(n302) );
  BUFFD0 U190 ( .I(OldReadAr[0]), .Z(n303) );
  BUFFD0 U191 ( .I(n305), .Z(n304) );
  BUFFD0 U192 ( .I(n273), .Z(n305) );
  MOAI22D0 U193 ( .A1(n167), .A2(n45), .B1(n45), .B2(n311), .ZN(n155) );
  BUFFD0 U194 ( .I(n308), .Z(n306) );
  BUFFD0 U195 ( .I(n155), .Z(n307) );
  BUFFD0 U196 ( .I(n309), .Z(n308) );
  BUFFD0 U197 ( .I(n310), .Z(n309) );
  BUFFD0 U198 ( .I(n312), .Z(n310) );
  BUFFD0 U199 ( .I(n313), .Z(n311) );
  BUFFD0 U200 ( .I(n314), .Z(n312) );
  BUFFD0 U201 ( .I(n315), .Z(n313) );
  BUFFD0 U202 ( .I(n307), .Z(n314) );
  BUFFD0 U203 ( .I(n492), .Z(n315) );
  MOAI22D0 U204 ( .A1(n45), .A2(n46), .B1(n45), .B2(n321), .ZN(n154) );
  BUFFD0 U205 ( .I(n318), .Z(n316) );
  BUFFD0 U206 ( .I(n154), .Z(n317) );
  BUFFD0 U207 ( .I(n319), .Z(n318) );
  BUFFD0 U208 ( .I(n320), .Z(n319) );
  BUFFD0 U209 ( .I(n322), .Z(n320) );
  BUFFD0 U210 ( .I(n323), .Z(n321) );
  BUFFD0 U211 ( .I(n324), .Z(n322) );
  BUFFD0 U212 ( .I(n325), .Z(n323) );
  BUFFD0 U213 ( .I(n317), .Z(n324) );
  BUFFD0 U214 ( .I(n494), .Z(n325) );
  MOAI22D0 U215 ( .A1(n169), .A2(n45), .B1(n45), .B2(n330), .ZN(n153) );
  BUFFD0 U216 ( .I(n328), .Z(n326) );
  BUFFD0 U217 ( .I(n153), .Z(n327) );
  BUFFD0 U218 ( .I(n329), .Z(n328) );
  BUFFD0 U219 ( .I(n331), .Z(n329) );
  BUFFD0 U220 ( .I(n332), .Z(n330) );
  BUFFD0 U221 ( .I(n333), .Z(n331) );
  BUFFD0 U222 ( .I(n334), .Z(n332) );
  BUFFD0 U223 ( .I(n327), .Z(n333) );
  BUFFD0 U224 ( .I(n495), .Z(n334) );
  MOAI22D0 U225 ( .A1(n168), .A2(n45), .B1(n45), .B2(n339), .ZN(n152) );
  BUFFD0 U226 ( .I(n337), .Z(n335) );
  BUFFD0 U227 ( .I(n152), .Z(n336) );
  BUFFD0 U228 ( .I(n338), .Z(n337) );
  BUFFD0 U229 ( .I(n340), .Z(n338) );
  BUFFD0 U230 ( .I(n341), .Z(n339) );
  BUFFD0 U231 ( .I(n342), .Z(n340) );
  BUFFD0 U232 ( .I(n343), .Z(n341) );
  BUFFD0 U233 ( .I(n336), .Z(n342) );
  BUFFD0 U234 ( .I(n491), .Z(n343) );
  BUFFD0 U235 ( .I(n346), .Z(n344) );
  BUFFD0 U236 ( .I(n149), .Z(n345) );
  BUFFD0 U237 ( .I(n347), .Z(n346) );
  BUFFD0 U238 ( .I(n348), .Z(n347) );
  BUFFD0 U239 ( .I(n349), .Z(n348) );
  BUFFD0 U240 ( .I(n350), .Z(n349) );
  BUFFD0 U241 ( .I(n351), .Z(n350) );
  BUFFD0 U242 ( .I(n352), .Z(n351) );
  BUFFD0 U243 ( .I(n353), .Z(n352) );
  BUFFD0 U244 ( .I(n354), .Z(n353) );
  BUFFD0 U245 ( .I(n355), .Z(n354) );
  BUFFD0 U246 ( .I(n356), .Z(n355) );
  BUFFD0 U247 ( .I(n357), .Z(n356) );
  BUFFD0 U248 ( .I(n358), .Z(n357) );
  BUFFD0 U249 ( .I(n359), .Z(n358) );
  BUFFD0 U250 ( .I(n360), .Z(n359) );
  BUFFD0 U251 ( .I(n361), .Z(n360) );
  BUFFD0 U252 ( .I(n362), .Z(n361) );
  BUFFD0 U253 ( .I(n363), .Z(n362) );
  BUFFD0 U254 ( .I(n364), .Z(n363) );
  BUFFD0 U255 ( .I(n365), .Z(n364) );
  BUFFD0 U256 ( .I(n366), .Z(n365) );
  BUFFD0 U257 ( .I(n367), .Z(n366) );
  BUFFD0 U258 ( .I(n368), .Z(n367) );
  BUFFD0 U259 ( .I(n369), .Z(n368) );
  BUFFD0 U260 ( .I(n370), .Z(n369) );
  BUFFD0 U261 ( .I(n371), .Z(n370) );
  BUFFD0 U262 ( .I(n372), .Z(n371) );
  BUFFD0 U263 ( .I(n374), .Z(n372) );
  BUFFD0 U264 ( .I(OldReadAr[1]), .Z(n373) );
  BUFFD0 U265 ( .I(n375), .Z(n374) );
  BUFFD0 U266 ( .I(n376), .Z(n375) );
  BUFFD0 U267 ( .I(n377), .Z(n376) );
  BUFFD0 U268 ( .I(n345), .Z(n377) );
  IOA22D0 U269 ( .B1(n165), .B2(n40), .A1(n40), .A2(n667), .ZN(n149) );
  BUFFD0 U270 ( .I(n1036), .Z(n378) );
  BUFFD0 U271 ( .I(n378), .Z(n379) );
  BUFFD0 U272 ( .I(n379), .Z(n380) );
  BUFFD0 U273 ( .I(n380), .Z(n381) );
  BUFFD0 U274 ( .I(n381), .Z(n382) );
  BUFFD0 U275 ( .I(n385), .Z(n383) );
  BUFFD0 U276 ( .I(n386), .Z(n384) );
  BUFFD0 U277 ( .I(n387), .Z(n385) );
  BUFFD0 U278 ( .I(n388), .Z(n386) );
  BUFFD0 U279 ( .I(n389), .Z(n387) );
  BUFFD0 U280 ( .I(n390), .Z(n388) );
  BUFFD0 U281 ( .I(n391), .Z(n389) );
  BUFFD0 U282 ( .I(n392), .Z(n390) );
  BUFFD0 U283 ( .I(n393), .Z(n391) );
  BUFFD0 U284 ( .I(n394), .Z(n392) );
  BUFFD0 U285 ( .I(n395), .Z(n393) );
  BUFFD0 U286 ( .I(n396), .Z(n394) );
  BUFFD0 U287 ( .I(n397), .Z(n395) );
  BUFFD0 U288 ( .I(n398), .Z(n396) );
  BUFFD0 U289 ( .I(n399), .Z(n397) );
  BUFFD0 U290 ( .I(n400), .Z(n398) );
  BUFFD0 U291 ( .I(n401), .Z(n399) );
  BUFFD0 U292 ( .I(n402), .Z(n400) );
  BUFFD0 U293 ( .I(n403), .Z(n401) );
  BUFFD0 U294 ( .I(n404), .Z(n402) );
  BUFFD0 U295 ( .I(n405), .Z(n403) );
  BUFFD0 U296 ( .I(n406), .Z(n404) );
  BUFFD0 U297 ( .I(n407), .Z(n405) );
  BUFFD0 U298 ( .I(n408), .Z(n406) );
  BUFFD0 U299 ( .I(n409), .Z(n407) );
  BUFFD0 U300 ( .I(n410), .Z(n408) );
  BUFFD0 U301 ( .I(n411), .Z(n409) );
  BUFFD0 U302 ( .I(n412), .Z(n410) );
  BUFFD0 U303 ( .I(n159), .Z(n411) );
  BUFFD0 U304 ( .I(n413), .Z(n412) );
  BUFFD0 U305 ( .I(n414), .Z(n413) );
  BUFFD0 U306 ( .I(n415), .Z(n414) );
  BUFFD0 U307 ( .I(n416), .Z(n415) );
  BUFFD0 U308 ( .I(n417), .Z(n416) );
  BUFFD0 U309 ( .I(n418), .Z(n417) );
  BUFFD0 U310 ( .I(n144), .Z(n418) );
  BUFFD0 U311 ( .I(n421), .Z(n419) );
  BUFFD0 U312 ( .I(n422), .Z(n420) );
  BUFFD0 U313 ( .I(n423), .Z(n421) );
  BUFFD0 U314 ( .I(n424), .Z(n422) );
  BUFFD0 U315 ( .I(n425), .Z(n423) );
  BUFFD0 U316 ( .I(n426), .Z(n424) );
  BUFFD0 U317 ( .I(n427), .Z(n425) );
  BUFFD0 U318 ( .I(n428), .Z(n426) );
  BUFFD0 U319 ( .I(n429), .Z(n427) );
  BUFFD0 U320 ( .I(n430), .Z(n428) );
  BUFFD0 U321 ( .I(n431), .Z(n429) );
  BUFFD0 U322 ( .I(n432), .Z(n430) );
  BUFFD0 U323 ( .I(n433), .Z(n431) );
  BUFFD0 U324 ( .I(n434), .Z(n432) );
  BUFFD0 U325 ( .I(n435), .Z(n433) );
  BUFFD0 U326 ( .I(n436), .Z(n434) );
  BUFFD0 U327 ( .I(n437), .Z(n435) );
  BUFFD0 U328 ( .I(n438), .Z(n436) );
  BUFFD0 U329 ( .I(n439), .Z(n437) );
  BUFFD0 U330 ( .I(n440), .Z(n438) );
  BUFFD0 U331 ( .I(n441), .Z(n439) );
  BUFFD0 U332 ( .I(n442), .Z(n440) );
  BUFFD0 U333 ( .I(n443), .Z(n441) );
  BUFFD0 U334 ( .I(n444), .Z(n442) );
  BUFFD0 U335 ( .I(n445), .Z(n443) );
  BUFFD0 U336 ( .I(n446), .Z(n444) );
  BUFFD0 U337 ( .I(n447), .Z(n445) );
  BUFFD0 U338 ( .I(n448), .Z(n446) );
  BUFFD0 U339 ( .I(n158), .Z(n447) );
  BUFFD0 U340 ( .I(n449), .Z(n448) );
  BUFFD0 U341 ( .I(n450), .Z(n449) );
  BUFFD0 U342 ( .I(n451), .Z(n450) );
  BUFFD0 U343 ( .I(n452), .Z(n451) );
  BUFFD0 U344 ( .I(n453), .Z(n452) );
  BUFFD0 U345 ( .I(n454), .Z(n453) );
  BUFFD0 U346 ( .I(n143), .Z(n454) );
  BUFFD0 U347 ( .I(n457), .Z(n455) );
  BUFFD0 U348 ( .I(n458), .Z(n456) );
  BUFFD0 U349 ( .I(n459), .Z(n457) );
  BUFFD0 U350 ( .I(n460), .Z(n458) );
  BUFFD0 U351 ( .I(n461), .Z(n459) );
  BUFFD0 U352 ( .I(n462), .Z(n460) );
  BUFFD0 U353 ( .I(n463), .Z(n461) );
  BUFFD0 U354 ( .I(n464), .Z(n462) );
  BUFFD0 U355 ( .I(n465), .Z(n463) );
  BUFFD0 U356 ( .I(n466), .Z(n464) );
  BUFFD0 U357 ( .I(n467), .Z(n465) );
  BUFFD0 U358 ( .I(n468), .Z(n466) );
  BUFFD0 U359 ( .I(n469), .Z(n467) );
  BUFFD0 U360 ( .I(n470), .Z(n468) );
  BUFFD0 U361 ( .I(n471), .Z(n469) );
  BUFFD0 U362 ( .I(n472), .Z(n470) );
  BUFFD0 U363 ( .I(n473), .Z(n471) );
  BUFFD0 U364 ( .I(n474), .Z(n472) );
  BUFFD0 U365 ( .I(n475), .Z(n473) );
  BUFFD0 U366 ( .I(n476), .Z(n474) );
  BUFFD0 U367 ( .I(n477), .Z(n475) );
  BUFFD0 U368 ( .I(n478), .Z(n476) );
  BUFFD0 U369 ( .I(n479), .Z(n477) );
  BUFFD0 U370 ( .I(n480), .Z(n478) );
  BUFFD0 U371 ( .I(n481), .Z(n479) );
  BUFFD0 U372 ( .I(n482), .Z(n480) );
  BUFFD0 U373 ( .I(n483), .Z(n481) );
  BUFFD0 U374 ( .I(n484), .Z(n482) );
  BUFFD0 U375 ( .I(n156), .Z(n483) );
  BUFFD0 U376 ( .I(n485), .Z(n484) );
  BUFFD0 U377 ( .I(n486), .Z(n485) );
  BUFFD0 U378 ( .I(n487), .Z(n486) );
  BUFFD0 U379 ( .I(n488), .Z(n487) );
  BUFFD0 U380 ( .I(n489), .Z(n488) );
  BUFFD0 U381 ( .I(n490), .Z(n489) );
  BUFFD0 U382 ( .I(n141), .Z(n490) );
  CKBD0 U383 ( .CLK(n157), .C(n630) );
  ND4D0 U384 ( .A1(n58), .A2(n47), .A3(n59), .A4(n60), .ZN(n57) );
  BUFFD0 U385 ( .I(n496), .Z(n491) );
  BUFFD0 U386 ( .I(n497), .Z(n492) );
  BUFFD0 U387 ( .I(n382), .Z(n493) );
  BUFFD0 U388 ( .I(n499), .Z(n494) );
  BUFFD0 U389 ( .I(n500), .Z(n495) );
  BUFFD0 U390 ( .I(n501), .Z(n496) );
  BUFFD0 U391 ( .I(n502), .Z(n497) );
  BUFFD0 U392 ( .I(n493), .Z(n498) );
  BUFFD0 U393 ( .I(n504), .Z(n499) );
  BUFFD0 U394 ( .I(n505), .Z(n500) );
  BUFFD0 U395 ( .I(n506), .Z(n501) );
  BUFFD0 U396 ( .I(n507), .Z(n502) );
  BUFFD0 U397 ( .I(n498), .Z(n503) );
  BUFFD0 U398 ( .I(n509), .Z(n504) );
  BUFFD0 U399 ( .I(n510), .Z(n505) );
  BUFFD0 U400 ( .I(n511), .Z(n506) );
  BUFFD0 U401 ( .I(n512), .Z(n507) );
  BUFFD0 U402 ( .I(n503), .Z(n508) );
  BUFFD0 U403 ( .I(n514), .Z(n509) );
  BUFFD0 U404 ( .I(n515), .Z(n510) );
  BUFFD0 U405 ( .I(n516), .Z(n511) );
  BUFFD0 U406 ( .I(n517), .Z(n512) );
  BUFFD0 U407 ( .I(n508), .Z(n513) );
  BUFFD0 U408 ( .I(n519), .Z(n514) );
  BUFFD0 U409 ( .I(n520), .Z(n515) );
  BUFFD0 U410 ( .I(n521), .Z(n516) );
  BUFFD0 U411 ( .I(n522), .Z(n517) );
  BUFFD0 U412 ( .I(n513), .Z(n518) );
  BUFFD0 U413 ( .I(n524), .Z(n519) );
  BUFFD0 U414 ( .I(n525), .Z(n520) );
  BUFFD0 U415 ( .I(n526), .Z(n521) );
  BUFFD0 U416 ( .I(n527), .Z(n522) );
  BUFFD0 U417 ( .I(n518), .Z(n523) );
  BUFFD0 U418 ( .I(n529), .Z(n524) );
  BUFFD0 U419 ( .I(n530), .Z(n525) );
  BUFFD0 U420 ( .I(n531), .Z(n526) );
  BUFFD0 U421 ( .I(n532), .Z(n527) );
  BUFFD0 U422 ( .I(n523), .Z(n528) );
  BUFFD0 U423 ( .I(n534), .Z(n529) );
  BUFFD0 U424 ( .I(n535), .Z(n530) );
  BUFFD0 U425 ( .I(n536), .Z(n531) );
  BUFFD0 U426 ( .I(n537), .Z(n532) );
  BUFFD0 U427 ( .I(n528), .Z(n533) );
  BUFFD0 U428 ( .I(n539), .Z(n534) );
  BUFFD0 U429 ( .I(n540), .Z(n535) );
  BUFFD0 U430 ( .I(n541), .Z(n536) );
  BUFFD0 U431 ( .I(n542), .Z(n537) );
  BUFFD0 U432 ( .I(n533), .Z(n538) );
  BUFFD0 U433 ( .I(n544), .Z(n539) );
  BUFFD0 U434 ( .I(n545), .Z(n540) );
  BUFFD0 U435 ( .I(n546), .Z(n541) );
  BUFFD0 U436 ( .I(n547), .Z(n542) );
  BUFFD0 U437 ( .I(n538), .Z(n543) );
  BUFFD0 U438 ( .I(n549), .Z(n544) );
  BUFFD0 U439 ( .I(n550), .Z(n545) );
  BUFFD0 U440 ( .I(n551), .Z(n546) );
  BUFFD0 U441 ( .I(n552), .Z(n547) );
  BUFFD0 U442 ( .I(n543), .Z(n548) );
  BUFFD0 U443 ( .I(n554), .Z(n549) );
  BUFFD0 U444 ( .I(n555), .Z(n550) );
  BUFFD0 U445 ( .I(n556), .Z(n551) );
  BUFFD0 U446 ( .I(n557), .Z(n552) );
  BUFFD0 U447 ( .I(n548), .Z(n553) );
  BUFFD0 U448 ( .I(n559), .Z(n554) );
  BUFFD0 U449 ( .I(n560), .Z(n555) );
  BUFFD0 U450 ( .I(n561), .Z(n556) );
  BUFFD0 U451 ( .I(n562), .Z(n557) );
  BUFFD0 U452 ( .I(n553), .Z(n558) );
  BUFFD0 U453 ( .I(n564), .Z(n559) );
  BUFFD0 U454 ( .I(n565), .Z(n560) );
  BUFFD0 U455 ( .I(n566), .Z(n561) );
  BUFFD0 U456 ( .I(n567), .Z(n562) );
  BUFFD0 U457 ( .I(n558), .Z(n563) );
  BUFFD0 U458 ( .I(n569), .Z(n564) );
  BUFFD0 U459 ( .I(n570), .Z(n565) );
  BUFFD0 U460 ( .I(n571), .Z(n566) );
  BUFFD0 U461 ( .I(n572), .Z(n567) );
  BUFFD0 U462 ( .I(n563), .Z(n568) );
  BUFFD0 U463 ( .I(n574), .Z(n569) );
  BUFFD0 U464 ( .I(n575), .Z(n570) );
  BUFFD0 U465 ( .I(n576), .Z(n571) );
  BUFFD0 U466 ( .I(n577), .Z(n572) );
  BUFFD0 U467 ( .I(n568), .Z(n573) );
  BUFFD0 U468 ( .I(n579), .Z(n574) );
  BUFFD0 U469 ( .I(n580), .Z(n575) );
  BUFFD0 U470 ( .I(n581), .Z(n576) );
  BUFFD0 U471 ( .I(n582), .Z(n577) );
  BUFFD0 U472 ( .I(n573), .Z(n578) );
  BUFFD0 U473 ( .I(n584), .Z(n579) );
  BUFFD0 U474 ( .I(n585), .Z(n580) );
  BUFFD0 U475 ( .I(n586), .Z(n581) );
  BUFFD0 U476 ( .I(n587), .Z(n582) );
  BUFFD0 U477 ( .I(n578), .Z(n583) );
  BUFFD0 U478 ( .I(n589), .Z(n584) );
  BUFFD0 U479 ( .I(n590), .Z(n585) );
  BUFFD0 U480 ( .I(n591), .Z(n586) );
  BUFFD0 U481 ( .I(n592), .Z(n587) );
  BUFFD0 U482 ( .I(n583), .Z(n588) );
  BUFFD0 U483 ( .I(n594), .Z(n589) );
  BUFFD0 U484 ( .I(n595), .Z(n590) );
  BUFFD0 U485 ( .I(n596), .Z(n591) );
  BUFFD0 U486 ( .I(n597), .Z(n592) );
  BUFFD0 U487 ( .I(n588), .Z(n593) );
  BUFFD0 U488 ( .I(n599), .Z(n594) );
  BUFFD0 U489 ( .I(n600), .Z(n595) );
  BUFFD0 U490 ( .I(n601), .Z(n596) );
  BUFFD0 U491 ( .I(n602), .Z(n597) );
  BUFFD0 U492 ( .I(n593), .Z(n598) );
  BUFFD0 U493 ( .I(n604), .Z(n599) );
  BUFFD0 U494 ( .I(n605), .Z(n600) );
  BUFFD0 U495 ( .I(n606), .Z(n601) );
  BUFFD0 U496 ( .I(n607), .Z(n602) );
  BUFFD0 U497 ( .I(n598), .Z(n603) );
  BUFFD0 U498 ( .I(n609), .Z(n604) );
  BUFFD0 U499 ( .I(n610), .Z(n605) );
  BUFFD0 U500 ( .I(n611), .Z(n606) );
  BUFFD0 U501 ( .I(n612), .Z(n607) );
  BUFFD0 U502 ( .I(n603), .Z(n608) );
  BUFFD0 U503 ( .I(n614), .Z(n609) );
  BUFFD0 U504 ( .I(n615), .Z(n610) );
  BUFFD0 U505 ( .I(n616), .Z(n611) );
  BUFFD0 U506 ( .I(n617), .Z(n612) );
  BUFFD0 U507 ( .I(n608), .Z(n613) );
  BUFFD0 U508 ( .I(n619), .Z(n614) );
  BUFFD0 U509 ( .I(n625), .Z(n615) );
  BUFFD0 U510 ( .I(n627), .Z(n616) );
  BUFFD0 U511 ( .I(n628), .Z(n617) );
  BUFFD0 U512 ( .I(n613), .Z(n618) );
  BUFFD0 U513 ( .I(n632), .Z(n619) );
  BUFFD0 U514 ( .I(n622), .Z(n620) );
  BUFFD0 U515 ( .I(n57), .Z(n621) );
  BUFFD0 U516 ( .I(n623), .Z(n622) );
  BUFFD0 U517 ( .I(n624), .Z(n623) );
  BUFFD0 U518 ( .I(n629), .Z(n624) );
  BUFFD0 U519 ( .I(n631), .Z(n625) );
  CKBXD0 U520 ( .I(n618), .Z(WriteCmd) );
  BUFFD0 U521 ( .I(n633), .Z(n627) );
  BUFFD0 U522 ( .I(OldWriteAr[3]), .Z(n628) );
  BUFFD0 U523 ( .I(n630), .Z(n629) );
  OAI21D0 U524 ( .A1(n56), .A2(n47), .B(n621), .ZN(n157) );
  BUFFD0 U525 ( .I(n634), .Z(n631) );
  BUFFD0 U526 ( .I(OldWriteAr[1]), .Z(n632) );
  BUFFD0 U527 ( .I(OldWriteAr[2]), .Z(n633) );
  BUFFD0 U528 ( .I(OldWriteAr[0]), .Z(n634) );
  ND4D0 U529 ( .A1(n121), .A2(n119), .A3(n122), .A4(n123), .ZN(n120) );
  BUFFD0 U530 ( .I(n120), .Z(n635) );
  ND2D0 U531 ( .A1(ReadCmd), .A2(n868), .ZN(n118) );
  BUFFD0 U532 ( .I(n637), .Z(n636) );
  BUFFD0 U533 ( .I(n638), .Z(n637) );
  BUFFD0 U534 ( .I(n639), .Z(n638) );
  BUFFD0 U535 ( .I(n640), .Z(n639) );
  BUFFD0 U536 ( .I(n641), .Z(n640) );
  BUFFD0 U537 ( .I(n642), .Z(n641) );
  BUFFD0 U538 ( .I(n643), .Z(n642) );
  BUFFD0 U539 ( .I(n644), .Z(n643) );
  BUFFD0 U540 ( .I(n645), .Z(n644) );
  BUFFD0 U541 ( .I(n646), .Z(n645) );
  BUFFD0 U542 ( .I(n647), .Z(n646) );
  BUFFD0 U543 ( .I(n648), .Z(n647) );
  BUFFD0 U544 ( .I(n649), .Z(n648) );
  BUFFD0 U545 ( .I(n650), .Z(n649) );
  BUFFD0 U546 ( .I(n651), .Z(n650) );
  BUFFD0 U547 ( .I(n652), .Z(n651) );
  BUFFD0 U548 ( .I(n653), .Z(n652) );
  BUFFD0 U549 ( .I(n654), .Z(n653) );
  BUFFD0 U550 ( .I(n655), .Z(n654) );
  BUFFD0 U551 ( .I(n656), .Z(n655) );
  BUFFD0 U552 ( .I(n657), .Z(n656) );
  BUFFD0 U553 ( .I(n658), .Z(n657) );
  BUFFD0 U554 ( .I(n659), .Z(n658) );
  BUFFD0 U555 ( .I(n660), .Z(n659) );
  BUFFD0 U556 ( .I(n661), .Z(n660) );
  BUFFD0 U557 ( .I(n662), .Z(n661) );
  BUFFD0 U558 ( .I(n663), .Z(n662) );
  BUFFD0 U559 ( .I(n664), .Z(n663) );
  BUFFD0 U560 ( .I(n672), .Z(n664) );
  OAI21D0 U561 ( .A1(n118), .A2(n119), .B(n635), .ZN(n160) );
  BUFFD0 U562 ( .I(OldReadAr[3]), .Z(n665) );
  BUFFD0 U563 ( .I(OldReadAr[2]), .Z(n666) );
  BUFFD0 U564 ( .I(n669), .Z(n667) );
  BUFFD0 U565 ( .I(n674), .Z(n668) );
  BUFFD0 U566 ( .I(n675), .Z(n669) );
  BUFFD0 U567 ( .I(n41), .Z(n670) );
  BUFFD0 U568 ( .I(n39), .Z(n671) );
  BUFFD0 U569 ( .I(n673), .Z(n672) );
  BUFFD0 U570 ( .I(n160), .Z(n673) );
  BUFFD0 U571 ( .I(n676), .Z(n674) );
  BUFFD0 U572 ( .I(n373), .Z(n675) );
  BUFFD0 U573 ( .I(n303), .Z(n676) );
  BUFFD0 U574 ( .I(n678), .Z(EmptyFIFO) );
  BUFFD0 U575 ( .I(n679), .Z(n678) );
  BUFFD0 U576 ( .I(n680), .Z(n679) );
  BUFFD0 U577 ( .I(n681), .Z(n680) );
  BUFFD0 U578 ( .I(n682), .Z(n681) );
  BUFFD0 U579 ( .I(n683), .Z(n682) );
  BUFFD0 U580 ( .I(n684), .Z(n683) );
  BUFFD0 U581 ( .I(n685), .Z(n684) );
  BUFFD0 U582 ( .I(n686), .Z(n685) );
  BUFFD0 U583 ( .I(n687), .Z(n686) );
  BUFFD0 U584 ( .I(n688), .Z(n687) );
  BUFFD0 U585 ( .I(n689), .Z(n688) );
  BUFFD0 U586 ( .I(n690), .Z(n689) );
  BUFFD0 U587 ( .I(n691), .Z(n690) );
  BUFFD0 U588 ( .I(n692), .Z(n691) );
  BUFFD0 U589 ( .I(n693), .Z(n692) );
  BUFFD0 U590 ( .I(n694), .Z(n693) );
  BUFFD0 U591 ( .I(n695), .Z(n694) );
  BUFFD0 U592 ( .I(n696), .Z(n695) );
  BUFFD0 U593 ( .I(n697), .Z(n696) );
  BUFFD0 U594 ( .I(n698), .Z(n697) );
  BUFFD0 U595 ( .I(n699), .Z(n698) );
  BUFFD0 U596 ( .I(n700), .Z(n699) );
  BUFFD0 U597 ( .I(n701), .Z(n700) );
  BUFFD0 U598 ( .I(n702), .Z(n701) );
  BUFFD0 U599 ( .I(n703), .Z(n702) );
  BUFFD0 U600 ( .I(n704), .Z(n703) );
  BUFFD0 U601 ( .I(n705), .Z(n704) );
  BUFFD0 U602 ( .I(n706), .Z(n705) );
  BUFFD0 U603 ( .I(n1034), .Z(n706) );
  BUFFD0 U604 ( .I(n1035), .Z(n707) );
  CKBD0 U605 ( .CLK(n707), .C(ReadCmd) );
  BUFFD0 U606 ( .I(n712), .Z(n709) );
  BUFFD0 U607 ( .I(N68), .Z(n710) );
  BUFFD0 U608 ( .I(n710), .Z(n711) );
  BUFFD0 U609 ( .I(n713), .Z(n712) );
  BUFFD0 U610 ( .I(n714), .Z(n713) );
  BUFFD0 U611 ( .I(n715), .Z(n714) );
  BUFFD0 U612 ( .I(n716), .Z(n715) );
  BUFFD0 U613 ( .I(n717), .Z(n716) );
  BUFFD0 U614 ( .I(n718), .Z(n717) );
  BUFFD0 U615 ( .I(n719), .Z(n718) );
  BUFFD0 U616 ( .I(n720), .Z(n719) );
  BUFFD0 U617 ( .I(n721), .Z(n720) );
  BUFFD0 U618 ( .I(n722), .Z(n721) );
  BUFFD0 U619 ( .I(n723), .Z(n722) );
  BUFFD0 U620 ( .I(n724), .Z(n723) );
  BUFFD0 U621 ( .I(n725), .Z(n724) );
  BUFFD0 U622 ( .I(n726), .Z(n725) );
  BUFFD0 U623 ( .I(n727), .Z(n726) );
  BUFFD0 U624 ( .I(n728), .Z(n727) );
  BUFFD0 U625 ( .I(n729), .Z(n728) );
  BUFFD0 U626 ( .I(n730), .Z(n729) );
  BUFFD0 U627 ( .I(n731), .Z(n730) );
  BUFFD0 U628 ( .I(n732), .Z(n731) );
  BUFFD0 U629 ( .I(n733), .Z(n732) );
  BUFFD0 U630 ( .I(n734), .Z(n733) );
  BUFFD0 U631 ( .I(n735), .Z(n734) );
  BUFFD0 U632 ( .I(n736), .Z(n735) );
  BUFFD0 U633 ( .I(n737), .Z(n736) );
  BUFFD0 U634 ( .I(n738), .Z(n737) );
  BUFFD0 U635 ( .I(n739), .Z(n738) );
  BUFFD0 U636 ( .I(n740), .Z(n739) );
  BUFFD0 U637 ( .I(n741), .Z(n740) );
  BUFFD0 U638 ( .I(n742), .Z(n741) );
  BUFFD0 U639 ( .I(n743), .Z(n742) );
  BUFFD0 U640 ( .I(n711), .Z(n743) );
  BUFFD0 U641 ( .I(n745), .Z(n744) );
  BUFFD0 U642 ( .I(n751), .Z(n745) );
  BUFFD0 U643 ( .I(n747), .Z(n746) );
  BUFFD0 U644 ( .I(n748), .Z(n747) );
  BUFFD0 U645 ( .I(n749), .Z(n748) );
  BUFFD0 U646 ( .I(n750), .Z(n749) );
  CKBD0 U647 ( .CLK(n163), .C(n924) );
  BUFFD0 U648 ( .I(n752), .Z(n750) );
  BUFFD0 U649 ( .I(N51), .Z(n751) );
  BUFFD0 U650 ( .I(n753), .Z(n752) );
  BUFFD0 U651 ( .I(n754), .Z(n753) );
  BUFFD0 U652 ( .I(n755), .Z(n754) );
  BUFFD0 U653 ( .I(n756), .Z(n755) );
  BUFFD0 U654 ( .I(n757), .Z(n756) );
  BUFFD0 U655 ( .I(n758), .Z(n757) );
  BUFFD0 U656 ( .I(n759), .Z(n758) );
  BUFFD0 U657 ( .I(n760), .Z(n759) );
  BUFFD0 U658 ( .I(n761), .Z(n760) );
  BUFFD0 U659 ( .I(n762), .Z(n761) );
  BUFFD0 U660 ( .I(n763), .Z(n762) );
  BUFFD0 U661 ( .I(n764), .Z(n763) );
  BUFFD0 U662 ( .I(n765), .Z(n764) );
  BUFFD0 U663 ( .I(n766), .Z(n765) );
  BUFFD0 U664 ( .I(n767), .Z(n766) );
  BUFFD0 U665 ( .I(n768), .Z(n767) );
  BUFFD0 U666 ( .I(n769), .Z(n768) );
  BUFFD0 U667 ( .I(n770), .Z(n769) );
  BUFFD0 U668 ( .I(n771), .Z(n770) );
  BUFFD0 U669 ( .I(n772), .Z(n771) );
  BUFFD0 U670 ( .I(n773), .Z(n772) );
  BUFFD0 U671 ( .I(n112), .Z(n773) );
  XNR2D0 U672 ( .A1(n924), .A2(n129), .ZN(n112) );
  BUFFD0 U673 ( .I(n775), .Z(n774) );
  BUFFD0 U674 ( .I(n776), .Z(n775) );
  BUFFD0 U675 ( .I(n777), .Z(n776) );
  BUFFD0 U676 ( .I(n778), .Z(n777) );
  BUFFD0 U677 ( .I(n779), .Z(n778) );
  BUFFD0 U678 ( .I(n780), .Z(n779) );
  BUFFD0 U679 ( .I(n781), .Z(n780) );
  BUFFD0 U680 ( .I(n782), .Z(n781) );
  BUFFD0 U681 ( .I(n783), .Z(n782) );
  BUFFD0 U682 ( .I(n784), .Z(n783) );
  BUFFD0 U683 ( .I(n785), .Z(n784) );
  BUFFD0 U684 ( .I(n786), .Z(n785) );
  BUFFD0 U685 ( .I(n787), .Z(n786) );
  BUFFD0 U686 ( .I(n788), .Z(n787) );
  BUFFD0 U687 ( .I(n789), .Z(n788) );
  BUFFD0 U688 ( .I(n790), .Z(n789) );
  BUFFD0 U689 ( .I(n791), .Z(n790) );
  BUFFD0 U690 ( .I(n792), .Z(n791) );
  BUFFD0 U691 ( .I(n793), .Z(n792) );
  BUFFD0 U692 ( .I(n794), .Z(n793) );
  BUFFD0 U693 ( .I(n795), .Z(n794) );
  BUFFD0 U694 ( .I(n796), .Z(n795) );
  BUFFD0 U695 ( .I(n797), .Z(n796) );
  BUFFD0 U696 ( .I(n798), .Z(n797) );
  BUFFD0 U697 ( .I(n799), .Z(n798) );
  BUFFD0 U698 ( .I(n800), .Z(n799) );
  BUFFD0 U699 ( .I(n801), .Z(n800) );
  BUFFD0 U700 ( .I(n802), .Z(n801) );
  BUFFD0 U701 ( .I(n803), .Z(n802) );
  BUFFD0 U702 ( .I(n804), .Z(n803) );
  BUFFD0 U703 ( .I(n805), .Z(n804) );
  BUFFD0 U704 ( .I(N49), .Z(n805) );
  CKBD0 U705 ( .CLK(ReadAddr[2]), .C(n806) );
  OAI21D0 U706 ( .A1(n130), .A2(n806), .B(n129), .ZN(n114) );
  BUFFD0 U707 ( .I(n809), .Z(n807) );
  BUFFD0 U708 ( .I(n810), .Z(n808) );
  BUFFD0 U709 ( .I(N48), .Z(n809) );
  BUFFD0 U710 ( .I(n811), .Z(n810) );
  BUFFD0 U711 ( .I(n812), .Z(n811) );
  BUFFD0 U712 ( .I(n813), .Z(n812) );
  BUFFD0 U713 ( .I(n814), .Z(n813) );
  BUFFD0 U714 ( .I(n815), .Z(n814) );
  BUFFD0 U715 ( .I(n816), .Z(n815) );
  BUFFD0 U716 ( .I(n817), .Z(n816) );
  BUFFD0 U717 ( .I(n818), .Z(n817) );
  BUFFD0 U718 ( .I(n819), .Z(n818) );
  BUFFD0 U719 ( .I(n820), .Z(n819) );
  BUFFD0 U720 ( .I(n821), .Z(n820) );
  BUFFD0 U721 ( .I(n822), .Z(n821) );
  BUFFD0 U722 ( .I(n823), .Z(n822) );
  BUFFD0 U723 ( .I(n824), .Z(n823) );
  BUFFD0 U724 ( .I(n825), .Z(n824) );
  BUFFD0 U725 ( .I(n826), .Z(n825) );
  BUFFD0 U726 ( .I(n827), .Z(n826) );
  BUFFD0 U727 ( .I(n828), .Z(n827) );
  BUFFD0 U728 ( .I(n829), .Z(n828) );
  BUFFD0 U729 ( .I(n830), .Z(n829) );
  BUFFD0 U730 ( .I(n831), .Z(n830) );
  BUFFD0 U731 ( .I(n832), .Z(n831) );
  BUFFD0 U732 ( .I(n833), .Z(n832) );
  BUFFD0 U733 ( .I(n834), .Z(n833) );
  BUFFD0 U734 ( .I(n835), .Z(n834) );
  BUFFD0 U735 ( .I(n131), .Z(n835) );
  BUFFD0 U736 ( .I(ReadAddr[1]), .Z(n836) );
  XNR2D0 U737 ( .A1(n836), .A2(n838), .ZN(n131) );
  BUFFD0 U738 ( .I(n839), .Z(n837) );
  BUFFD0 U739 ( .I(n840), .Z(n838) );
  BUFFD0 U740 ( .I(n841), .Z(n839) );
  BUFFD0 U741 ( .I(n842), .Z(n840) );
  BUFFD0 U742 ( .I(n843), .Z(n841) );
  BUFFD0 U743 ( .I(n844), .Z(n842) );
  BUFFD0 U744 ( .I(n845), .Z(n843) );
  BUFFD0 U745 ( .I(n846), .Z(n844) );
  BUFFD0 U746 ( .I(n847), .Z(n845) );
  BUFFD0 U747 ( .I(n848), .Z(n846) );
  BUFFD0 U748 ( .I(n849), .Z(n847) );
  BUFFD0 U749 ( .I(n850), .Z(n848) );
  BUFFD0 U750 ( .I(N47), .Z(n849) );
  BUFFD0 U751 ( .I(n851), .Z(n850) );
  BUFFD0 U752 ( .I(n852), .Z(n851) );
  BUFFD0 U753 ( .I(n853), .Z(n852) );
  BUFFD0 U754 ( .I(n854), .Z(n853) );
  BUFFD0 U755 ( .I(n855), .Z(n854) );
  BUFFD0 U756 ( .I(n856), .Z(n855) );
  BUFFD0 U757 ( .I(n857), .Z(n856) );
  BUFFD0 U758 ( .I(n858), .Z(n857) );
  BUFFD0 U759 ( .I(n859), .Z(n858) );
  BUFFD0 U760 ( .I(n860), .Z(n859) );
  BUFFD0 U761 ( .I(n861), .Z(n860) );
  BUFFD0 U762 ( .I(n862), .Z(n861) );
  BUFFD0 U763 ( .I(n863), .Z(n862) );
  BUFFD0 U764 ( .I(n864), .Z(n863) );
  BUFFD0 U765 ( .I(n865), .Z(n864) );
  BUFFD0 U766 ( .I(n866), .Z(n865) );
  BUFFD0 U767 ( .I(ReadAddr[0]), .Z(n866) );
  BUFFD0 U768 ( .I(n871), .Z(n867) );
  BUFFD0 U769 ( .I(n869), .Z(n868) );
  BUFFD0 U770 ( .I(n870), .Z(n869) );
  BUFFD0 U771 ( .I(n2), .Z(n870) );
  BUFFD0 U772 ( .I(N50), .Z(n871) );
  BUFFD0 U773 ( .I(n35), .Z(n872) );
  BUFFD0 U774 ( .I(n872), .Z(n873) );
  BUFFD0 U775 ( .I(n873), .Z(n874) );
  BUFFD0 U776 ( .I(n874), .Z(n875) );
  BUFFD0 U777 ( .I(n875), .Z(n876) );
  BUFFD0 U778 ( .I(n876), .Z(n877) );
  BUFFD0 U779 ( .I(n877), .Z(n878) );
  BUFFD0 U780 ( .I(n878), .Z(n879) );
  BUFFD0 U781 ( .I(n879), .Z(n880) );
  BUFFD0 U782 ( .I(n880), .Z(n881) );
  BUFFD0 U783 ( .I(n881), .Z(n882) );
  BUFFD0 U784 ( .I(n882), .Z(n883) );
  BUFFD0 U785 ( .I(n883), .Z(n884) );
  BUFFD0 U786 ( .I(n884), .Z(n885) );
  BUFFD0 U787 ( .I(n885), .Z(n886) );
  BUFFD0 U788 ( .I(n886), .Z(n887) );
  BUFFD0 U789 ( .I(n887), .Z(n888) );
  BUFFD0 U790 ( .I(n888), .Z(n889) );
  BUFFD0 U791 ( .I(n893), .Z(n890) );
  BUFFD0 U792 ( .I(N70), .Z(n891) );
  BUFFD0 U793 ( .I(n891), .Z(n892) );
  BUFFD0 U794 ( .I(n894), .Z(n893) );
  BUFFD0 U795 ( .I(n895), .Z(n894) );
  BUFFD0 U796 ( .I(n896), .Z(n895) );
  BUFFD0 U797 ( .I(n897), .Z(n896) );
  BUFFD0 U798 ( .I(n898), .Z(n897) );
  BUFFD0 U799 ( .I(n899), .Z(n898) );
  BUFFD0 U800 ( .I(n900), .Z(n899) );
  BUFFD0 U801 ( .I(n901), .Z(n900) );
  BUFFD0 U802 ( .I(n902), .Z(n901) );
  BUFFD0 U803 ( .I(n903), .Z(n902) );
  BUFFD0 U804 ( .I(n904), .Z(n903) );
  BUFFD0 U805 ( .I(n905), .Z(n904) );
  BUFFD0 U806 ( .I(n906), .Z(n905) );
  BUFFD0 U807 ( .I(n907), .Z(n906) );
  BUFFD0 U808 ( .I(n908), .Z(n907) );
  BUFFD0 U809 ( .I(n909), .Z(n908) );
  BUFFD0 U810 ( .I(n910), .Z(n909) );
  BUFFD0 U811 ( .I(n911), .Z(n910) );
  BUFFD0 U812 ( .I(n912), .Z(n911) );
  BUFFD0 U813 ( .I(n913), .Z(n912) );
  BUFFD0 U814 ( .I(n914), .Z(n913) );
  BUFFD0 U815 ( .I(n915), .Z(n914) );
  BUFFD0 U816 ( .I(n916), .Z(n915) );
  BUFFD0 U817 ( .I(n917), .Z(n916) );
  BUFFD0 U818 ( .I(n918), .Z(n917) );
  BUFFD0 U819 ( .I(n919), .Z(n918) );
  BUFFD0 U820 ( .I(n920), .Z(n919) );
  BUFFD0 U821 ( .I(n921), .Z(n920) );
  BUFFD0 U822 ( .I(n922), .Z(n921) );
  BUFFD0 U823 ( .I(n923), .Z(n922) );
  BUFFD0 U824 ( .I(n892), .Z(n923) );
  XNR2D0 U825 ( .A1(n126), .A2(WriteAddr[3]), .ZN(n99) );
  BUFFD0 U826 ( .I(n928), .Z(n925) );
  BUFFD0 U827 ( .I(N69), .Z(n926) );
  BUFFD0 U828 ( .I(n926), .Z(n927) );
  BUFFD0 U829 ( .I(n929), .Z(n928) );
  BUFFD0 U830 ( .I(n930), .Z(n929) );
  BUFFD0 U831 ( .I(n931), .Z(n930) );
  BUFFD0 U832 ( .I(n932), .Z(n931) );
  BUFFD0 U833 ( .I(n933), .Z(n932) );
  BUFFD0 U834 ( .I(n934), .Z(n933) );
  BUFFD0 U835 ( .I(n935), .Z(n934) );
  BUFFD0 U836 ( .I(n936), .Z(n935) );
  BUFFD0 U837 ( .I(n937), .Z(n936) );
  BUFFD0 U838 ( .I(n938), .Z(n937) );
  BUFFD0 U839 ( .I(n939), .Z(n938) );
  BUFFD0 U840 ( .I(n940), .Z(n939) );
  BUFFD0 U841 ( .I(n941), .Z(n940) );
  BUFFD0 U842 ( .I(n942), .Z(n941) );
  BUFFD0 U843 ( .I(n943), .Z(n942) );
  BUFFD0 U844 ( .I(n944), .Z(n943) );
  BUFFD0 U845 ( .I(n945), .Z(n944) );
  BUFFD0 U846 ( .I(n946), .Z(n945) );
  BUFFD0 U847 ( .I(n947), .Z(n946) );
  BUFFD0 U848 ( .I(n948), .Z(n947) );
  BUFFD0 U849 ( .I(n949), .Z(n948) );
  BUFFD0 U850 ( .I(n950), .Z(n949) );
  BUFFD0 U851 ( .I(n951), .Z(n950) );
  BUFFD0 U852 ( .I(n952), .Z(n951) );
  BUFFD0 U853 ( .I(n953), .Z(n952) );
  BUFFD0 U854 ( .I(n954), .Z(n953) );
  BUFFD0 U855 ( .I(n955), .Z(n954) );
  BUFFD0 U856 ( .I(n956), .Z(n955) );
  BUFFD0 U857 ( .I(n957), .Z(n956) );
  BUFFD0 U858 ( .I(n958), .Z(n957) );
  BUFFD0 U859 ( .I(n959), .Z(n958) );
  BUFFD0 U860 ( .I(n927), .Z(n959) );
  BUFFD0 U861 ( .I(n963), .Z(n960) );
  BUFFD0 U862 ( .I(N67), .Z(n961) );
  BUFFD0 U863 ( .I(n961), .Z(n962) );
  BUFFD0 U864 ( .I(n964), .Z(n963) );
  BUFFD0 U865 ( .I(n965), .Z(n964) );
  BUFFD0 U866 ( .I(n966), .Z(n965) );
  BUFFD0 U867 ( .I(n967), .Z(n966) );
  BUFFD0 U868 ( .I(n968), .Z(n967) );
  BUFFD0 U869 ( .I(n969), .Z(n968) );
  BUFFD0 U870 ( .I(n970), .Z(n969) );
  BUFFD0 U871 ( .I(n971), .Z(n970) );
  BUFFD0 U872 ( .I(n972), .Z(n971) );
  BUFFD0 U873 ( .I(n973), .Z(n972) );
  BUFFD0 U874 ( .I(n974), .Z(n973) );
  BUFFD0 U875 ( .I(n975), .Z(n974) );
  BUFFD0 U876 ( .I(n976), .Z(n975) );
  BUFFD0 U877 ( .I(n977), .Z(n976) );
  BUFFD0 U878 ( .I(n978), .Z(n977) );
  BUFFD0 U879 ( .I(n979), .Z(n978) );
  BUFFD0 U880 ( .I(n980), .Z(n979) );
  BUFFD0 U881 ( .I(n981), .Z(n980) );
  BUFFD0 U882 ( .I(n982), .Z(n981) );
  BUFFD0 U883 ( .I(n983), .Z(n982) );
  BUFFD0 U884 ( .I(n984), .Z(n983) );
  BUFFD0 U885 ( .I(n985), .Z(n984) );
  BUFFD0 U886 ( .I(n986), .Z(n985) );
  BUFFD0 U887 ( .I(n987), .Z(n986) );
  BUFFD0 U888 ( .I(n988), .Z(n987) );
  BUFFD0 U889 ( .I(n989), .Z(n988) );
  BUFFD0 U890 ( .I(n990), .Z(n989) );
  BUFFD0 U891 ( .I(n991), .Z(n990) );
  BUFFD0 U892 ( .I(n992), .Z(n991) );
  BUFFD0 U893 ( .I(n993), .Z(n992) );
  BUFFD0 U894 ( .I(n994), .Z(n993) );
  BUFFD0 U895 ( .I(n962), .Z(n994) );
  BUFFD0 U896 ( .I(n996), .Z(n995) );
  BUFFD0 U897 ( .I(n997), .Z(n996) );
  BUFFD0 U898 ( .I(n998), .Z(n997) );
  BUFFD0 U899 ( .I(n999), .Z(n998) );
  BUFFD0 U900 ( .I(n1000), .Z(n999) );
  BUFFD0 U901 ( .I(n1001), .Z(n1000) );
  BUFFD0 U902 ( .I(n1002), .Z(n1001) );
  BUFFD0 U903 ( .I(n1003), .Z(n1002) );
  BUFFD0 U904 ( .I(n1004), .Z(n1003) );
  BUFFD0 U905 ( .I(n1005), .Z(n1004) );
  BUFFD0 U906 ( .I(n1006), .Z(n1005) );
  BUFFD0 U907 ( .I(n1007), .Z(n1006) );
  BUFFD0 U908 ( .I(n1008), .Z(n1007) );
  BUFFD0 U909 ( .I(n1009), .Z(n1008) );
  BUFFD0 U910 ( .I(n1010), .Z(n1009) );
  BUFFD0 U911 ( .I(n1011), .Z(n1010) );
  BUFFD0 U912 ( .I(n1012), .Z(n1011) );
  BUFFD0 U913 ( .I(n1013), .Z(n1012) );
  BUFFD0 U914 ( .I(n1014), .Z(n1013) );
  BUFFD0 U915 ( .I(n1015), .Z(n1014) );
  BUFFD0 U916 ( .I(n1016), .Z(n1015) );
  BUFFD0 U917 ( .I(n1017), .Z(n1016) );
  BUFFD0 U918 ( .I(n1018), .Z(n1017) );
  BUFFD0 U919 ( .I(n1019), .Z(n1018) );
  BUFFD0 U920 ( .I(N71), .Z(n1019) );
  ND3D0 U921 ( .A1(n171), .A2(n170), .A3(n172), .ZN(n35) );
  INVD0 U922 ( .I(n53), .ZN(n42) );
  BUFFD0 U923 ( .I(n889), .Z(n1020) );
  INVD1 U924 ( .I(Reset), .ZN(n1033) );
  INVD1 U925 ( .I(Reset), .ZN(n1032) );
  INVD1 U926 ( .I(n48), .ZN(n49) );
  ND2D1 U927 ( .A1(n66), .A2(n42), .ZN(n119) );
  OAI211D1 U928 ( .A1(n35), .A2(n63), .B(n66), .C(n115), .ZN(n48) );
  INR2D1 U929 ( .A1(n71), .B1(n116), .ZN(n115) );
  AOI21D1 U930 ( .A1(n52), .A2(n117), .B(n170), .ZN(n116) );
  MAOI22D0 U931 ( .A1(n5), .A2(n170), .B1(n170), .B2(n71), .ZN(n66) );
  ND2D1 U932 ( .A1(n66), .A2(n35), .ZN(n47) );
  INVD1 U933 ( .I(n106), .ZN(n76) );
  OA211D0 U934 ( .A1(n75), .A2(n76), .B(n77), .C(n78), .Z(n55) );
  INVD1 U935 ( .I(n85), .ZN(n77) );
  NR3D0 U936 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n78) );
  NR3D0 U937 ( .A1(WriteAddr[2]), .A2(n46), .A3(ReadAddr[2]), .ZN(n80) );
  ND2D1 U938 ( .A1(n130), .A2(n806), .ZN(n129) );
  INVD1 U939 ( .I(n40), .ZN(n38) );
  ND2D1 U940 ( .A1(n107), .A2(n108), .ZN(n85) );
  XNR2D1 U941 ( .A1(ReadAddr[1]), .A2(n46), .ZN(n107) );
  INVD1 U942 ( .I(n90), .ZN(n84) );
  INVD1 U943 ( .I(n97), .ZN(n108) );
  AOI21D1 U944 ( .A1(n76), .A2(n83), .B(ReadAddr[1]), .ZN(n105) );
  NR3D0 U945 ( .A1(n117), .A2(n124), .A3(n125), .ZN(n123) );
  XNR2D1 U946 ( .A1(ReadAddr[3]), .A2(n670), .ZN(n125) );
  XNR2D1 U947 ( .A1(ReadAddr[2]), .A2(n671), .ZN(n124) );
  XNR2D1 U948 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n104) );
  NR2D1 U949 ( .A1(n114), .A2(n118), .ZN(N49) );
  NR2D1 U950 ( .A1(n808), .A2(n118), .ZN(N48) );
  NR2D1 U951 ( .A1(n746), .A2(n118), .ZN(N51) );
  NR2D1 U952 ( .A1(n838), .A2(n118), .ZN(N47) );
  ND2D1 U953 ( .A1(WriteReq), .A2(n47), .ZN(n45) );
  OAI32D1 U954 ( .A1(n35), .A2(WriteReq), .A3(Reset), .B1(n36), .B2(n7), .ZN(
        n147) );
  AOI21D1 U955 ( .A1(n37), .A2(n35), .B(Reset), .ZN(n36) );
  OAI22D0 U956 ( .A1(n48), .A2(n456), .B1(n49), .B2(n50), .ZN(n156) );
  AOI21D1 U957 ( .A1(n51), .A2(n52), .B(n53), .ZN(n50) );
  OAI22D0 U958 ( .A1(n171), .A2(n54), .B1(n170), .B2(n55), .ZN(n51) );
  OAI22D0 U959 ( .A1(n48), .A2(n420), .B1(n49), .B2(n67), .ZN(n158) );
  AOI31D0 U960 ( .A1(n68), .A2(n5), .A3(n170), .B(n70), .ZN(n67) );
  IOA21D1 U961 ( .A1(n52), .A2(n54), .B(n86), .ZN(n68) );
  OAI31D0 U962 ( .A1(n71), .A2(n170), .A3(n72), .B(n35), .ZN(n70) );
  OAI22D0 U963 ( .A1(n48), .A2(n384), .B1(n49), .B2(n100), .ZN(n159) );
  AOI22D0 U964 ( .A1(n101), .A2(n52), .B1(n102), .B2(n103), .ZN(n100) );
  AOI211D1 U965 ( .A1(n164), .A2(n106), .B(n37), .C(n85), .ZN(n102) );
  AOI221D0 U966 ( .A1(n90), .A2(n76), .B1(n104), .B2(ReadAddr[1]), .C(n105), 
        .ZN(n103) );
  NR3D0 U967 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n60) );
  XNR2D1 U968 ( .A1(n167), .A2(n492), .ZN(n62) );
  XNR2D1 U969 ( .A1(n46), .A2(n494), .ZN(n61) );
  XNR2D1 U970 ( .A1(WriteAddr[0]), .A2(n495), .ZN(n58) );
  XNR2D1 U971 ( .A1(WriteAddr[2]), .A2(n491), .ZN(n59) );
  INVD1 U972 ( .I(WriteReq), .ZN(n63) );
  CKND2D0 U973 ( .A1(ReadReq), .A2(n119), .ZN(n40) );
  ND2D1 U974 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .ZN(n128) );
  AOI21D1 U975 ( .A1(n128), .A2(n168), .B(n126), .ZN(n98) );
  ND2D1 U976 ( .A1(n171), .A2(n52), .ZN(n71) );
  OAI22D0 U977 ( .A1(n38), .A2(n671), .B1(n164), .B2(n40), .ZN(n148) );
  OAI22D0 U978 ( .A1(n38), .A2(n670), .B1(n163), .B2(n40), .ZN(n150) );
  AOI21D1 U979 ( .A1(n83), .A2(n84), .B(WriteAddr[1]), .ZN(n79) );
  NR2D1 U980 ( .A1(WriteAddr[2]), .A2(n164), .ZN(n90) );
  OAI21D1 U981 ( .A1(n171), .A2(n109), .B(n170), .ZN(n101) );
  NR4D0 U982 ( .A1(n108), .A2(n110), .A3(n95), .A4(n111), .ZN(n109) );
  XNR2D1 U983 ( .A1(WriteAddr[2]), .A2(n114), .ZN(n110) );
  XNR2D1 U984 ( .A1(WriteAddr[3]), .A2(n112), .ZN(n111) );
  ND4D1 U985 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(n54) );
  XNR2D1 U986 ( .A1(n99), .A2(n163), .ZN(n94) );
  XNR2D1 U987 ( .A1(ReadAddr[2]), .A2(n98), .ZN(n96) );
  NR2D1 U988 ( .A1(n128), .A2(n168), .ZN(n126) );
  NR2D1 U989 ( .A1(n46), .A2(n168), .ZN(n75) );
  XNR2D1 U990 ( .A1(ReadAddr[3]), .A2(n167), .ZN(n106) );
  XNR2D1 U991 ( .A1(WriteAddr[0]), .A2(n166), .ZN(n97) );
  ND2D1 U992 ( .A1(WriteCmd), .A2(n42), .ZN(n56) );
  OAI211D1 U993 ( .A1(n46), .A2(ReadAddr[1]), .B(n83), .C(n92), .ZN(n74) );
  AOI22D0 U994 ( .A1(n163), .A2(WriteAddr[3]), .B1(n166), .B2(WriteAddr[0]), 
        .ZN(n92) );
  OAI21D1 U995 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n128), .ZN(n113) );
  OAI211D1 U996 ( .A1(n165), .A2(WriteAddr[1]), .B(n84), .C(n87), .ZN(n73) );
  AOI22D0 U997 ( .A1(n167), .A2(ReadAddr[3]), .B1(n169), .B2(ReadAddr[0]), 
        .ZN(n87) );
  OAI22D0 U998 ( .A1(n165), .A2(n42), .B1(n113), .B2(n56), .ZN(N68) );
  OAI22D0 U999 ( .A1(n924), .A2(n42), .B1(n99), .B2(n56), .ZN(N70) );
  OAI22D0 U1000 ( .A1(n164), .A2(n42), .B1(n127), .B2(n56), .ZN(N69) );
  INVD1 U1001 ( .I(n98), .ZN(n127) );
  OAI22D0 U1002 ( .A1(n166), .A2(n42), .B1(WriteAddr[0]), .B2(n56), .ZN(N67)
         );
  NR3D0 U1003 ( .A1(n171), .A2(n172), .A3(n170), .ZN(n53) );
  ND2D1 U1004 ( .A1(n164), .A2(WriteAddr[2]), .ZN(n83) );
  ND3D1 U1005 ( .A1(n170), .A2(n5), .A3(n172), .ZN(n37) );
  XNR2D1 U1006 ( .A1(ReadAddr[0]), .A2(n668), .ZN(n121) );
  XNR2D1 U1007 ( .A1(ReadAddr[1]), .A2(n667), .ZN(n122) );
  OAI21D1 U1008 ( .A1(n74), .A2(n73), .B(n172), .ZN(n86) );
  NR2D1 U1009 ( .A1(n166), .A2(n165), .ZN(n130) );
  XNR2D1 U1010 ( .A1(n113), .A2(n165), .ZN(n95) );
  OAI31D0 U1011 ( .A1(n42), .A2(Reset), .A3(ReadReq), .B(n138), .ZN(n151) );
  INVD1 U1012 ( .I(n666), .ZN(n39) );
  INVD1 U1013 ( .I(n665), .ZN(n41) );
  ND2D1 U1014 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  INVD0 U1015 ( .I(ReadReq), .ZN(n117) );
endmodule


module DPMem1kx32_AWid4_DWid32_0 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [3:0] AddrR;
  input [3:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N9, N44, N45, N46, N47, ClockR, ClockW, Dreadyr, \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N84, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n103, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n85, n102, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];

  XNR4D1 U13 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n76) );
  XOR4D1 U14 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n75) );
  XOR4D1 U15 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n72) );
  XOR4D1 U16 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n69) );
  XNR4D1 U17 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n66) );
  XOR4D1 U21 ( .A1(n81), .A2(n4002), .A3(n82), .A4(n4001), .Z(n80) );
  XNR4D1 U22 ( .A1(n3965), .A2(n3971), .A3(n3963), .A4(n3961), .ZN(n82) );
  XNR4D1 U27 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n88) );
  XOR4D1 U28 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n87) );
  XNR4D1 U29 ( .A1(n3924), .A2(n3932), .A3(n3935), .A4(n3931), .ZN(n84) );
  XNR4D1 U30 ( .A1(n4006), .A2(n4008), .A3(n4007), .A4(n4004), .ZN(n78) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N84), .E(n4248), .CP(n4284), .CDN(n4349), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(n4248), .CP(n4284), .CDN(
        n4356), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(n4249), .CP(n4284), .CDN(
        n4348), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(DataI[29]), .E(n4248), .CP(n4285), .CDN(
        n4358), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(n4249), .CP(n4285), .CDN(
        n4352), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(n4248), .CP(n4285), .CDN(
        n4339), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(DataI[22]), .E(n4248), .CP(n4285), .CDN(
        n4358), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(n4248), .CP(n4285), .CDN(
        n4351), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(DataI[20]), .E(n4248), .CP(n4286), .CDN(
        n4360), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(n4248), .CP(n4286), .CDN(
        n4357), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(n4248), .CP(n4286), .CDN(
        n4358), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(DataI[17]), .E(n4248), .CP(n4286), .CDN(
        n4354), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(n4248), .CP(n4286), .CDN(
        n4356), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(DataI[15]), .E(n4248), .CP(n4286), .CDN(
        n4354), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(n4248), .CP(n4286), .CDN(
        n4352), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(n4248), .CP(n4286), .CDN(
        n4358), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(DataI[12]), .E(n4249), .CP(n4286), .CDN(
        n4362), .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(n4249), .CP(n4287), .CDN(
        n4353), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(DataI[10]), .E(n4249), .CP(n4287), .CDN(
        n4361), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(DataI[9]), .E(n4249), .CP(n4287), .CDN(
        n4340), .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(n4249), .CP(n4287), .CDN(
        n4354), .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(DataI[7]), .E(n4249), .CP(n4287), .CDN(
        n4356), .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(DataI[6]), .E(n4249), .CP(n4287), .CDN(
        n4355), .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(DataI[5]), .E(n4249), .CP(n4287), .CDN(
        n4356), .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(DataI[4]), .E(n4249), .CP(n4287), .CDN(
        n4357), .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(DataI[3]), .E(n4249), .CP(n4287), .CDN(
        n4361), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(DataI[2]), .E(n4249), .CP(n4288), .CDN(
        n4360), .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(DataI[1]), .E(n4249), .CP(n4288), .CDN(
        n4335), .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(DataI[0]), .E(n4248), .CP(n4288), .CDN(
        n4359), .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N84), .E(n4250), .CP(n4288), .CDN(n4346), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(DataI[31]), .E(n4250), .CP(n4288), .CDN(
        n4347), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(DataI[30]), .E(n4251), .CP(n4288), .CDN(
        n4360), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(n4250), .CP(n4288), .CDN(
        n4363), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(DataI[24]), .E(n4251), .CP(n4289), .CDN(
        n4350), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(DataI[23]), .E(n4250), .CP(n4289), .CDN(
        n4353), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(DataI[22]), .E(n4250), .CP(n4289), .CDN(
        n4351), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(DataI[21]), .E(n4250), .CP(n4289), .CDN(
        n4356), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(n4250), .CP(n4289), .CDN(
        n4362), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(DataI[19]), .E(n4250), .CP(n4289), .CDN(
        n4361), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(DataI[18]), .E(n4250), .CP(n4289), .CDN(
        n4358), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(n4250), .CP(n4290), .CDN(
        n4351), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(DataI[16]), .E(n4250), .CP(n4290), .CDN(
        n4357), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(n4250), .CP(n4290), .CDN(
        n4335), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(DataI[14]), .E(n4250), .CP(n4290), .CDN(
        n4350), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(DataI[13]), .E(n4250), .CP(n4290), .CDN(
        n4351), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(DataI[12]), .E(n4251), .CP(n4290), .CDN(
        n4352), .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(DataI[11]), .E(n4251), .CP(n4290), .CDN(
        n4360), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(n4251), .CP(n4290), .CDN(
        n4357), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(DataI[9]), .E(n4251), .CP(n4290), .CDN(
        n4345), .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(DataI[8]), .E(n4251), .CP(n4291), .CDN(
        n4360), .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(n4251), .CP(n4291), .CDN(
        n4361), .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(DataI[6]), .E(n4251), .CP(n4291), .CDN(
        n4363), .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(DataI[5]), .E(n4251), .CP(n4291), .CDN(
        n4354), .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(DataI[4]), .E(n4251), .CP(n4291), .CDN(
        n4353), .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(n4251), .CP(n4291), .CDN(
        n4362), .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(DataI[2]), .E(n4251), .CP(n4291), .CDN(
        n4362), .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(n4250), .CP(n4291), .CDN(
        n4347), .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(DataI[0]), .E(n4251), .CP(n4291), .CDN(
        n4363), .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N84), .E(n4256), .CP(n4299), .CDN(n4353), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(DataI[31]), .E(n4256), .CP(n4299), .CDN(
        n4359), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(DataI[30]), .E(n4257), .CP(n4299), .CDN(
        n4350), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(DataI[29]), .E(n4256), .CP(n4299), .CDN(
        n4354), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(DataI[24]), .E(n4257), .CP(n4300), .CDN(
        n4353), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(DataI[23]), .E(n4256), .CP(n4300), .CDN(
        n4359), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(DataI[22]), .E(n4256), .CP(n4300), .CDN(
        n4363), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(DataI[21]), .E(n4256), .CP(n4300), .CDN(
        n4355), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(DataI[20]), .E(n4256), .CP(n4300), .CDN(
        n4357), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(DataI[19]), .E(n4256), .CP(n4300), .CDN(
        n4356), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(DataI[18]), .E(n4256), .CP(n4300), .CDN(
        n4349), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(DataI[17]), .E(n4256), .CP(n4301), .CDN(
        n4355), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(DataI[16]), .E(n4256), .CP(n4301), .CDN(
        n4355), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(DataI[15]), .E(n4256), .CP(n4301), .CDN(
        n4361), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(DataI[14]), .E(n4256), .CP(n4301), .CDN(
        n4334), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(DataI[13]), .E(n4256), .CP(n4301), .CDN(
        n4342), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(DataI[12]), .E(n4257), .CP(n4301), .CDN(
        n4356), .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(DataI[11]), .E(n4257), .CP(n4301), .CDN(
        n4335), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(DataI[10]), .E(n4257), .CP(n4301), .CDN(
        n4358), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(DataI[9]), .E(n4257), .CP(n4301), .CDN(
        n4360), .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(DataI[8]), .E(n4257), .CP(n4302), .CDN(
        n4358), .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(DataI[7]), .E(n4257), .CP(n4302), .CDN(
        n4355), .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(DataI[6]), .E(n4257), .CP(n4302), .CDN(
        n4354), .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(DataI[5]), .E(n4257), .CP(n4302), .CDN(
        n4357), .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(DataI[4]), .E(n4257), .CP(n4302), .CDN(
        n4362), .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(DataI[3]), .E(n4257), .CP(n4302), .CDN(
        n4344), .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(DataI[2]), .E(n4257), .CP(n4302), .CDN(
        n4363), .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(DataI[1]), .E(n4256), .CP(n4302), .CDN(
        n4354), .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(DataI[0]), .E(n4257), .CP(n4302), .CDN(
        n4353), .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N84), .E(n4258), .CP(n4303), .CDN(n4355), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(DataI[31]), .E(n4258), .CP(n4310), .CDN(
        n4349), .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(DataI[30]), .E(n4258), .CP(n4307), .CDN(
        n4349), .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(DataI[29]), .E(n4258), .CP(n4286), .CDN(
        n4349), .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(DataI[24]), .E(n4258), .CP(n4287), .CDN(
        n4349), .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(DataI[23]), .E(n4258), .CP(n4303), .CDN(
        n4349), .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(n4259), .CP(n4303), .CDN(
        n4349), .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(DataI[21]), .E(n4259), .CP(n4303), .CDN(
        n4349), .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(DataI[20]), .E(n4259), .CP(n4303), .CDN(
        n4348), .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(DataI[19]), .E(n4259), .CP(n4303), .CDN(
        n4348), .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(DataI[18]), .E(n4259), .CP(n4303), .CDN(
        n4348), .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(DataI[17]), .E(n4259), .CP(n4303), .CDN(
        n4348), .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(DataI[16]), .E(n4259), .CP(n4303), .CDN(
        n4348), .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(DataI[15]), .E(n4259), .CP(n4303), .CDN(
        n4348), .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(DataI[14]), .E(n4259), .CP(n4304), .CDN(
        n4348), .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(DataI[13]), .E(n4259), .CP(n4304), .CDN(
        n4348), .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(n4258), .CP(n4304), .CDN(
        n4348), .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(DataI[11]), .E(n4259), .CP(n4304), .CDN(
        n4348), .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(DataI[10]), .E(n4258), .CP(n4304), .CDN(
        n4348), .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(n4259), .CP(n4304), .CDN(
        n4347), .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(DataI[8]), .E(n4258), .CP(n4304), .CDN(
        n4347), .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(DataI[7]), .E(n4259), .CP(n4304), .CDN(
        n4347), .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(DataI[6]), .E(n4258), .CP(n4304), .CDN(
        n4347), .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(DataI[5]), .E(n4259), .CP(n4305), .CDN(
        n4347), .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(n4258), .CP(n4305), .CDN(
        n4347), .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(DataI[3]), .E(n4259), .CP(n4305), .CDN(
        n4347), .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(DataI[2]), .E(n4259), .CP(n4305), .CDN(
        n4347), .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(DataI[1]), .E(n4259), .CP(n4305), .CDN(
        n4347), .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(n4258), .CP(n4305), .CDN(
        n4347), .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N84), .E(n4264), .CP(n4285), .CDN(n4343), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(n4264), .CP(n4281), .CDN(
        n4342), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(n4265), .CP(n4283), .CDN(
        n4342), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n4264), .CP(n4282), .CDN(
        n4342), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n4265), .CP(ClockW), .CDN(
        n4342), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n4264), .CP(n4310), .CDN(
        n4342), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n4264), .CP(n4281), .CDN(
        n4342), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(n4264), .CP(n4321), .CDN(
        n4342), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n4264), .CP(n4322), .CDN(
        n4341), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n4264), .CP(n4314), .CDN(
        n4341), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n4264), .CP(n4317), .CDN(
        n4341), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n4264), .CP(n4323), .CDN(
        n4341), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n4264), .CP(n4324), .CDN(
        n4341), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n4264), .CP(n4325), .CDN(
        n4341), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(n4264), .CP(n4320), .CDN(
        n4341), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(n4264), .CP(n4322), .CDN(
        n4341), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n4265), .CP(n4308), .CDN(
        n4341), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n4265), .CP(n4309), .CDN(
        n4341), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n4265), .CP(n4310), .CDN(
        n4341), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n4265), .CP(n4279), .CDN(
        n4340), .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(n4265), .CP(n4322), .CDN(
        n4340), .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(n4265), .CP(n4324), .CDN(
        n4340), .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(n4265), .CP(n4325), .CDN(
        n4340), .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(n4265), .CP(n4310), .CDN(
        n4340), .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n4265), .CP(n4312), .CDN(
        n4340), .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n4265), .CP(n4324), .CDN(
        n4340), .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n4265), .CP(n4319), .CDN(
        n4340), .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n4265), .CP(ClockW), .CDN(
        n4340), .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n4264), .CP(n4280), .CDN(
        n4340), .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N84), .E(n4266), .CP(n4297), .CDN(n4340), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(n4266), .CP(n4278), .CDN(
        n4351), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(n4267), .CP(n4291), .CDN(
        n4358), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(n4266), .CP(n4287), .CDN(
        n4339), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n4267), .CP(n4309), .CDN(
        n4344), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(n4266), .CP(n4308), .CDN(
        n4357), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n4266), .CP(n4320), .CDN(
        n4352), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(n4266), .CP(n4321), .CDN(
        n4347), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n4266), .CP(n4282), .CDN(
        n4360), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n4266), .CP(n4292), .CDN(
        n4339), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n4266), .CP(n4290), .CDN(
        n4352), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n4266), .CP(n4291), .CDN(
        n4363), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n4266), .CP(n4279), .CDN(
        n4363), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n4266), .CP(n4283), .CDN(
        n4363), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(n4266), .CP(n4284), .CDN(
        n4348), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n4266), .CP(n4285), .CDN(
        n4350), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n4267), .CP(n4283), .CDN(
        n4355), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n4267), .CP(n4317), .CDN(
        n4351), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n4267), .CP(n4279), .CDN(
        n4361), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n4267), .CP(n4316), .CDN(
        n4346), .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(n4267), .CP(n4310), .CDN(
        n4361), .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(n4267), .CP(n4292), .CDN(
        n4361), .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n4267), .CP(n4320), .CDN(
        n4334), .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(n4267), .CP(n4278), .CDN(
        n4347), .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n4267), .CP(ClockW), .CDN(
        n4339), .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n4267), .CP(n4321), .CDN(
        n4349), .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n4267), .CP(n4323), .CDN(
        n4338), .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(n4267), .CP(n4311), .CDN(
        n4338), .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n4266), .CP(n4310), .CDN(
        n4345), .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N84), .E(n4272), .CP(n4312), .CDN(n4351), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(n4272), .CP(n4316), .CDN(
        n4343), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(n4273), .CP(n4319), .CDN(
        n4355), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(n4272), .CP(n4315), .CDN(
        n4350), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n4273), .CP(n4319), .CDN(
        n4346), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(n4272), .CP(n4320), .CDN(
        n4349), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n4272), .CP(n4279), .CDN(
        n4341), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n4272), .CP(n4312), .CDN(
        n4347), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n4272), .CP(n4311), .CDN(
        n4341), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n4272), .CP(n4313), .CDN(
        n4345), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n4272), .CP(n4278), .CDN(
        n4351), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n4272), .CP(n4278), .CDN(
        n4363), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n4272), .CP(n4280), .CDN(
        n4341), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(n4272), .CP(n4278), .CDN(
        n4336), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n4272), .CP(n4315), .CDN(
        n4337), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n4272), .CP(n4314), .CDN(
        n4356), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n4273), .CP(n4313), .CDN(
        n4335), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n4273), .CP(n4308), .CDN(
        n4357), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n4273), .CP(n4315), .CDN(
        n4358), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n4273), .CP(n4321), .CDN(
        n4350), .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n4273), .CP(n4320), .CDN(
        n4359), .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(n4273), .CP(n4312), .CDN(
        n4353), .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n4273), .CP(n4297), .CDN(
        n4348), .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(n4273), .CP(n4314), .CDN(
        n4354), .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n4273), .CP(n4318), .CDN(
        n4342), .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(n4273), .CP(n4309), .CDN(
        n4341), .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n4273), .CP(n4314), .CDN(
        n4340), .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(n4273), .CP(n4318), .CDN(
        n4348), .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(n4272), .CP(n4324), .CDN(
        n4342), .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N84), .E(n4274), .CP(n4279), .CDN(n4343), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(n4274), .CP(n4320), .CDN(
        n4339), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(n4275), .CP(n4312), .CDN(
        n4339), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(n4274), .CP(n4311), .CDN(
        n4339), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n4275), .CP(n4317), .CDN(
        n4339), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n4274), .CP(n4316), .CDN(
        n4339), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n4274), .CP(n4323), .CDN(
        n4339), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(n4274), .CP(n4315), .CDN(
        n4339), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n4274), .CP(n4295), .CDN(
        n4338), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n4274), .CP(n4316), .CDN(
        n4338), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n4274), .CP(n4317), .CDN(
        n4338), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n4274), .CP(n4294), .CDN(
        n4338), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n4274), .CP(n4309), .CDN(
        n4338), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n4274), .CP(n4308), .CDN(
        n4338), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(n4274), .CP(n4304), .CDN(
        n4338), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(n4274), .CP(n4295), .CDN(
        n4338), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n4275), .CP(n4280), .CDN(
        n4338), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n4275), .CP(n4323), .CDN(
        n4338), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n4275), .CP(n4325), .CDN(
        n4338), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n4275), .CP(n4318), .CDN(
        n4337), .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(n4275), .CP(n4321), .CDN(
        n4337), .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(n4275), .CP(n4321), .CDN(
        n4337), .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(n4275), .CP(n4307), .CDN(
        n4337), .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(n4275), .CP(n4318), .CDN(
        n4337), .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n4275), .CP(n4314), .CDN(
        n4337), .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n4275), .CP(n4310), .CDN(
        n4337), .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n4275), .CP(n4317), .CDN(
        n4337), .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n4275), .CP(ClockW), .CDN(
        n4337), .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n4274), .CP(n4305), .CDN(
        n4337), .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N84), .E(n4246), .CP(n4281), .CDN(n4356), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(n4246), .CP(n4281), .CDN(
        n4359), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(n4247), .CP(n4281), .CDN(
        n4362), .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(DataI[29]), .E(n4247), .CP(n4281), .CDN(
        n4353), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(n4247), .CP(n4281), .CDN(
        n4359), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(n4247), .CP(n4282), .CDN(
        n4354), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(DataI[22]), .E(n4246), .CP(n4282), .CDN(
        n4354), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(n4246), .CP(n4282), .CDN(
        n4351), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(DataI[20]), .E(n4246), .CP(n4282), .CDN(
        n4337), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(n4246), .CP(n4282), .CDN(
        n4336), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(n4246), .CP(n4282), .CDN(
        n4338), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(DataI[17]), .E(n4246), .CP(n4282), .CDN(
        n4339), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(n4246), .CP(n4282), .CDN(
        n4355), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(DataI[15]), .E(n4246), .CP(n4282), .CDN(
        n4356), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(n4246), .CP(n4283), .CDN(
        n4360), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(n4246), .CP(n4283), .CDN(
        n4350), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(DataI[12]), .E(n4247), .CP(n4283), .CDN(
        n4343), .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(n4247), .CP(n4283), .CDN(
        n4354), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(DataI[10]), .E(n4247), .CP(n4283), .CDN(
        n4349), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(DataI[9]), .E(n4247), .CP(n4283), .CDN(
        n4342), .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(n4247), .CP(n4283), .CDN(
        n4335), .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(DataI[7]), .E(n4247), .CP(n4283), .CDN(
        n4355), .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(DataI[6]), .E(n4247), .CP(n4283), .CDN(
        n4353), .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(DataI[5]), .E(n4247), .CP(n4284), .CDN(
        n4363), .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(DataI[4]), .E(n4247), .CP(n4284), .CDN(
        n4344), .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(DataI[3]), .E(n4247), .CP(n4284), .CDN(
        n4362), .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(DataI[2]), .E(n4246), .CP(n4284), .CDN(
        n4350), .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(DataI[1]), .E(n4247), .CP(n4284), .CDN(
        n4362), .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(DataI[0]), .E(n4246), .CP(n4284), .CDN(
        n4355), .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N84), .E(n4252), .CP(n4292), .CDN(n4363), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(DataI[31]), .E(n4252), .CP(n4292), .CDN(
        n4363), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(DataI[30]), .E(n4253), .CP(n4292), .CDN(
        n4336), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(DataI[29]), .E(n4252), .CP(n4292), .CDN(
        n4359), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(DataI[24]), .E(n4253), .CP(n4292), .CDN(
        n4361), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(DataI[23]), .E(n4252), .CP(n4293), .CDN(
        n4362), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(DataI[22]), .E(n4252), .CP(n4293), .CDN(
        n4358), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(DataI[21]), .E(n4252), .CP(n4293), .CDN(
        n4357), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(DataI[20]), .E(n4252), .CP(n4293), .CDN(
        n4352), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(DataI[19]), .E(n4252), .CP(n4293), .CDN(
        n4355), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(DataI[18]), .E(n4252), .CP(n4293), .CDN(
        n4360), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(DataI[17]), .E(n4252), .CP(n4293), .CDN(
        n4359), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(DataI[16]), .E(n4252), .CP(n4293), .CDN(
        n4351), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(DataI[15]), .E(n4252), .CP(n4293), .CDN(
        n4334), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(DataI[14]), .E(n4252), .CP(n4294), .CDN(
        n4355), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(DataI[13]), .E(n4252), .CP(n4294), .CDN(
        n4360), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(DataI[12]), .E(n4253), .CP(n4294), .CDN(
        n4356), .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(DataI[11]), .E(n4253), .CP(n4294), .CDN(
        n4355), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(DataI[10]), .E(n4253), .CP(n4294), .CDN(
        n4356), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(DataI[9]), .E(n4253), .CP(n4294), .CDN(
        n4355), .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(DataI[8]), .E(n4253), .CP(n4294), .CDN(
        n4356), .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(DataI[7]), .E(n4253), .CP(n4294), .CDN(
        n4362), .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(DataI[6]), .E(n4253), .CP(n4294), .CDN(
        n4353), .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(DataI[5]), .E(n4253), .CP(n4295), .CDN(
        n4362), .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(DataI[4]), .E(n4253), .CP(n4295), .CDN(
        n4358), .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(DataI[3]), .E(n4253), .CP(n4295), .CDN(
        n4361), .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(DataI[2]), .E(n4253), .CP(n4295), .CDN(
        n4352), .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(DataI[1]), .E(n4252), .CP(n4295), .CDN(
        n4359), .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(DataI[0]), .E(n4253), .CP(n4295), .CDN(
        n4343), .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N84), .E(n4254), .CP(n4295), .CDN(n4350), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(DataI[31]), .E(n4254), .CP(n4295), .CDN(
        n4360), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(DataI[30]), .E(n4255), .CP(n4295), .CDN(
        n4335), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(DataI[29]), .E(n4254), .CP(n4296), .CDN(
        n4357), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(DataI[24]), .E(n4255), .CP(n4296), .CDN(
        n4358), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(DataI[23]), .E(n4254), .CP(n4296), .CDN(
        n4346), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(DataI[22]), .E(n4254), .CP(n4296), .CDN(
        n4353), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(DataI[21]), .E(n4254), .CP(n4296), .CDN(
        n4354), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(DataI[20]), .E(n4254), .CP(n4297), .CDN(
        n4334), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(DataI[19]), .E(n4254), .CP(n4297), .CDN(
        n4357), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(DataI[18]), .E(n4254), .CP(n4297), .CDN(
        n4363), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(DataI[17]), .E(n4254), .CP(n4297), .CDN(
        n4338), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(DataI[16]), .E(n4254), .CP(n4297), .CDN(
        n4341), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(DataI[15]), .E(n4254), .CP(n4297), .CDN(
        n4359), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(DataI[14]), .E(n4254), .CP(n4297), .CDN(
        n4359), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(DataI[13]), .E(n4254), .CP(n4297), .CDN(
        n4354), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(DataI[12]), .E(n4255), .CP(n4297), .CDN(
        n4353), .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(DataI[11]), .E(n4255), .CP(n4298), .CDN(
        n4362), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(DataI[10]), .E(n4255), .CP(n4298), .CDN(
        n4358), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(DataI[9]), .E(n4255), .CP(n4298), .CDN(
        n4351), .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(DataI[8]), .E(n4255), .CP(n4298), .CDN(
        n4363), .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(DataI[7]), .E(n4255), .CP(n4298), .CDN(
        n4338), .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(DataI[6]), .E(n4255), .CP(n4298), .CDN(
        n4356), .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(DataI[5]), .E(n4255), .CP(n4298), .CDN(
        n4337), .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(DataI[4]), .E(n4255), .CP(n4298), .CDN(
        n4344), .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(DataI[3]), .E(n4255), .CP(n4298), .CDN(
        n4348), .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(DataI[2]), .E(n4255), .CP(n4299), .CDN(
        n4338), .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(DataI[1]), .E(n4254), .CP(n4299), .CDN(
        n4359), .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(DataI[0]), .E(n4255), .CP(n4299), .CDN(
        n4352), .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N84), .E(n4260), .CP(n4305), .CDN(n4347), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(DataI[31]), .E(n4260), .CP(n4305), .CDN(
        n4346), .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(DataI[30]), .E(n4261), .CP(n4305), .CDN(
        n4346), .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(DataI[29]), .E(n4260), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(DataI[24]), .E(n4261), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(DataI[23]), .E(n4260), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(n4260), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(DataI[21]), .E(n4260), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(DataI[20]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(DataI[19]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(DataI[18]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(DataI[17]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(DataI[16]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(DataI[15]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(DataI[14]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(DataI[13]), .E(n4260), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(n4261), .CP(n4307), .CDN(
        n4345), .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(DataI[11]), .E(n4261), .CP(n4303), .CDN(
        n4345), .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(DataI[10]), .E(n4261), .CP(n4280), .CDN(
        n4345), .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(n4261), .CP(n4293), .CDN(
        n4344), .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(DataI[8]), .E(n4261), .CP(n4298), .CDN(
        n4344), .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(DataI[7]), .E(n4261), .CP(n4299), .CDN(
        n4344), .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(DataI[6]), .E(n4261), .CP(n4300), .CDN(
        n4344), .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(DataI[5]), .E(n4261), .CP(n4301), .CDN(
        n4344), .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(n4261), .CP(n4302), .CDN(
        n4344), .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(DataI[3]), .E(n4261), .CP(n4290), .CDN(
        n4344), .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(DataI[2]), .E(n4261), .CP(n4321), .CDN(
        n4344), .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(DataI[1]), .E(n4261), .CP(n4313), .CDN(
        n4344), .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(n4260), .CP(n4314), .CDN(
        n4344), .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N84), .E(n4262), .CP(n4311), .CDN(n4344), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(n4262), .CP(n4315), .CDN(
        n4343), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(n4263), .CP(n4309), .CDN(
        n4343), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n4262), .CP(n4312), .CDN(
        n4343), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(n4263), .CP(n4296), .CDN(
        n4343), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(n4262), .CP(n4305), .CDN(
        n4343), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n4262), .CP(n4284), .CDN(
        n4343), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(n4262), .CP(n4291), .CDN(
        n4343), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n4262), .CP(n4302), .CDN(
        n4343), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n4262), .CP(n4298), .CDN(
        n4341), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n4262), .CP(n4299), .CDN(
        n4342), .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n4262), .CP(n4285), .CDN(
        n4340), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(n4262), .CP(n4319), .CDN(
        n4343), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(n4262), .CP(n4306), .CDN(
        n4341), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(n4262), .CP(n4288), .CDN(
        n4342), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(n4262), .CP(n4289), .CDN(
        n4340), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n4263), .CP(n4286), .CDN(
        n4353), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n4263), .CP(n4287), .CDN(
        n4354), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n4263), .CP(n4281), .CDN(
        n4353), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n4263), .CP(n4282), .CDN(
        n4345), .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(n4263), .CP(n4317), .CDN(
        n4346), .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(n4263), .CP(n4284), .CDN(
        n4347), .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(n4263), .CP(n4307), .CDN(
        n4348), .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(n4263), .CP(n4312), .CDN(
        n4349), .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n4263), .CP(n4319), .CDN(
        n4336), .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n4263), .CP(n4322), .CDN(
        n4337), .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n4263), .CP(n4324), .CDN(
        n4357), .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(n4263), .CP(n4323), .CDN(
        n4345), .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(n4262), .CP(n4316), .CDN(
        n4344), .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N84), .E(n4268), .CP(n4319), .CDN(n4349), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(n4268), .CP(n4322), .CDN(
        n4359), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(n4269), .CP(n4278), .CDN(
        n4363), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(n4268), .CP(n4280), .CDN(
        n4334), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n4269), .CP(n4278), .CDN(
        n4363), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(n4268), .CP(n4313), .CDN(
        n4336), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n4268), .CP(n4308), .CDN(
        n4337), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(n4268), .CP(n4316), .CDN(
        n4356), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n4268), .CP(n4318), .CDN(
        n4362), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n4268), .CP(n4325), .CDN(
        n4359), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n4268), .CP(n4309), .CDN(
        n4344), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n4268), .CP(n4280), .CDN(
        n4353), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n4268), .CP(n4324), .CDN(
        n4354), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(n4268), .CP(n4280), .CDN(
        n4343), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(n4268), .CP(n4320), .CDN(
        n4344), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(n4268), .CP(n4317), .CDN(
        n4349), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n4269), .CP(n4319), .CDN(
        n4342), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n4269), .CP(ClockW), .CDN(
        n4341), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n4269), .CP(n4321), .CDN(
        n4340), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n4269), .CP(n4313), .CDN(
        n4350), .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(n4269), .CP(n4311), .CDN(
        n4356), .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(n4269), .CP(n4325), .CDN(
        n4336), .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(n4269), .CP(n4322), .CDN(
        n4337), .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(n4269), .CP(n4323), .CDN(
        n4352), .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n4269), .CP(n4280), .CDN(
        n4351), .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(n4269), .CP(n4279), .CDN(
        n4350), .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n4269), .CP(n4308), .CDN(
        n4352), .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(n4269), .CP(n4311), .CDN(
        n4351), .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(n4268), .CP(n4312), .CDN(
        n4350), .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N84), .E(n4270), .CP(n4309), .CDN(n4345), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(n4270), .CP(n4313), .CDN(
        n4339), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(n4270), .CP(n4314), .CDN(
        n4337), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(n4270), .CP(n4315), .CDN(
        n4343), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(n4270), .CP(n4319), .CDN(
        n4358), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(n4270), .CP(n4318), .CDN(
        n4362), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n4271), .CP(ClockW), .CDN(
        n4342), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n4271), .CP(n4322), .CDN(
        n4352), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n4270), .CP(n4318), .CDN(
        n4360), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n4271), .CP(n4317), .CDN(
        n4351), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n4270), .CP(n4316), .CDN(
        n4348), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n4271), .CP(n4320), .CDN(
        n4346), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n4270), .CP(n4323), .CDN(
        n4353), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(n4271), .CP(n4293), .CDN(
        n4363), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n4270), .CP(n4278), .CDN(
        n4347), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(n4271), .CP(n4321), .CDN(
        n4354), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n4271), .CP(n4290), .CDN(
        n4334), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n4271), .CP(n4306), .CDN(
        n4339), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n4271), .CP(n4308), .CDN(
        n4340), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n4271), .CP(n4309), .CDN(
        n4352), .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n4271), .CP(n4315), .CDN(
        n4357), .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(n4271), .CP(n4296), .CDN(
        n4358), .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(n4271), .CP(n4279), .CDN(
        n4352), .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(n4271), .CP(n4278), .CDN(
        n4352), .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n4271), .CP(n4280), .CDN(
        n4361), .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(n4271), .CP(n4324), .CDN(
        n4362), .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n4270), .CP(n4325), .CDN(
        n4335), .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(n4271), .CP(n4323), .CDN(
        n4338), .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(n4270), .CP(n4315), .CDN(
        n4350), .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N84), .E(n4276), .CP(n4314), .CDN(n4337), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(n4277), .CP(n4318), .CDN(
        n4336), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n4277), .CP(n4312), .CDN(
        n4336), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(n4276), .CP(n4308), .CDN(
        n4336), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n4277), .CP(n4322), .CDN(
        n4336), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n4276), .CP(n4322), .CDN(
        n4336), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(n4276), .CP(n4309), .CDN(
        n4336), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n4276), .CP(n4294), .CDN(
        n4336), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(n4276), .CP(n4313), .CDN(
        n4335), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(n4276), .CP(ClockW), .CDN(
        n4335), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(n4276), .CP(n4315), .CDN(
        n4335), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n4276), .CP(ClockW), .CDN(
        n4335), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n4276), .CP(n4321), .CDN(
        n4335), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(n4276), .CP(n4311), .CDN(
        n4335), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(n4276), .CP(n4318), .CDN(
        n4335), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(n4276), .CP(n4317), .CDN(
        n4335), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n4277), .CP(n4279), .CDN(
        n4335), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(n4277), .CP(n4315), .CDN(
        n4335), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(n4277), .CP(n4314), .CDN(
        n4335), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n4277), .CP(n4313), .CDN(
        n4334), .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(n4277), .CP(n4312), .CDN(
        n4334), .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(n4277), .CP(n4311), .CDN(
        n4334), .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(n4277), .CP(n4310), .CDN(
        n4334), .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(n4277), .CP(n4320), .CDN(
        n4334), .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n4277), .CP(n4316), .CDN(
        n4334), .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(n4277), .CP(ClockW), .CDN(
        n4334), .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n4277), .CP(n4280), .CDN(
        n4334), .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(n4276), .CP(n4278), .CDN(
        n4334), .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n4276), .CP(n4319), .CDN(
        n4334), .Q(\Storage[0][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n1797), .CP(ClockR), .CDN(n4334), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(n4249), .CP(n4285), .CDN(
        n4350), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(n4248), .CP(n4285), .CDN(
        n4359), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(n4249), .CP(n4285), .CDN(
        n4354), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(n4248), .CP(n4285), .CDN(
        n4351), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(DataI[28]), .E(n4251), .CP(n4288), .CDN(
        n4352), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(DataI[27]), .E(n4250), .CP(n4288), .CDN(
        n4363), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(DataI[26]), .E(n4251), .CP(n4289), .CDN(
        n4340), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(DataI[25]), .E(n4250), .CP(n4289), .CDN(
        n4340), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(DataI[28]), .E(n4257), .CP(n4299), .CDN(
        n4353), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(DataI[27]), .E(n4256), .CP(n4299), .CDN(
        n4334), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(DataI[26]), .E(n4257), .CP(n4300), .CDN(
        n4362), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(DataI[25]), .E(n4256), .CP(n4300), .CDN(
        n4361), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(DataI[28]), .E(n4258), .CP(n4288), .CDN(
        n4349), .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(DataI[27]), .E(n4258), .CP(n4289), .CDN(
        n4349), .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(DataI[26]), .E(n4258), .CP(n4305), .CDN(
        n4349), .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(DataI[25]), .E(n4258), .CP(n4306), .CDN(
        n4349), .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(n4265), .CP(n4321), .CDN(
        n4342), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(n4264), .CP(n4279), .CDN(
        n4342), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(n4265), .CP(n4311), .CDN(
        n4342), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(n4264), .CP(n4309), .CDN(
        n4342), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n4267), .CP(ClockW), .CDN(
        n4340), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n4266), .CP(n4289), .CDN(
        n4345), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(n4267), .CP(n4288), .CDN(
        n4362), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(n4266), .CP(n4286), .CDN(
        n4338), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n4273), .CP(n4311), .CDN(
        n4350), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n4272), .CP(n4310), .CDN(
        n4350), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n4273), .CP(n4313), .CDN(
        n4360), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(n4272), .CP(n4314), .CDN(
        n4362), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(n4275), .CP(n4310), .CDN(
        n4339), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(n4274), .CP(n4313), .CDN(
        n4339), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(n4275), .CP(ClockW), .CDN(
        n4339), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(n4274), .CP(n4304), .CDN(
        n4339), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(n4246), .CP(n4281), .CDN(
        n4353), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(n4247), .CP(n4281), .CDN(
        n4360), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(n4246), .CP(n4281), .CDN(
        n4361), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(n4247), .CP(n4281), .CDN(
        n4362), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(DataI[28]), .E(n4253), .CP(n4292), .CDN(
        n4361), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(DataI[27]), .E(n4252), .CP(n4292), .CDN(
        n4357), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(DataI[26]), .E(n4253), .CP(n4292), .CDN(
        n4335), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(DataI[25]), .E(n4252), .CP(n4292), .CDN(
        n4348), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(DataI[28]), .E(n4255), .CP(n4296), .CDN(
        n4361), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(DataI[27]), .E(n4254), .CP(n4296), .CDN(
        n4336), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(DataI[26]), .E(n4255), .CP(n4296), .CDN(
        n4334), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(DataI[25]), .E(n4254), .CP(n4296), .CDN(
        n4361), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(DataI[28]), .E(n4261), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(DataI[27]), .E(n4260), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(DataI[26]), .E(n4261), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(DataI[25]), .E(n4260), .CP(n4306), .CDN(
        n4346), .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n4263), .CP(n4310), .CDN(
        n4343), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(n4262), .CP(n4308), .CDN(
        n4343), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(n4263), .CP(n4300), .CDN(
        n4343), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(n4262), .CP(n4301), .CDN(
        n4343), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n4269), .CP(n4325), .CDN(
        n4344), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n4268), .CP(n4324), .CDN(
        n4345), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n4269), .CP(n4308), .CDN(
        n4346), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(n4268), .CP(n4303), .CDN(
        n4347), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(n4270), .CP(n4320), .CDN(
        n4352), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(n4270), .CP(n4318), .CDN(
        n4355), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n4270), .CP(n4316), .CDN(
        n4355), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(n4270), .CP(n4279), .CDN(
        n4345), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(n4277), .CP(n4324), .CDN(
        n4336), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(n4276), .CP(n4325), .CDN(
        n4336), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(n4277), .CP(n4323), .CDN(
        n4336), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(n4276), .CP(n4325), .CDN(
        n4336), .Q(\Storage[0][25] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n1860), .E(n4328), .CP(n4326), .CDN(n4358), 
        .Q(DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n1), .E(n4328), .CP(ClockR), .CDN(n4356), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n2), .E(n4329), .CP(n4326), .CDN(n4357), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n3), .E(n4328), .CP(ClockR), .CDN(n4351), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n2124), .E(n4329), .CP(n4326), .CDN(n4357), 
        .Q(DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n4), .E(n4328), .CP(ClockR), .CDN(n4360), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n5), .E(n4329), .CP(n4326), .CDN(n4344), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n2322), .E(n4328), .CP(n4326), .CDN(n4357), 
        .Q(DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n2388), .E(n4329), .CP(ClockR), .CDN(n4350), 
        .Q(DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n2454), .E(n4328), .CP(n4326), .CDN(n4335), 
        .Q(DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n2519), .E(n4328), .CP(ClockR), .CDN(n4351), 
        .Q(DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n2585), .E(n4328), .CP(n4326), .CDN(n4352), 
        .Q(DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n2651), .E(n4328), .CP(ClockR), .CDN(n4353), 
        .Q(DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n2717), .E(n4328), .CP(n4326), .CDN(n4360), 
        .Q(DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n6), .E(n4328), .CP(ClockR), .CDN(n4350), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n2846), .E(n4328), .CP(n4326), .CDN(n4352), 
        .Q(DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n2909), .E(n4328), .CP(ClockR), .CDN(n4351), 
        .Q(DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n2972), .E(n4328), .CP(n4326), .CDN(n4355), 
        .Q(DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n3034), .E(n4328), .CP(n4326), .CDN(n4361), 
        .Q(DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n3096), .E(n4328), .CP(n4326), .CDN(n4336), 
        .Q(DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n3159), .E(n4329), .CP(n4326), .CDN(n4337), 
        .Q(DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n3222), .E(n4329), .CP(n4326), .CDN(n4341), 
        .Q(DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n3283), .E(n4329), .CP(n4326), .CDN(n4356), 
        .Q(DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n3341), .E(n4329), .CP(n4326), .CDN(n4354), 
        .Q(DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n3398), .E(n4329), .CP(n4326), .CDN(n4346), 
        .Q(DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n3458), .E(n4329), .CP(n4326), .CDN(n4359), 
        .Q(DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n3517), .E(n4329), .CP(n4326), .CDN(n4361), 
        .Q(DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n7), .E(n4329), .CP(ClockR), .CDN(n4339), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n3635), .E(n4329), .CP(ClockR), .CDN(n4360), 
        .Q(DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n3691), .E(n4329), .CP(ClockR), .CDN(n4342), 
        .Q(DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n3750), .E(n9), .CP(ClockR), .CDN(n4358), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n8), .E(n9), .CP(ClockR), .CDN(n4334), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(n3873), .E(n9), .CP(ClockR), .CDN(n4359), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(n1742), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(n1687), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(n1632), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(n1577), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(n1522), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(n1468), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(n1414), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(n1360), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(n1306), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(n1252), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(n1198), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(n1144), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(n1090), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(n1036), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(n982), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(n928), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(n874), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(n820), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(n766), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(n712), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(n658), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(n604), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(n550), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(n496), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(n442), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(n388), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(n334), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(n280), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(n226), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(n172), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(n118), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(n27), .OE(ChipEna), .Z(DataO[31]) );
  CKBD0 U3 ( .CLK(N50), .C(n1861) );
  BUFFD0 U4 ( .I(n1926), .Z(n1) );
  BUFFD0 U5 ( .I(n1992), .Z(n2) );
  BUFFD0 U6 ( .I(n2058), .Z(n3) );
  CKBD0 U7 ( .CLK(N54), .C(n2125) );
  BUFFD0 U8 ( .I(n2190), .Z(n4) );
  BUFFD0 U9 ( .I(n2256), .Z(n5) );
  CKBD0 U10 ( .CLK(N57), .C(n2323) );
  BUFFD0 U11 ( .I(n2783), .Z(n6) );
  BUFFD0 U12 ( .I(n3576), .Z(n7) );
  CKBD0 U18 ( .CLK(n4027), .C(n4017) );
  CKBD0 U19 ( .CLK(n4026), .C(n4016) );
  BUFFD0 U20 ( .I(n3809), .Z(n8) );
  XOR3D4 U23 ( .A1(n4038), .A2(n4037), .A3(n77), .Z(N82) );
  XOR3D0 U24 ( .A1(n4031), .A2(n78), .A3(n79), .Z(n77) );
  BUFFD0 U25 ( .I(n4044), .Z(n9) );
  XNR3D1 U26 ( .A1(n3933), .A2(n84), .A3(n10), .ZN(n83) );
  XNR3D1 U31 ( .A1(n3925), .A2(n3943), .A3(n86), .ZN(n10) );
  CKBXD0 U32 ( .I(N44), .Z(n4332) );
  OR2D1 U33 ( .A1(n89), .A2(n93), .Z(n11) );
  OR2D1 U34 ( .A1(n91), .A2(n92), .Z(n12) );
  OR2D1 U35 ( .A1(n91), .A2(n93), .Z(n13) );
  OR2D1 U36 ( .A1(n89), .A2(n92), .Z(n14) );
  OR2D1 U37 ( .A1(n89), .A2(n90), .Z(n15) );
  OR2D1 U38 ( .A1(n94), .A2(n98), .Z(n16) );
  INVD0 U39 ( .I(N47), .ZN(n4231) );
  OR2D1 U40 ( .A1(n89), .A2(n94), .Z(n17) );
  OR2D1 U41 ( .A1(n91), .A2(n94), .Z(n18) );
  OR2D1 U42 ( .A1(n92), .A2(n98), .Z(n19) );
  OR2D1 U43 ( .A1(n94), .A2(n97), .Z(n20) );
  OR2D1 U44 ( .A1(n92), .A2(n97), .Z(n21) );
  OR2D1 U45 ( .A1(n93), .A2(n97), .Z(n22) );
  OR2D1 U46 ( .A1(n90), .A2(n97), .Z(n23) );
  OR2D1 U47 ( .A1(n90), .A2(n91), .Z(n24) );
  OR2D1 U48 ( .A1(n93), .A2(n98), .Z(n25) );
  OR2D1 U49 ( .A1(n90), .A2(n98), .Z(n26) );
  BUFFD0 U50 ( .I(n28), .Z(n27) );
  BUFFD0 U51 ( .I(n29), .Z(n28) );
  BUFFD0 U52 ( .I(n30), .Z(n29) );
  BUFFD0 U53 ( .I(n31), .Z(n30) );
  BUFFD0 U54 ( .I(n32), .Z(n31) );
  BUFFD0 U55 ( .I(n33), .Z(n32) );
  BUFFD0 U56 ( .I(n34), .Z(n33) );
  BUFFD0 U57 ( .I(n35), .Z(n34) );
  BUFFD0 U58 ( .I(n36), .Z(n35) );
  BUFFD0 U59 ( .I(n37), .Z(n36) );
  BUFFD0 U60 ( .I(n38), .Z(n37) );
  BUFFD0 U61 ( .I(n39), .Z(n38) );
  BUFFD0 U62 ( .I(n40), .Z(n39) );
  BUFFD0 U63 ( .I(n41), .Z(n40) );
  BUFFD0 U64 ( .I(n42), .Z(n41) );
  BUFFD0 U65 ( .I(n43), .Z(n42) );
  BUFFD0 U66 ( .I(n44), .Z(n43) );
  BUFFD0 U67 ( .I(n45), .Z(n44) );
  BUFFD0 U68 ( .I(n46), .Z(n45) );
  BUFFD0 U69 ( .I(n47), .Z(n46) );
  BUFFD0 U70 ( .I(n48), .Z(n47) );
  BUFFD0 U71 ( .I(n49), .Z(n48) );
  BUFFD0 U72 ( .I(n50), .Z(n49) );
  BUFFD0 U73 ( .I(n51), .Z(n50) );
  BUFFD0 U74 ( .I(n52), .Z(n51) );
  BUFFD0 U75 ( .I(n53), .Z(n52) );
  BUFFD0 U76 ( .I(n54), .Z(n53) );
  BUFFD0 U77 ( .I(n55), .Z(n54) );
  BUFFD0 U78 ( .I(n56), .Z(n55) );
  BUFFD0 U79 ( .I(n57), .Z(n56) );
  BUFFD0 U80 ( .I(n58), .Z(n57) );
  BUFFD0 U81 ( .I(n59), .Z(n58) );
  BUFFD0 U82 ( .I(n60), .Z(n59) );
  BUFFD0 U83 ( .I(n61), .Z(n60) );
  BUFFD0 U84 ( .I(n62), .Z(n61) );
  BUFFD0 U85 ( .I(n63), .Z(n62) );
  BUFFD0 U86 ( .I(n64), .Z(n63) );
  BUFFD0 U87 ( .I(n85), .Z(n64) );
  BUFFD0 U88 ( .I(n102), .Z(n85) );
  BUFFD0 U89 ( .I(n104), .Z(n102) );
  BUFFD0 U90 ( .I(n105), .Z(n104) );
  BUFFD0 U91 ( .I(n106), .Z(n105) );
  BUFFD0 U92 ( .I(n107), .Z(n106) );
  BUFFD0 U93 ( .I(n108), .Z(n107) );
  BUFFD0 U94 ( .I(n109), .Z(n108) );
  BUFFD0 U95 ( .I(n110), .Z(n109) );
  BUFFD0 U96 ( .I(n111), .Z(n110) );
  BUFFD0 U97 ( .I(n112), .Z(n111) );
  BUFFD0 U98 ( .I(n113), .Z(n112) );
  BUFFD0 U99 ( .I(n114), .Z(n113) );
  BUFFD0 U100 ( .I(n115), .Z(n114) );
  BUFFD0 U101 ( .I(n116), .Z(n115) );
  BUFFD0 U102 ( .I(n117), .Z(n116) );
  BUFFD0 U103 ( .I(DataOr[31]), .Z(n117) );
  BUFFD0 U104 ( .I(n119), .Z(n118) );
  BUFFD0 U105 ( .I(n120), .Z(n119) );
  BUFFD0 U106 ( .I(n121), .Z(n120) );
  BUFFD0 U107 ( .I(n122), .Z(n121) );
  BUFFD0 U108 ( .I(n123), .Z(n122) );
  BUFFD0 U109 ( .I(n124), .Z(n123) );
  BUFFD0 U110 ( .I(n125), .Z(n124) );
  BUFFD0 U111 ( .I(n126), .Z(n125) );
  BUFFD0 U112 ( .I(n127), .Z(n126) );
  BUFFD0 U113 ( .I(n128), .Z(n127) );
  BUFFD0 U114 ( .I(n129), .Z(n128) );
  BUFFD0 U115 ( .I(n130), .Z(n129) );
  BUFFD0 U116 ( .I(n131), .Z(n130) );
  BUFFD0 U117 ( .I(n132), .Z(n131) );
  BUFFD0 U118 ( .I(n133), .Z(n132) );
  BUFFD0 U119 ( .I(n134), .Z(n133) );
  BUFFD0 U120 ( .I(n135), .Z(n134) );
  BUFFD0 U121 ( .I(n136), .Z(n135) );
  BUFFD0 U122 ( .I(n137), .Z(n136) );
  BUFFD0 U123 ( .I(n138), .Z(n137) );
  BUFFD0 U124 ( .I(n139), .Z(n138) );
  BUFFD0 U125 ( .I(n140), .Z(n139) );
  BUFFD0 U126 ( .I(n141), .Z(n140) );
  BUFFD0 U127 ( .I(n142), .Z(n141) );
  BUFFD0 U128 ( .I(n143), .Z(n142) );
  BUFFD0 U129 ( .I(n144), .Z(n143) );
  BUFFD0 U130 ( .I(n145), .Z(n144) );
  BUFFD0 U131 ( .I(n146), .Z(n145) );
  BUFFD0 U132 ( .I(n147), .Z(n146) );
  BUFFD0 U133 ( .I(n148), .Z(n147) );
  BUFFD0 U134 ( .I(n149), .Z(n148) );
  BUFFD0 U135 ( .I(n150), .Z(n149) );
  BUFFD0 U136 ( .I(n151), .Z(n150) );
  BUFFD0 U137 ( .I(n152), .Z(n151) );
  BUFFD0 U138 ( .I(n153), .Z(n152) );
  BUFFD0 U139 ( .I(n154), .Z(n153) );
  BUFFD0 U140 ( .I(n155), .Z(n154) );
  BUFFD0 U141 ( .I(n156), .Z(n155) );
  BUFFD0 U142 ( .I(n157), .Z(n156) );
  BUFFD0 U143 ( .I(n158), .Z(n157) );
  BUFFD0 U144 ( .I(n159), .Z(n158) );
  BUFFD0 U145 ( .I(n160), .Z(n159) );
  BUFFD0 U146 ( .I(n161), .Z(n160) );
  BUFFD0 U147 ( .I(n162), .Z(n161) );
  BUFFD0 U148 ( .I(n163), .Z(n162) );
  BUFFD0 U149 ( .I(n164), .Z(n163) );
  BUFFD0 U150 ( .I(n165), .Z(n164) );
  BUFFD0 U151 ( .I(n166), .Z(n165) );
  BUFFD0 U152 ( .I(n167), .Z(n166) );
  BUFFD0 U153 ( .I(n168), .Z(n167) );
  BUFFD0 U154 ( .I(n169), .Z(n168) );
  BUFFD0 U155 ( .I(n170), .Z(n169) );
  BUFFD0 U156 ( .I(n171), .Z(n170) );
  BUFFD0 U157 ( .I(DataOr[30]), .Z(n171) );
  BUFFD0 U158 ( .I(n173), .Z(n172) );
  BUFFD0 U159 ( .I(n174), .Z(n173) );
  BUFFD0 U160 ( .I(n175), .Z(n174) );
  BUFFD0 U161 ( .I(n176), .Z(n175) );
  BUFFD0 U162 ( .I(n177), .Z(n176) );
  BUFFD0 U163 ( .I(n178), .Z(n177) );
  BUFFD0 U164 ( .I(n179), .Z(n178) );
  BUFFD0 U165 ( .I(n180), .Z(n179) );
  BUFFD0 U166 ( .I(n181), .Z(n180) );
  BUFFD0 U167 ( .I(n182), .Z(n181) );
  BUFFD0 U168 ( .I(n183), .Z(n182) );
  BUFFD0 U169 ( .I(n184), .Z(n183) );
  BUFFD0 U170 ( .I(n185), .Z(n184) );
  BUFFD0 U171 ( .I(n186), .Z(n185) );
  BUFFD0 U172 ( .I(n187), .Z(n186) );
  BUFFD0 U173 ( .I(n188), .Z(n187) );
  BUFFD0 U174 ( .I(n189), .Z(n188) );
  BUFFD0 U175 ( .I(n190), .Z(n189) );
  BUFFD0 U176 ( .I(n191), .Z(n190) );
  BUFFD0 U177 ( .I(n192), .Z(n191) );
  BUFFD0 U178 ( .I(n193), .Z(n192) );
  BUFFD0 U179 ( .I(n194), .Z(n193) );
  BUFFD0 U180 ( .I(n195), .Z(n194) );
  BUFFD0 U181 ( .I(n196), .Z(n195) );
  BUFFD0 U182 ( .I(n197), .Z(n196) );
  BUFFD0 U183 ( .I(n198), .Z(n197) );
  BUFFD0 U184 ( .I(n199), .Z(n198) );
  BUFFD0 U185 ( .I(n200), .Z(n199) );
  BUFFD0 U186 ( .I(n201), .Z(n200) );
  BUFFD0 U187 ( .I(n202), .Z(n201) );
  BUFFD0 U188 ( .I(n203), .Z(n202) );
  BUFFD0 U189 ( .I(n204), .Z(n203) );
  BUFFD0 U190 ( .I(n205), .Z(n204) );
  BUFFD0 U191 ( .I(n206), .Z(n205) );
  BUFFD0 U192 ( .I(n207), .Z(n206) );
  BUFFD0 U193 ( .I(n208), .Z(n207) );
  BUFFD0 U194 ( .I(n209), .Z(n208) );
  BUFFD0 U195 ( .I(n210), .Z(n209) );
  BUFFD0 U196 ( .I(n211), .Z(n210) );
  BUFFD0 U197 ( .I(n212), .Z(n211) );
  BUFFD0 U198 ( .I(n213), .Z(n212) );
  BUFFD0 U199 ( .I(n214), .Z(n213) );
  BUFFD0 U200 ( .I(n215), .Z(n214) );
  BUFFD0 U201 ( .I(n216), .Z(n215) );
  BUFFD0 U202 ( .I(n217), .Z(n216) );
  BUFFD0 U203 ( .I(n218), .Z(n217) );
  BUFFD0 U204 ( .I(n219), .Z(n218) );
  BUFFD0 U205 ( .I(n220), .Z(n219) );
  BUFFD0 U206 ( .I(n221), .Z(n220) );
  BUFFD0 U207 ( .I(n222), .Z(n221) );
  BUFFD0 U208 ( .I(n223), .Z(n222) );
  BUFFD0 U209 ( .I(n224), .Z(n223) );
  BUFFD0 U210 ( .I(n225), .Z(n224) );
  BUFFD0 U211 ( .I(DataOr[29]), .Z(n225) );
  BUFFD0 U212 ( .I(n227), .Z(n226) );
  BUFFD0 U213 ( .I(n228), .Z(n227) );
  BUFFD0 U214 ( .I(n229), .Z(n228) );
  BUFFD0 U215 ( .I(n230), .Z(n229) );
  BUFFD0 U216 ( .I(n231), .Z(n230) );
  BUFFD0 U217 ( .I(n232), .Z(n231) );
  BUFFD0 U218 ( .I(n233), .Z(n232) );
  BUFFD0 U219 ( .I(n234), .Z(n233) );
  BUFFD0 U220 ( .I(n235), .Z(n234) );
  BUFFD0 U221 ( .I(n236), .Z(n235) );
  BUFFD0 U222 ( .I(n237), .Z(n236) );
  BUFFD0 U223 ( .I(n238), .Z(n237) );
  BUFFD0 U224 ( .I(n239), .Z(n238) );
  BUFFD0 U225 ( .I(n240), .Z(n239) );
  BUFFD0 U226 ( .I(n241), .Z(n240) );
  BUFFD0 U227 ( .I(n242), .Z(n241) );
  BUFFD0 U228 ( .I(n243), .Z(n242) );
  BUFFD0 U229 ( .I(n244), .Z(n243) );
  BUFFD0 U230 ( .I(n245), .Z(n244) );
  BUFFD0 U231 ( .I(n246), .Z(n245) );
  BUFFD0 U232 ( .I(n247), .Z(n246) );
  BUFFD0 U233 ( .I(n248), .Z(n247) );
  BUFFD0 U234 ( .I(n249), .Z(n248) );
  BUFFD0 U235 ( .I(n250), .Z(n249) );
  BUFFD0 U236 ( .I(n251), .Z(n250) );
  BUFFD0 U237 ( .I(n252), .Z(n251) );
  BUFFD0 U238 ( .I(n253), .Z(n252) );
  BUFFD0 U239 ( .I(n254), .Z(n253) );
  BUFFD0 U240 ( .I(n255), .Z(n254) );
  BUFFD0 U241 ( .I(n256), .Z(n255) );
  BUFFD0 U242 ( .I(n257), .Z(n256) );
  BUFFD0 U243 ( .I(n258), .Z(n257) );
  BUFFD0 U244 ( .I(n259), .Z(n258) );
  BUFFD0 U245 ( .I(n260), .Z(n259) );
  BUFFD0 U246 ( .I(n261), .Z(n260) );
  BUFFD0 U247 ( .I(n262), .Z(n261) );
  BUFFD0 U248 ( .I(n263), .Z(n262) );
  BUFFD0 U249 ( .I(n264), .Z(n263) );
  BUFFD0 U250 ( .I(n265), .Z(n264) );
  BUFFD0 U251 ( .I(n266), .Z(n265) );
  BUFFD0 U252 ( .I(n267), .Z(n266) );
  BUFFD0 U253 ( .I(n268), .Z(n267) );
  BUFFD0 U254 ( .I(n269), .Z(n268) );
  BUFFD0 U255 ( .I(n270), .Z(n269) );
  BUFFD0 U256 ( .I(n271), .Z(n270) );
  BUFFD0 U257 ( .I(n272), .Z(n271) );
  BUFFD0 U258 ( .I(n273), .Z(n272) );
  BUFFD0 U259 ( .I(n274), .Z(n273) );
  BUFFD0 U260 ( .I(n275), .Z(n274) );
  BUFFD0 U261 ( .I(n276), .Z(n275) );
  BUFFD0 U262 ( .I(n277), .Z(n276) );
  BUFFD0 U263 ( .I(n278), .Z(n277) );
  BUFFD0 U264 ( .I(n279), .Z(n278) );
  BUFFD0 U265 ( .I(DataOr[28]), .Z(n279) );
  BUFFD0 U266 ( .I(n281), .Z(n280) );
  BUFFD0 U267 ( .I(n282), .Z(n281) );
  BUFFD0 U268 ( .I(n283), .Z(n282) );
  BUFFD0 U269 ( .I(n284), .Z(n283) );
  BUFFD0 U270 ( .I(n285), .Z(n284) );
  BUFFD0 U271 ( .I(n286), .Z(n285) );
  BUFFD0 U272 ( .I(n287), .Z(n286) );
  BUFFD0 U273 ( .I(n288), .Z(n287) );
  BUFFD0 U274 ( .I(n289), .Z(n288) );
  BUFFD0 U275 ( .I(n290), .Z(n289) );
  BUFFD0 U276 ( .I(n291), .Z(n290) );
  BUFFD0 U277 ( .I(n292), .Z(n291) );
  BUFFD0 U278 ( .I(n293), .Z(n292) );
  BUFFD0 U279 ( .I(n294), .Z(n293) );
  BUFFD0 U280 ( .I(n295), .Z(n294) );
  BUFFD0 U281 ( .I(n296), .Z(n295) );
  BUFFD0 U282 ( .I(n297), .Z(n296) );
  BUFFD0 U283 ( .I(n298), .Z(n297) );
  BUFFD0 U284 ( .I(n299), .Z(n298) );
  BUFFD0 U285 ( .I(n300), .Z(n299) );
  BUFFD0 U286 ( .I(n301), .Z(n300) );
  BUFFD0 U287 ( .I(n302), .Z(n301) );
  BUFFD0 U288 ( .I(n303), .Z(n302) );
  BUFFD0 U289 ( .I(n304), .Z(n303) );
  BUFFD0 U290 ( .I(n305), .Z(n304) );
  BUFFD0 U291 ( .I(n306), .Z(n305) );
  BUFFD0 U292 ( .I(n307), .Z(n306) );
  BUFFD0 U293 ( .I(n308), .Z(n307) );
  BUFFD0 U294 ( .I(n309), .Z(n308) );
  BUFFD0 U295 ( .I(n310), .Z(n309) );
  BUFFD0 U296 ( .I(n311), .Z(n310) );
  BUFFD0 U297 ( .I(n312), .Z(n311) );
  BUFFD0 U298 ( .I(n313), .Z(n312) );
  BUFFD0 U299 ( .I(n314), .Z(n313) );
  BUFFD0 U300 ( .I(n315), .Z(n314) );
  BUFFD0 U301 ( .I(n316), .Z(n315) );
  BUFFD0 U302 ( .I(n317), .Z(n316) );
  BUFFD0 U303 ( .I(n318), .Z(n317) );
  BUFFD0 U304 ( .I(n319), .Z(n318) );
  BUFFD0 U305 ( .I(n320), .Z(n319) );
  BUFFD0 U306 ( .I(n321), .Z(n320) );
  BUFFD0 U307 ( .I(n322), .Z(n321) );
  BUFFD0 U308 ( .I(n323), .Z(n322) );
  BUFFD0 U309 ( .I(n324), .Z(n323) );
  BUFFD0 U310 ( .I(n325), .Z(n324) );
  BUFFD0 U311 ( .I(n326), .Z(n325) );
  BUFFD0 U312 ( .I(n327), .Z(n326) );
  BUFFD0 U313 ( .I(n328), .Z(n327) );
  BUFFD0 U314 ( .I(n329), .Z(n328) );
  BUFFD0 U315 ( .I(n330), .Z(n329) );
  BUFFD0 U316 ( .I(n331), .Z(n330) );
  BUFFD0 U317 ( .I(n332), .Z(n331) );
  BUFFD0 U318 ( .I(n333), .Z(n332) );
  BUFFD0 U319 ( .I(DataOr[27]), .Z(n333) );
  BUFFD0 U320 ( .I(n335), .Z(n334) );
  BUFFD0 U321 ( .I(n336), .Z(n335) );
  BUFFD0 U322 ( .I(n337), .Z(n336) );
  BUFFD0 U323 ( .I(n338), .Z(n337) );
  BUFFD0 U324 ( .I(n339), .Z(n338) );
  BUFFD0 U325 ( .I(n340), .Z(n339) );
  BUFFD0 U326 ( .I(n341), .Z(n340) );
  BUFFD0 U327 ( .I(n342), .Z(n341) );
  BUFFD0 U328 ( .I(n343), .Z(n342) );
  BUFFD0 U329 ( .I(n344), .Z(n343) );
  BUFFD0 U330 ( .I(n345), .Z(n344) );
  BUFFD0 U331 ( .I(n346), .Z(n345) );
  BUFFD0 U332 ( .I(n347), .Z(n346) );
  BUFFD0 U333 ( .I(n348), .Z(n347) );
  BUFFD0 U334 ( .I(n349), .Z(n348) );
  BUFFD0 U335 ( .I(n350), .Z(n349) );
  BUFFD0 U336 ( .I(n351), .Z(n350) );
  BUFFD0 U337 ( .I(n352), .Z(n351) );
  BUFFD0 U338 ( .I(n353), .Z(n352) );
  BUFFD0 U339 ( .I(n354), .Z(n353) );
  BUFFD0 U340 ( .I(n355), .Z(n354) );
  BUFFD0 U341 ( .I(n356), .Z(n355) );
  BUFFD0 U342 ( .I(n357), .Z(n356) );
  BUFFD0 U343 ( .I(n358), .Z(n357) );
  BUFFD0 U344 ( .I(n359), .Z(n358) );
  BUFFD0 U345 ( .I(n360), .Z(n359) );
  BUFFD0 U346 ( .I(n361), .Z(n360) );
  BUFFD0 U347 ( .I(n362), .Z(n361) );
  BUFFD0 U348 ( .I(n363), .Z(n362) );
  BUFFD0 U349 ( .I(n364), .Z(n363) );
  BUFFD0 U350 ( .I(n365), .Z(n364) );
  BUFFD0 U351 ( .I(n366), .Z(n365) );
  BUFFD0 U352 ( .I(n367), .Z(n366) );
  BUFFD0 U353 ( .I(n368), .Z(n367) );
  BUFFD0 U354 ( .I(n369), .Z(n368) );
  BUFFD0 U355 ( .I(n370), .Z(n369) );
  BUFFD0 U356 ( .I(n371), .Z(n370) );
  BUFFD0 U357 ( .I(n372), .Z(n371) );
  BUFFD0 U358 ( .I(n373), .Z(n372) );
  BUFFD0 U359 ( .I(n374), .Z(n373) );
  BUFFD0 U360 ( .I(n375), .Z(n374) );
  BUFFD0 U361 ( .I(n376), .Z(n375) );
  BUFFD0 U362 ( .I(n377), .Z(n376) );
  BUFFD0 U363 ( .I(n378), .Z(n377) );
  BUFFD0 U364 ( .I(n379), .Z(n378) );
  BUFFD0 U365 ( .I(n380), .Z(n379) );
  BUFFD0 U366 ( .I(n381), .Z(n380) );
  BUFFD0 U367 ( .I(n382), .Z(n381) );
  BUFFD0 U368 ( .I(n383), .Z(n382) );
  BUFFD0 U369 ( .I(n384), .Z(n383) );
  BUFFD0 U370 ( .I(n385), .Z(n384) );
  BUFFD0 U371 ( .I(n386), .Z(n385) );
  BUFFD0 U372 ( .I(n387), .Z(n386) );
  BUFFD0 U373 ( .I(DataOr[26]), .Z(n387) );
  BUFFD0 U374 ( .I(n389), .Z(n388) );
  BUFFD0 U375 ( .I(n390), .Z(n389) );
  BUFFD0 U376 ( .I(n391), .Z(n390) );
  BUFFD0 U377 ( .I(n392), .Z(n391) );
  BUFFD0 U378 ( .I(n393), .Z(n392) );
  BUFFD0 U379 ( .I(n394), .Z(n393) );
  BUFFD0 U380 ( .I(n395), .Z(n394) );
  BUFFD0 U381 ( .I(n396), .Z(n395) );
  BUFFD0 U382 ( .I(n397), .Z(n396) );
  BUFFD0 U383 ( .I(n398), .Z(n397) );
  BUFFD0 U384 ( .I(n399), .Z(n398) );
  BUFFD0 U385 ( .I(n400), .Z(n399) );
  BUFFD0 U386 ( .I(n401), .Z(n400) );
  BUFFD0 U387 ( .I(n402), .Z(n401) );
  BUFFD0 U388 ( .I(n403), .Z(n402) );
  BUFFD0 U389 ( .I(n404), .Z(n403) );
  BUFFD0 U390 ( .I(n405), .Z(n404) );
  BUFFD0 U391 ( .I(n406), .Z(n405) );
  BUFFD0 U392 ( .I(n407), .Z(n406) );
  BUFFD0 U393 ( .I(n408), .Z(n407) );
  BUFFD0 U394 ( .I(n409), .Z(n408) );
  BUFFD0 U395 ( .I(n410), .Z(n409) );
  BUFFD0 U396 ( .I(n411), .Z(n410) );
  BUFFD0 U397 ( .I(n412), .Z(n411) );
  BUFFD0 U398 ( .I(n413), .Z(n412) );
  BUFFD0 U399 ( .I(n414), .Z(n413) );
  BUFFD0 U400 ( .I(n415), .Z(n414) );
  BUFFD0 U401 ( .I(n416), .Z(n415) );
  BUFFD0 U402 ( .I(n417), .Z(n416) );
  BUFFD0 U403 ( .I(n418), .Z(n417) );
  BUFFD0 U404 ( .I(n419), .Z(n418) );
  BUFFD0 U405 ( .I(n420), .Z(n419) );
  BUFFD0 U406 ( .I(n421), .Z(n420) );
  BUFFD0 U407 ( .I(n422), .Z(n421) );
  BUFFD0 U408 ( .I(n423), .Z(n422) );
  BUFFD0 U409 ( .I(n424), .Z(n423) );
  BUFFD0 U410 ( .I(n425), .Z(n424) );
  BUFFD0 U411 ( .I(n426), .Z(n425) );
  BUFFD0 U412 ( .I(n427), .Z(n426) );
  BUFFD0 U413 ( .I(n428), .Z(n427) );
  BUFFD0 U414 ( .I(n429), .Z(n428) );
  BUFFD0 U415 ( .I(n430), .Z(n429) );
  BUFFD0 U416 ( .I(n431), .Z(n430) );
  BUFFD0 U417 ( .I(n432), .Z(n431) );
  BUFFD0 U418 ( .I(n433), .Z(n432) );
  BUFFD0 U419 ( .I(n434), .Z(n433) );
  BUFFD0 U420 ( .I(n435), .Z(n434) );
  BUFFD0 U421 ( .I(n436), .Z(n435) );
  BUFFD0 U422 ( .I(n437), .Z(n436) );
  BUFFD0 U423 ( .I(n438), .Z(n437) );
  BUFFD0 U424 ( .I(n439), .Z(n438) );
  BUFFD0 U425 ( .I(n440), .Z(n439) );
  BUFFD0 U426 ( .I(n441), .Z(n440) );
  BUFFD0 U427 ( .I(DataOr[25]), .Z(n441) );
  BUFFD0 U428 ( .I(n443), .Z(n442) );
  BUFFD0 U429 ( .I(n444), .Z(n443) );
  BUFFD0 U430 ( .I(n445), .Z(n444) );
  BUFFD0 U431 ( .I(n446), .Z(n445) );
  BUFFD0 U432 ( .I(n447), .Z(n446) );
  BUFFD0 U433 ( .I(n448), .Z(n447) );
  BUFFD0 U434 ( .I(n449), .Z(n448) );
  BUFFD0 U435 ( .I(n450), .Z(n449) );
  BUFFD0 U436 ( .I(n451), .Z(n450) );
  BUFFD0 U437 ( .I(n452), .Z(n451) );
  BUFFD0 U438 ( .I(n453), .Z(n452) );
  BUFFD0 U439 ( .I(n454), .Z(n453) );
  BUFFD0 U440 ( .I(n455), .Z(n454) );
  BUFFD0 U441 ( .I(n456), .Z(n455) );
  BUFFD0 U442 ( .I(n457), .Z(n456) );
  BUFFD0 U443 ( .I(n458), .Z(n457) );
  BUFFD0 U444 ( .I(n459), .Z(n458) );
  BUFFD0 U445 ( .I(n460), .Z(n459) );
  BUFFD0 U446 ( .I(n461), .Z(n460) );
  BUFFD0 U447 ( .I(n462), .Z(n461) );
  BUFFD0 U448 ( .I(n463), .Z(n462) );
  BUFFD0 U449 ( .I(n464), .Z(n463) );
  BUFFD0 U450 ( .I(n465), .Z(n464) );
  BUFFD0 U451 ( .I(n466), .Z(n465) );
  BUFFD0 U452 ( .I(n467), .Z(n466) );
  BUFFD0 U453 ( .I(n468), .Z(n467) );
  BUFFD0 U454 ( .I(n469), .Z(n468) );
  BUFFD0 U455 ( .I(n470), .Z(n469) );
  BUFFD0 U456 ( .I(n471), .Z(n470) );
  BUFFD0 U457 ( .I(n472), .Z(n471) );
  BUFFD0 U458 ( .I(n473), .Z(n472) );
  BUFFD0 U459 ( .I(n474), .Z(n473) );
  BUFFD0 U460 ( .I(n475), .Z(n474) );
  BUFFD0 U461 ( .I(n476), .Z(n475) );
  BUFFD0 U462 ( .I(n477), .Z(n476) );
  BUFFD0 U463 ( .I(n478), .Z(n477) );
  BUFFD0 U464 ( .I(n479), .Z(n478) );
  BUFFD0 U465 ( .I(n480), .Z(n479) );
  BUFFD0 U466 ( .I(n481), .Z(n480) );
  BUFFD0 U467 ( .I(n482), .Z(n481) );
  BUFFD0 U468 ( .I(n483), .Z(n482) );
  BUFFD0 U469 ( .I(n484), .Z(n483) );
  BUFFD0 U470 ( .I(n485), .Z(n484) );
  BUFFD0 U471 ( .I(n486), .Z(n485) );
  BUFFD0 U472 ( .I(n487), .Z(n486) );
  BUFFD0 U473 ( .I(n488), .Z(n487) );
  BUFFD0 U474 ( .I(n489), .Z(n488) );
  BUFFD0 U475 ( .I(n490), .Z(n489) );
  BUFFD0 U476 ( .I(n491), .Z(n490) );
  BUFFD0 U477 ( .I(n492), .Z(n491) );
  BUFFD0 U478 ( .I(n493), .Z(n492) );
  BUFFD0 U479 ( .I(n494), .Z(n493) );
  BUFFD0 U480 ( .I(n495), .Z(n494) );
  BUFFD0 U481 ( .I(DataOr[24]), .Z(n495) );
  BUFFD0 U482 ( .I(n497), .Z(n496) );
  BUFFD0 U483 ( .I(n498), .Z(n497) );
  BUFFD0 U484 ( .I(n499), .Z(n498) );
  BUFFD0 U485 ( .I(n500), .Z(n499) );
  BUFFD0 U486 ( .I(n501), .Z(n500) );
  BUFFD0 U487 ( .I(n502), .Z(n501) );
  BUFFD0 U488 ( .I(n503), .Z(n502) );
  BUFFD0 U489 ( .I(n504), .Z(n503) );
  BUFFD0 U490 ( .I(n505), .Z(n504) );
  BUFFD0 U491 ( .I(n506), .Z(n505) );
  BUFFD0 U492 ( .I(n507), .Z(n506) );
  BUFFD0 U493 ( .I(n508), .Z(n507) );
  BUFFD0 U494 ( .I(n509), .Z(n508) );
  BUFFD0 U495 ( .I(n510), .Z(n509) );
  BUFFD0 U496 ( .I(n511), .Z(n510) );
  BUFFD0 U497 ( .I(n512), .Z(n511) );
  BUFFD0 U498 ( .I(n513), .Z(n512) );
  BUFFD0 U499 ( .I(n514), .Z(n513) );
  BUFFD0 U500 ( .I(n515), .Z(n514) );
  BUFFD0 U501 ( .I(n516), .Z(n515) );
  BUFFD0 U502 ( .I(n517), .Z(n516) );
  BUFFD0 U503 ( .I(n518), .Z(n517) );
  BUFFD0 U504 ( .I(n519), .Z(n518) );
  BUFFD0 U505 ( .I(n520), .Z(n519) );
  BUFFD0 U506 ( .I(n521), .Z(n520) );
  BUFFD0 U507 ( .I(n522), .Z(n521) );
  BUFFD0 U508 ( .I(n523), .Z(n522) );
  BUFFD0 U509 ( .I(n524), .Z(n523) );
  BUFFD0 U510 ( .I(n525), .Z(n524) );
  BUFFD0 U511 ( .I(n526), .Z(n525) );
  BUFFD0 U512 ( .I(n527), .Z(n526) );
  BUFFD0 U513 ( .I(n528), .Z(n527) );
  BUFFD0 U514 ( .I(n529), .Z(n528) );
  BUFFD0 U515 ( .I(n530), .Z(n529) );
  BUFFD0 U516 ( .I(n531), .Z(n530) );
  BUFFD0 U517 ( .I(n532), .Z(n531) );
  BUFFD0 U518 ( .I(n533), .Z(n532) );
  BUFFD0 U519 ( .I(n534), .Z(n533) );
  BUFFD0 U520 ( .I(n535), .Z(n534) );
  BUFFD0 U521 ( .I(n536), .Z(n535) );
  BUFFD0 U522 ( .I(n537), .Z(n536) );
  BUFFD0 U523 ( .I(n538), .Z(n537) );
  BUFFD0 U524 ( .I(n539), .Z(n538) );
  BUFFD0 U525 ( .I(n540), .Z(n539) );
  BUFFD0 U526 ( .I(n541), .Z(n540) );
  BUFFD0 U527 ( .I(n542), .Z(n541) );
  BUFFD0 U528 ( .I(n543), .Z(n542) );
  BUFFD0 U529 ( .I(n544), .Z(n543) );
  BUFFD0 U530 ( .I(n545), .Z(n544) );
  BUFFD0 U531 ( .I(n546), .Z(n545) );
  BUFFD0 U532 ( .I(n547), .Z(n546) );
  BUFFD0 U533 ( .I(n548), .Z(n547) );
  BUFFD0 U534 ( .I(n549), .Z(n548) );
  BUFFD0 U535 ( .I(DataOr[23]), .Z(n549) );
  BUFFD0 U536 ( .I(n551), .Z(n550) );
  BUFFD0 U537 ( .I(n552), .Z(n551) );
  BUFFD0 U538 ( .I(n553), .Z(n552) );
  BUFFD0 U539 ( .I(n554), .Z(n553) );
  BUFFD0 U540 ( .I(n555), .Z(n554) );
  BUFFD0 U541 ( .I(n556), .Z(n555) );
  BUFFD0 U542 ( .I(n557), .Z(n556) );
  BUFFD0 U543 ( .I(n558), .Z(n557) );
  BUFFD0 U544 ( .I(n559), .Z(n558) );
  BUFFD0 U545 ( .I(n560), .Z(n559) );
  BUFFD0 U546 ( .I(n561), .Z(n560) );
  BUFFD0 U547 ( .I(n562), .Z(n561) );
  BUFFD0 U548 ( .I(n563), .Z(n562) );
  BUFFD0 U549 ( .I(n564), .Z(n563) );
  BUFFD0 U550 ( .I(n565), .Z(n564) );
  BUFFD0 U551 ( .I(n566), .Z(n565) );
  BUFFD0 U552 ( .I(n567), .Z(n566) );
  BUFFD0 U553 ( .I(n568), .Z(n567) );
  BUFFD0 U554 ( .I(n569), .Z(n568) );
  BUFFD0 U555 ( .I(n570), .Z(n569) );
  BUFFD0 U556 ( .I(n571), .Z(n570) );
  BUFFD0 U557 ( .I(n572), .Z(n571) );
  BUFFD0 U558 ( .I(n573), .Z(n572) );
  BUFFD0 U559 ( .I(n574), .Z(n573) );
  BUFFD0 U560 ( .I(n575), .Z(n574) );
  BUFFD0 U561 ( .I(n576), .Z(n575) );
  BUFFD0 U562 ( .I(n577), .Z(n576) );
  BUFFD0 U563 ( .I(n578), .Z(n577) );
  BUFFD0 U564 ( .I(n579), .Z(n578) );
  BUFFD0 U565 ( .I(n580), .Z(n579) );
  BUFFD0 U566 ( .I(n581), .Z(n580) );
  BUFFD0 U567 ( .I(n582), .Z(n581) );
  BUFFD0 U568 ( .I(n583), .Z(n582) );
  BUFFD0 U569 ( .I(n584), .Z(n583) );
  BUFFD0 U570 ( .I(n585), .Z(n584) );
  BUFFD0 U571 ( .I(n586), .Z(n585) );
  BUFFD0 U572 ( .I(n587), .Z(n586) );
  BUFFD0 U573 ( .I(n588), .Z(n587) );
  BUFFD0 U574 ( .I(n589), .Z(n588) );
  BUFFD0 U575 ( .I(n590), .Z(n589) );
  BUFFD0 U576 ( .I(n591), .Z(n590) );
  BUFFD0 U577 ( .I(n592), .Z(n591) );
  BUFFD0 U578 ( .I(n593), .Z(n592) );
  BUFFD0 U579 ( .I(n594), .Z(n593) );
  BUFFD0 U580 ( .I(n595), .Z(n594) );
  BUFFD0 U581 ( .I(n596), .Z(n595) );
  BUFFD0 U582 ( .I(n597), .Z(n596) );
  BUFFD0 U583 ( .I(n598), .Z(n597) );
  BUFFD0 U584 ( .I(n599), .Z(n598) );
  BUFFD0 U585 ( .I(n600), .Z(n599) );
  BUFFD0 U586 ( .I(n601), .Z(n600) );
  BUFFD0 U587 ( .I(n602), .Z(n601) );
  BUFFD0 U588 ( .I(n603), .Z(n602) );
  BUFFD0 U589 ( .I(DataOr[22]), .Z(n603) );
  BUFFD0 U590 ( .I(n605), .Z(n604) );
  BUFFD0 U591 ( .I(n606), .Z(n605) );
  BUFFD0 U592 ( .I(n607), .Z(n606) );
  BUFFD0 U593 ( .I(n608), .Z(n607) );
  BUFFD0 U594 ( .I(n609), .Z(n608) );
  BUFFD0 U595 ( .I(n610), .Z(n609) );
  BUFFD0 U596 ( .I(n611), .Z(n610) );
  BUFFD0 U597 ( .I(n612), .Z(n611) );
  BUFFD0 U598 ( .I(n613), .Z(n612) );
  BUFFD0 U599 ( .I(n614), .Z(n613) );
  BUFFD0 U600 ( .I(n615), .Z(n614) );
  BUFFD0 U601 ( .I(n616), .Z(n615) );
  BUFFD0 U602 ( .I(n617), .Z(n616) );
  BUFFD0 U603 ( .I(n618), .Z(n617) );
  BUFFD0 U604 ( .I(n619), .Z(n618) );
  BUFFD0 U605 ( .I(n620), .Z(n619) );
  BUFFD0 U606 ( .I(n621), .Z(n620) );
  BUFFD0 U607 ( .I(n622), .Z(n621) );
  BUFFD0 U608 ( .I(n623), .Z(n622) );
  BUFFD0 U609 ( .I(n624), .Z(n623) );
  BUFFD0 U610 ( .I(n625), .Z(n624) );
  BUFFD0 U611 ( .I(n626), .Z(n625) );
  BUFFD0 U612 ( .I(n627), .Z(n626) );
  BUFFD0 U613 ( .I(n628), .Z(n627) );
  BUFFD0 U614 ( .I(n629), .Z(n628) );
  BUFFD0 U615 ( .I(n630), .Z(n629) );
  BUFFD0 U616 ( .I(n631), .Z(n630) );
  BUFFD0 U617 ( .I(n632), .Z(n631) );
  BUFFD0 U618 ( .I(n633), .Z(n632) );
  BUFFD0 U619 ( .I(n634), .Z(n633) );
  BUFFD0 U620 ( .I(n635), .Z(n634) );
  BUFFD0 U621 ( .I(n636), .Z(n635) );
  BUFFD0 U622 ( .I(n637), .Z(n636) );
  BUFFD0 U623 ( .I(n638), .Z(n637) );
  BUFFD0 U624 ( .I(n639), .Z(n638) );
  BUFFD0 U625 ( .I(n640), .Z(n639) );
  BUFFD0 U626 ( .I(n641), .Z(n640) );
  BUFFD0 U627 ( .I(n642), .Z(n641) );
  BUFFD0 U628 ( .I(n643), .Z(n642) );
  BUFFD0 U629 ( .I(n644), .Z(n643) );
  BUFFD0 U630 ( .I(n645), .Z(n644) );
  BUFFD0 U631 ( .I(n646), .Z(n645) );
  BUFFD0 U632 ( .I(n647), .Z(n646) );
  BUFFD0 U633 ( .I(n648), .Z(n647) );
  BUFFD0 U634 ( .I(n649), .Z(n648) );
  BUFFD0 U635 ( .I(n650), .Z(n649) );
  BUFFD0 U636 ( .I(n651), .Z(n650) );
  BUFFD0 U637 ( .I(n652), .Z(n651) );
  BUFFD0 U638 ( .I(n653), .Z(n652) );
  BUFFD0 U639 ( .I(n654), .Z(n653) );
  BUFFD0 U640 ( .I(n655), .Z(n654) );
  BUFFD0 U641 ( .I(n656), .Z(n655) );
  BUFFD0 U642 ( .I(n657), .Z(n656) );
  BUFFD0 U643 ( .I(DataOr[21]), .Z(n657) );
  BUFFD0 U644 ( .I(n659), .Z(n658) );
  BUFFD0 U645 ( .I(n660), .Z(n659) );
  BUFFD0 U646 ( .I(n661), .Z(n660) );
  BUFFD0 U647 ( .I(n662), .Z(n661) );
  BUFFD0 U648 ( .I(n663), .Z(n662) );
  BUFFD0 U649 ( .I(n664), .Z(n663) );
  BUFFD0 U650 ( .I(n665), .Z(n664) );
  BUFFD0 U651 ( .I(n666), .Z(n665) );
  BUFFD0 U652 ( .I(n667), .Z(n666) );
  BUFFD0 U653 ( .I(n668), .Z(n667) );
  BUFFD0 U654 ( .I(n669), .Z(n668) );
  BUFFD0 U655 ( .I(n670), .Z(n669) );
  BUFFD0 U656 ( .I(n671), .Z(n670) );
  BUFFD0 U657 ( .I(n672), .Z(n671) );
  BUFFD0 U658 ( .I(n673), .Z(n672) );
  BUFFD0 U659 ( .I(n674), .Z(n673) );
  BUFFD0 U660 ( .I(n675), .Z(n674) );
  BUFFD0 U661 ( .I(n676), .Z(n675) );
  BUFFD0 U662 ( .I(n677), .Z(n676) );
  BUFFD0 U663 ( .I(n678), .Z(n677) );
  BUFFD0 U664 ( .I(n679), .Z(n678) );
  BUFFD0 U665 ( .I(n680), .Z(n679) );
  BUFFD0 U666 ( .I(n681), .Z(n680) );
  BUFFD0 U667 ( .I(n682), .Z(n681) );
  BUFFD0 U668 ( .I(n683), .Z(n682) );
  BUFFD0 U669 ( .I(n684), .Z(n683) );
  BUFFD0 U670 ( .I(n685), .Z(n684) );
  BUFFD0 U671 ( .I(n686), .Z(n685) );
  BUFFD0 U672 ( .I(n687), .Z(n686) );
  BUFFD0 U673 ( .I(n688), .Z(n687) );
  BUFFD0 U674 ( .I(n689), .Z(n688) );
  BUFFD0 U675 ( .I(n690), .Z(n689) );
  BUFFD0 U676 ( .I(n691), .Z(n690) );
  BUFFD0 U677 ( .I(n692), .Z(n691) );
  BUFFD0 U678 ( .I(n693), .Z(n692) );
  BUFFD0 U679 ( .I(n694), .Z(n693) );
  BUFFD0 U680 ( .I(n695), .Z(n694) );
  BUFFD0 U681 ( .I(n696), .Z(n695) );
  BUFFD0 U682 ( .I(n697), .Z(n696) );
  BUFFD0 U683 ( .I(n698), .Z(n697) );
  BUFFD0 U684 ( .I(n699), .Z(n698) );
  BUFFD0 U685 ( .I(n700), .Z(n699) );
  BUFFD0 U686 ( .I(n701), .Z(n700) );
  BUFFD0 U687 ( .I(n702), .Z(n701) );
  BUFFD0 U688 ( .I(n703), .Z(n702) );
  BUFFD0 U689 ( .I(n704), .Z(n703) );
  BUFFD0 U690 ( .I(n705), .Z(n704) );
  BUFFD0 U691 ( .I(n706), .Z(n705) );
  BUFFD0 U692 ( .I(n707), .Z(n706) );
  BUFFD0 U693 ( .I(n708), .Z(n707) );
  BUFFD0 U694 ( .I(n709), .Z(n708) );
  BUFFD0 U695 ( .I(n710), .Z(n709) );
  BUFFD0 U696 ( .I(n711), .Z(n710) );
  BUFFD0 U697 ( .I(DataOr[20]), .Z(n711) );
  BUFFD0 U698 ( .I(n713), .Z(n712) );
  BUFFD0 U699 ( .I(n714), .Z(n713) );
  BUFFD0 U700 ( .I(n715), .Z(n714) );
  BUFFD0 U701 ( .I(n716), .Z(n715) );
  BUFFD0 U702 ( .I(n717), .Z(n716) );
  BUFFD0 U703 ( .I(n718), .Z(n717) );
  BUFFD0 U704 ( .I(n719), .Z(n718) );
  BUFFD0 U705 ( .I(n720), .Z(n719) );
  BUFFD0 U706 ( .I(n721), .Z(n720) );
  BUFFD0 U707 ( .I(n722), .Z(n721) );
  BUFFD0 U708 ( .I(n723), .Z(n722) );
  BUFFD0 U709 ( .I(n724), .Z(n723) );
  BUFFD0 U710 ( .I(n725), .Z(n724) );
  BUFFD0 U711 ( .I(n726), .Z(n725) );
  BUFFD0 U712 ( .I(n727), .Z(n726) );
  BUFFD0 U713 ( .I(n728), .Z(n727) );
  BUFFD0 U714 ( .I(n729), .Z(n728) );
  BUFFD0 U715 ( .I(n730), .Z(n729) );
  BUFFD0 U716 ( .I(n731), .Z(n730) );
  BUFFD0 U717 ( .I(n732), .Z(n731) );
  BUFFD0 U718 ( .I(n733), .Z(n732) );
  BUFFD0 U719 ( .I(n734), .Z(n733) );
  BUFFD0 U720 ( .I(n735), .Z(n734) );
  BUFFD0 U721 ( .I(n736), .Z(n735) );
  BUFFD0 U722 ( .I(n737), .Z(n736) );
  BUFFD0 U723 ( .I(n738), .Z(n737) );
  BUFFD0 U724 ( .I(n739), .Z(n738) );
  BUFFD0 U725 ( .I(n740), .Z(n739) );
  BUFFD0 U726 ( .I(n741), .Z(n740) );
  BUFFD0 U727 ( .I(n742), .Z(n741) );
  BUFFD0 U728 ( .I(n743), .Z(n742) );
  BUFFD0 U729 ( .I(n744), .Z(n743) );
  BUFFD0 U730 ( .I(n745), .Z(n744) );
  BUFFD0 U731 ( .I(n746), .Z(n745) );
  BUFFD0 U732 ( .I(n747), .Z(n746) );
  BUFFD0 U733 ( .I(n748), .Z(n747) );
  BUFFD0 U734 ( .I(n749), .Z(n748) );
  BUFFD0 U735 ( .I(n750), .Z(n749) );
  BUFFD0 U736 ( .I(n751), .Z(n750) );
  BUFFD0 U737 ( .I(n752), .Z(n751) );
  BUFFD0 U738 ( .I(n753), .Z(n752) );
  BUFFD0 U739 ( .I(n754), .Z(n753) );
  BUFFD0 U740 ( .I(n755), .Z(n754) );
  BUFFD0 U741 ( .I(n756), .Z(n755) );
  BUFFD0 U742 ( .I(n757), .Z(n756) );
  BUFFD0 U743 ( .I(n758), .Z(n757) );
  BUFFD0 U744 ( .I(n759), .Z(n758) );
  BUFFD0 U745 ( .I(n760), .Z(n759) );
  BUFFD0 U746 ( .I(n761), .Z(n760) );
  BUFFD0 U747 ( .I(n762), .Z(n761) );
  BUFFD0 U748 ( .I(n763), .Z(n762) );
  BUFFD0 U749 ( .I(n764), .Z(n763) );
  BUFFD0 U750 ( .I(n765), .Z(n764) );
  BUFFD0 U751 ( .I(DataOr[19]), .Z(n765) );
  BUFFD0 U752 ( .I(n767), .Z(n766) );
  BUFFD0 U753 ( .I(n768), .Z(n767) );
  BUFFD0 U754 ( .I(n769), .Z(n768) );
  BUFFD0 U755 ( .I(n770), .Z(n769) );
  BUFFD0 U756 ( .I(n771), .Z(n770) );
  BUFFD0 U757 ( .I(n772), .Z(n771) );
  BUFFD0 U758 ( .I(n773), .Z(n772) );
  BUFFD0 U759 ( .I(n774), .Z(n773) );
  BUFFD0 U760 ( .I(n775), .Z(n774) );
  BUFFD0 U761 ( .I(n776), .Z(n775) );
  BUFFD0 U762 ( .I(n777), .Z(n776) );
  BUFFD0 U763 ( .I(n778), .Z(n777) );
  BUFFD0 U764 ( .I(n779), .Z(n778) );
  BUFFD0 U765 ( .I(n780), .Z(n779) );
  BUFFD0 U766 ( .I(n781), .Z(n780) );
  BUFFD0 U767 ( .I(n782), .Z(n781) );
  BUFFD0 U768 ( .I(n783), .Z(n782) );
  BUFFD0 U769 ( .I(n784), .Z(n783) );
  BUFFD0 U770 ( .I(n785), .Z(n784) );
  BUFFD0 U771 ( .I(n786), .Z(n785) );
  BUFFD0 U772 ( .I(n787), .Z(n786) );
  BUFFD0 U773 ( .I(n788), .Z(n787) );
  BUFFD0 U774 ( .I(n789), .Z(n788) );
  BUFFD0 U775 ( .I(n790), .Z(n789) );
  BUFFD0 U776 ( .I(n791), .Z(n790) );
  BUFFD0 U777 ( .I(n792), .Z(n791) );
  BUFFD0 U778 ( .I(n793), .Z(n792) );
  BUFFD0 U779 ( .I(n794), .Z(n793) );
  BUFFD0 U780 ( .I(n795), .Z(n794) );
  BUFFD0 U781 ( .I(n796), .Z(n795) );
  BUFFD0 U782 ( .I(n797), .Z(n796) );
  BUFFD0 U783 ( .I(n798), .Z(n797) );
  BUFFD0 U784 ( .I(n799), .Z(n798) );
  BUFFD0 U785 ( .I(n800), .Z(n799) );
  BUFFD0 U786 ( .I(n801), .Z(n800) );
  BUFFD0 U787 ( .I(n802), .Z(n801) );
  BUFFD0 U788 ( .I(n803), .Z(n802) );
  BUFFD0 U789 ( .I(n804), .Z(n803) );
  BUFFD0 U790 ( .I(n805), .Z(n804) );
  BUFFD0 U791 ( .I(n806), .Z(n805) );
  BUFFD0 U792 ( .I(n807), .Z(n806) );
  BUFFD0 U793 ( .I(n808), .Z(n807) );
  BUFFD0 U794 ( .I(n809), .Z(n808) );
  BUFFD0 U795 ( .I(n810), .Z(n809) );
  BUFFD0 U796 ( .I(n811), .Z(n810) );
  BUFFD0 U797 ( .I(n812), .Z(n811) );
  BUFFD0 U798 ( .I(n813), .Z(n812) );
  BUFFD0 U799 ( .I(n814), .Z(n813) );
  BUFFD0 U800 ( .I(n815), .Z(n814) );
  BUFFD0 U801 ( .I(n816), .Z(n815) );
  BUFFD0 U802 ( .I(n817), .Z(n816) );
  BUFFD0 U803 ( .I(n818), .Z(n817) );
  BUFFD0 U804 ( .I(n819), .Z(n818) );
  BUFFD0 U805 ( .I(DataOr[18]), .Z(n819) );
  BUFFD0 U806 ( .I(n821), .Z(n820) );
  BUFFD0 U807 ( .I(n822), .Z(n821) );
  BUFFD0 U808 ( .I(n823), .Z(n822) );
  BUFFD0 U809 ( .I(n824), .Z(n823) );
  BUFFD0 U810 ( .I(n825), .Z(n824) );
  BUFFD0 U811 ( .I(n826), .Z(n825) );
  BUFFD0 U812 ( .I(n827), .Z(n826) );
  BUFFD0 U813 ( .I(n828), .Z(n827) );
  BUFFD0 U814 ( .I(n829), .Z(n828) );
  BUFFD0 U815 ( .I(n830), .Z(n829) );
  BUFFD0 U816 ( .I(n831), .Z(n830) );
  BUFFD0 U817 ( .I(n832), .Z(n831) );
  BUFFD0 U818 ( .I(n833), .Z(n832) );
  BUFFD0 U819 ( .I(n834), .Z(n833) );
  BUFFD0 U820 ( .I(n835), .Z(n834) );
  BUFFD0 U821 ( .I(n836), .Z(n835) );
  BUFFD0 U822 ( .I(n837), .Z(n836) );
  BUFFD0 U823 ( .I(n838), .Z(n837) );
  BUFFD0 U824 ( .I(n839), .Z(n838) );
  BUFFD0 U825 ( .I(n840), .Z(n839) );
  BUFFD0 U826 ( .I(n841), .Z(n840) );
  BUFFD0 U827 ( .I(n842), .Z(n841) );
  BUFFD0 U828 ( .I(n843), .Z(n842) );
  BUFFD0 U829 ( .I(n844), .Z(n843) );
  BUFFD0 U830 ( .I(n845), .Z(n844) );
  BUFFD0 U831 ( .I(n846), .Z(n845) );
  BUFFD0 U832 ( .I(n847), .Z(n846) );
  BUFFD0 U833 ( .I(n848), .Z(n847) );
  BUFFD0 U834 ( .I(n849), .Z(n848) );
  BUFFD0 U835 ( .I(n850), .Z(n849) );
  BUFFD0 U836 ( .I(n851), .Z(n850) );
  BUFFD0 U837 ( .I(n852), .Z(n851) );
  BUFFD0 U838 ( .I(n853), .Z(n852) );
  BUFFD0 U839 ( .I(n854), .Z(n853) );
  BUFFD0 U840 ( .I(n855), .Z(n854) );
  BUFFD0 U841 ( .I(n856), .Z(n855) );
  BUFFD0 U842 ( .I(n857), .Z(n856) );
  BUFFD0 U843 ( .I(n858), .Z(n857) );
  BUFFD0 U844 ( .I(n859), .Z(n858) );
  BUFFD0 U845 ( .I(n860), .Z(n859) );
  BUFFD0 U846 ( .I(n861), .Z(n860) );
  BUFFD0 U847 ( .I(n862), .Z(n861) );
  BUFFD0 U848 ( .I(n863), .Z(n862) );
  BUFFD0 U849 ( .I(n864), .Z(n863) );
  BUFFD0 U850 ( .I(n865), .Z(n864) );
  BUFFD0 U851 ( .I(n866), .Z(n865) );
  BUFFD0 U852 ( .I(n867), .Z(n866) );
  BUFFD0 U853 ( .I(n868), .Z(n867) );
  BUFFD0 U854 ( .I(n869), .Z(n868) );
  BUFFD0 U855 ( .I(n870), .Z(n869) );
  BUFFD0 U856 ( .I(n871), .Z(n870) );
  BUFFD0 U857 ( .I(n872), .Z(n871) );
  BUFFD0 U858 ( .I(n873), .Z(n872) );
  BUFFD0 U859 ( .I(DataOr[17]), .Z(n873) );
  BUFFD0 U860 ( .I(n875), .Z(n874) );
  BUFFD0 U861 ( .I(n876), .Z(n875) );
  BUFFD0 U862 ( .I(n877), .Z(n876) );
  BUFFD0 U863 ( .I(n878), .Z(n877) );
  BUFFD0 U864 ( .I(n879), .Z(n878) );
  BUFFD0 U865 ( .I(n880), .Z(n879) );
  BUFFD0 U866 ( .I(n881), .Z(n880) );
  BUFFD0 U867 ( .I(n882), .Z(n881) );
  BUFFD0 U868 ( .I(n883), .Z(n882) );
  BUFFD0 U869 ( .I(n884), .Z(n883) );
  BUFFD0 U870 ( .I(n885), .Z(n884) );
  BUFFD0 U871 ( .I(n886), .Z(n885) );
  BUFFD0 U872 ( .I(n887), .Z(n886) );
  BUFFD0 U873 ( .I(n888), .Z(n887) );
  BUFFD0 U874 ( .I(n889), .Z(n888) );
  BUFFD0 U875 ( .I(n890), .Z(n889) );
  BUFFD0 U876 ( .I(n891), .Z(n890) );
  BUFFD0 U877 ( .I(n892), .Z(n891) );
  BUFFD0 U878 ( .I(n893), .Z(n892) );
  BUFFD0 U879 ( .I(n894), .Z(n893) );
  BUFFD0 U880 ( .I(n895), .Z(n894) );
  BUFFD0 U881 ( .I(n896), .Z(n895) );
  BUFFD0 U882 ( .I(n897), .Z(n896) );
  BUFFD0 U883 ( .I(n898), .Z(n897) );
  BUFFD0 U884 ( .I(n899), .Z(n898) );
  BUFFD0 U885 ( .I(n900), .Z(n899) );
  BUFFD0 U886 ( .I(n901), .Z(n900) );
  BUFFD0 U887 ( .I(n902), .Z(n901) );
  BUFFD0 U888 ( .I(n903), .Z(n902) );
  BUFFD0 U889 ( .I(n904), .Z(n903) );
  BUFFD0 U890 ( .I(n905), .Z(n904) );
  BUFFD0 U891 ( .I(n906), .Z(n905) );
  BUFFD0 U892 ( .I(n907), .Z(n906) );
  BUFFD0 U893 ( .I(n908), .Z(n907) );
  BUFFD0 U894 ( .I(n909), .Z(n908) );
  BUFFD0 U895 ( .I(n910), .Z(n909) );
  BUFFD0 U896 ( .I(n911), .Z(n910) );
  BUFFD0 U897 ( .I(n912), .Z(n911) );
  BUFFD0 U898 ( .I(n913), .Z(n912) );
  BUFFD0 U899 ( .I(n914), .Z(n913) );
  BUFFD0 U900 ( .I(n915), .Z(n914) );
  BUFFD0 U901 ( .I(n916), .Z(n915) );
  BUFFD0 U902 ( .I(n917), .Z(n916) );
  BUFFD0 U903 ( .I(n918), .Z(n917) );
  BUFFD0 U904 ( .I(n919), .Z(n918) );
  BUFFD0 U905 ( .I(n920), .Z(n919) );
  BUFFD0 U906 ( .I(n921), .Z(n920) );
  BUFFD0 U907 ( .I(n922), .Z(n921) );
  BUFFD0 U908 ( .I(n923), .Z(n922) );
  BUFFD0 U909 ( .I(n924), .Z(n923) );
  BUFFD0 U910 ( .I(n925), .Z(n924) );
  BUFFD0 U911 ( .I(n926), .Z(n925) );
  BUFFD0 U912 ( .I(n927), .Z(n926) );
  BUFFD0 U913 ( .I(DataOr[16]), .Z(n927) );
  BUFFD0 U914 ( .I(n929), .Z(n928) );
  BUFFD0 U915 ( .I(n930), .Z(n929) );
  BUFFD0 U916 ( .I(n931), .Z(n930) );
  BUFFD0 U917 ( .I(n932), .Z(n931) );
  BUFFD0 U918 ( .I(n933), .Z(n932) );
  BUFFD0 U919 ( .I(n934), .Z(n933) );
  BUFFD0 U920 ( .I(n935), .Z(n934) );
  BUFFD0 U921 ( .I(n936), .Z(n935) );
  BUFFD0 U922 ( .I(n937), .Z(n936) );
  BUFFD0 U923 ( .I(n938), .Z(n937) );
  BUFFD0 U924 ( .I(n939), .Z(n938) );
  BUFFD0 U925 ( .I(n940), .Z(n939) );
  BUFFD0 U926 ( .I(n941), .Z(n940) );
  BUFFD0 U927 ( .I(n942), .Z(n941) );
  BUFFD0 U928 ( .I(n943), .Z(n942) );
  BUFFD0 U929 ( .I(n944), .Z(n943) );
  BUFFD0 U930 ( .I(n945), .Z(n944) );
  BUFFD0 U931 ( .I(n946), .Z(n945) );
  BUFFD0 U932 ( .I(n947), .Z(n946) );
  BUFFD0 U933 ( .I(n948), .Z(n947) );
  BUFFD0 U934 ( .I(n949), .Z(n948) );
  BUFFD0 U935 ( .I(n950), .Z(n949) );
  BUFFD0 U936 ( .I(n951), .Z(n950) );
  BUFFD0 U937 ( .I(n952), .Z(n951) );
  BUFFD0 U938 ( .I(n953), .Z(n952) );
  BUFFD0 U939 ( .I(n954), .Z(n953) );
  BUFFD0 U940 ( .I(n955), .Z(n954) );
  BUFFD0 U941 ( .I(n956), .Z(n955) );
  BUFFD0 U942 ( .I(n957), .Z(n956) );
  BUFFD0 U943 ( .I(n958), .Z(n957) );
  BUFFD0 U944 ( .I(n959), .Z(n958) );
  BUFFD0 U945 ( .I(n960), .Z(n959) );
  BUFFD0 U946 ( .I(n961), .Z(n960) );
  BUFFD0 U947 ( .I(n962), .Z(n961) );
  BUFFD0 U948 ( .I(n963), .Z(n962) );
  BUFFD0 U949 ( .I(n964), .Z(n963) );
  BUFFD0 U950 ( .I(n965), .Z(n964) );
  BUFFD0 U951 ( .I(n966), .Z(n965) );
  BUFFD0 U952 ( .I(n967), .Z(n966) );
  BUFFD0 U953 ( .I(n968), .Z(n967) );
  BUFFD0 U954 ( .I(n969), .Z(n968) );
  BUFFD0 U955 ( .I(n970), .Z(n969) );
  BUFFD0 U956 ( .I(n971), .Z(n970) );
  BUFFD0 U957 ( .I(n972), .Z(n971) );
  BUFFD0 U958 ( .I(n973), .Z(n972) );
  BUFFD0 U959 ( .I(n974), .Z(n973) );
  BUFFD0 U960 ( .I(n975), .Z(n974) );
  BUFFD0 U961 ( .I(n976), .Z(n975) );
  BUFFD0 U962 ( .I(n977), .Z(n976) );
  BUFFD0 U963 ( .I(n978), .Z(n977) );
  BUFFD0 U964 ( .I(n979), .Z(n978) );
  BUFFD0 U965 ( .I(n980), .Z(n979) );
  BUFFD0 U966 ( .I(n981), .Z(n980) );
  BUFFD0 U967 ( .I(DataOr[15]), .Z(n981) );
  BUFFD0 U968 ( .I(n983), .Z(n982) );
  BUFFD0 U969 ( .I(n984), .Z(n983) );
  BUFFD0 U970 ( .I(n985), .Z(n984) );
  BUFFD0 U971 ( .I(n986), .Z(n985) );
  BUFFD0 U972 ( .I(n987), .Z(n986) );
  BUFFD0 U973 ( .I(n988), .Z(n987) );
  BUFFD0 U974 ( .I(n989), .Z(n988) );
  BUFFD0 U975 ( .I(n990), .Z(n989) );
  BUFFD0 U976 ( .I(n991), .Z(n990) );
  BUFFD0 U977 ( .I(n992), .Z(n991) );
  BUFFD0 U978 ( .I(n993), .Z(n992) );
  BUFFD0 U979 ( .I(n994), .Z(n993) );
  BUFFD0 U980 ( .I(n995), .Z(n994) );
  BUFFD0 U981 ( .I(n996), .Z(n995) );
  BUFFD0 U982 ( .I(n997), .Z(n996) );
  BUFFD0 U983 ( .I(n998), .Z(n997) );
  BUFFD0 U984 ( .I(n999), .Z(n998) );
  BUFFD0 U985 ( .I(n1000), .Z(n999) );
  BUFFD0 U986 ( .I(n1001), .Z(n1000) );
  BUFFD0 U987 ( .I(n1002), .Z(n1001) );
  BUFFD0 U988 ( .I(n1003), .Z(n1002) );
  BUFFD0 U989 ( .I(n1004), .Z(n1003) );
  BUFFD0 U990 ( .I(n1005), .Z(n1004) );
  BUFFD0 U991 ( .I(n1006), .Z(n1005) );
  BUFFD0 U992 ( .I(n1007), .Z(n1006) );
  BUFFD0 U993 ( .I(n1008), .Z(n1007) );
  BUFFD0 U994 ( .I(n1009), .Z(n1008) );
  BUFFD0 U995 ( .I(n1010), .Z(n1009) );
  BUFFD0 U996 ( .I(n1011), .Z(n1010) );
  BUFFD0 U997 ( .I(n1012), .Z(n1011) );
  BUFFD0 U998 ( .I(n1013), .Z(n1012) );
  BUFFD0 U999 ( .I(n1014), .Z(n1013) );
  BUFFD0 U1000 ( .I(n1015), .Z(n1014) );
  BUFFD0 U1001 ( .I(n1016), .Z(n1015) );
  BUFFD0 U1002 ( .I(n1017), .Z(n1016) );
  BUFFD0 U1003 ( .I(n1018), .Z(n1017) );
  BUFFD0 U1004 ( .I(n1019), .Z(n1018) );
  BUFFD0 U1005 ( .I(n1020), .Z(n1019) );
  BUFFD0 U1006 ( .I(n1021), .Z(n1020) );
  BUFFD0 U1007 ( .I(n1022), .Z(n1021) );
  BUFFD0 U1008 ( .I(n1023), .Z(n1022) );
  BUFFD0 U1009 ( .I(n1024), .Z(n1023) );
  BUFFD0 U1010 ( .I(n1025), .Z(n1024) );
  BUFFD0 U1011 ( .I(n1026), .Z(n1025) );
  BUFFD0 U1012 ( .I(n1027), .Z(n1026) );
  BUFFD0 U1013 ( .I(n1028), .Z(n1027) );
  BUFFD0 U1014 ( .I(n1029), .Z(n1028) );
  BUFFD0 U1015 ( .I(n1030), .Z(n1029) );
  BUFFD0 U1016 ( .I(n1031), .Z(n1030) );
  BUFFD0 U1017 ( .I(n1032), .Z(n1031) );
  BUFFD0 U1018 ( .I(n1033), .Z(n1032) );
  BUFFD0 U1019 ( .I(n1034), .Z(n1033) );
  BUFFD0 U1020 ( .I(n1035), .Z(n1034) );
  BUFFD0 U1021 ( .I(DataOr[14]), .Z(n1035) );
  BUFFD0 U1022 ( .I(n1037), .Z(n1036) );
  BUFFD0 U1023 ( .I(n1038), .Z(n1037) );
  BUFFD0 U1024 ( .I(n1039), .Z(n1038) );
  BUFFD0 U1025 ( .I(n1040), .Z(n1039) );
  BUFFD0 U1026 ( .I(n1041), .Z(n1040) );
  BUFFD0 U1027 ( .I(n1042), .Z(n1041) );
  BUFFD0 U1028 ( .I(n1043), .Z(n1042) );
  BUFFD0 U1029 ( .I(n1044), .Z(n1043) );
  BUFFD0 U1030 ( .I(n1045), .Z(n1044) );
  BUFFD0 U1031 ( .I(n1046), .Z(n1045) );
  BUFFD0 U1032 ( .I(n1047), .Z(n1046) );
  BUFFD0 U1033 ( .I(n1048), .Z(n1047) );
  BUFFD0 U1034 ( .I(n1049), .Z(n1048) );
  BUFFD0 U1035 ( .I(n1050), .Z(n1049) );
  BUFFD0 U1036 ( .I(n1051), .Z(n1050) );
  BUFFD0 U1037 ( .I(n1052), .Z(n1051) );
  BUFFD0 U1038 ( .I(n1053), .Z(n1052) );
  BUFFD0 U1039 ( .I(n1054), .Z(n1053) );
  BUFFD0 U1040 ( .I(n1055), .Z(n1054) );
  BUFFD0 U1041 ( .I(n1056), .Z(n1055) );
  BUFFD0 U1042 ( .I(n1057), .Z(n1056) );
  BUFFD0 U1043 ( .I(n1058), .Z(n1057) );
  BUFFD0 U1044 ( .I(n1059), .Z(n1058) );
  BUFFD0 U1045 ( .I(n1060), .Z(n1059) );
  BUFFD0 U1046 ( .I(n1061), .Z(n1060) );
  BUFFD0 U1047 ( .I(n1062), .Z(n1061) );
  BUFFD0 U1048 ( .I(n1063), .Z(n1062) );
  BUFFD0 U1049 ( .I(n1064), .Z(n1063) );
  BUFFD0 U1050 ( .I(n1065), .Z(n1064) );
  BUFFD0 U1051 ( .I(n1066), .Z(n1065) );
  BUFFD0 U1052 ( .I(n1067), .Z(n1066) );
  BUFFD0 U1053 ( .I(n1068), .Z(n1067) );
  BUFFD0 U1054 ( .I(n1069), .Z(n1068) );
  BUFFD0 U1055 ( .I(n1070), .Z(n1069) );
  BUFFD0 U1056 ( .I(n1071), .Z(n1070) );
  BUFFD0 U1057 ( .I(n1072), .Z(n1071) );
  BUFFD0 U1058 ( .I(n1073), .Z(n1072) );
  BUFFD0 U1059 ( .I(n1074), .Z(n1073) );
  BUFFD0 U1060 ( .I(n1075), .Z(n1074) );
  BUFFD0 U1061 ( .I(n1076), .Z(n1075) );
  BUFFD0 U1062 ( .I(n1077), .Z(n1076) );
  BUFFD0 U1063 ( .I(n1078), .Z(n1077) );
  BUFFD0 U1064 ( .I(n1079), .Z(n1078) );
  BUFFD0 U1065 ( .I(n1080), .Z(n1079) );
  BUFFD0 U1066 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1067 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1068 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1069 ( .I(n1084), .Z(n1083) );
  BUFFD0 U1070 ( .I(n1085), .Z(n1084) );
  BUFFD0 U1071 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1072 ( .I(n1087), .Z(n1086) );
  BUFFD0 U1073 ( .I(n1088), .Z(n1087) );
  BUFFD0 U1074 ( .I(n1089), .Z(n1088) );
  BUFFD0 U1075 ( .I(DataOr[13]), .Z(n1089) );
  BUFFD0 U1076 ( .I(n1091), .Z(n1090) );
  BUFFD0 U1077 ( .I(n1092), .Z(n1091) );
  BUFFD0 U1078 ( .I(n1093), .Z(n1092) );
  BUFFD0 U1079 ( .I(n1094), .Z(n1093) );
  BUFFD0 U1080 ( .I(n1095), .Z(n1094) );
  BUFFD0 U1081 ( .I(n1096), .Z(n1095) );
  BUFFD0 U1082 ( .I(n1097), .Z(n1096) );
  BUFFD0 U1083 ( .I(n1098), .Z(n1097) );
  BUFFD0 U1084 ( .I(n1099), .Z(n1098) );
  BUFFD0 U1085 ( .I(n1100), .Z(n1099) );
  BUFFD0 U1086 ( .I(n1101), .Z(n1100) );
  BUFFD0 U1087 ( .I(n1102), .Z(n1101) );
  BUFFD0 U1088 ( .I(n1103), .Z(n1102) );
  BUFFD0 U1089 ( .I(n1104), .Z(n1103) );
  BUFFD0 U1090 ( .I(n1105), .Z(n1104) );
  BUFFD0 U1091 ( .I(n1106), .Z(n1105) );
  BUFFD0 U1092 ( .I(n1107), .Z(n1106) );
  BUFFD0 U1093 ( .I(n1108), .Z(n1107) );
  BUFFD0 U1094 ( .I(n1109), .Z(n1108) );
  BUFFD0 U1095 ( .I(n1110), .Z(n1109) );
  BUFFD0 U1096 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1097 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1098 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1099 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1100 ( .I(n1115), .Z(n1114) );
  BUFFD0 U1101 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1102 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1103 ( .I(n1118), .Z(n1117) );
  BUFFD0 U1104 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1105 ( .I(n1120), .Z(n1119) );
  BUFFD0 U1106 ( .I(n1121), .Z(n1120) );
  BUFFD0 U1107 ( .I(n1122), .Z(n1121) );
  BUFFD0 U1108 ( .I(n1123), .Z(n1122) );
  BUFFD0 U1109 ( .I(n1124), .Z(n1123) );
  BUFFD0 U1110 ( .I(n1125), .Z(n1124) );
  BUFFD0 U1111 ( .I(n1126), .Z(n1125) );
  BUFFD0 U1112 ( .I(n1127), .Z(n1126) );
  BUFFD0 U1113 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1114 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1115 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1116 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1117 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1118 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1119 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1120 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1121 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1122 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1123 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1124 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1125 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1126 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1127 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1128 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1129 ( .I(DataOr[12]), .Z(n1143) );
  BUFFD0 U1130 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1131 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1132 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1133 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1134 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1135 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1136 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1137 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1138 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1139 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1140 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1141 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1142 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1143 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1144 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1145 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1146 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1147 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1148 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1149 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1150 ( .I(n1165), .Z(n1164) );
  BUFFD0 U1151 ( .I(n1166), .Z(n1165) );
  BUFFD0 U1152 ( .I(n1167), .Z(n1166) );
  BUFFD0 U1153 ( .I(n1168), .Z(n1167) );
  BUFFD0 U1154 ( .I(n1169), .Z(n1168) );
  BUFFD0 U1155 ( .I(n1170), .Z(n1169) );
  BUFFD0 U1156 ( .I(n1171), .Z(n1170) );
  BUFFD0 U1157 ( .I(n1172), .Z(n1171) );
  BUFFD0 U1158 ( .I(n1173), .Z(n1172) );
  BUFFD0 U1159 ( .I(n1174), .Z(n1173) );
  BUFFD0 U1160 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1161 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1162 ( .I(n1177), .Z(n1176) );
  BUFFD0 U1163 ( .I(n1178), .Z(n1177) );
  BUFFD0 U1164 ( .I(n1179), .Z(n1178) );
  BUFFD0 U1165 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1166 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1167 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1168 ( .I(n1183), .Z(n1182) );
  BUFFD0 U1169 ( .I(n1184), .Z(n1183) );
  BUFFD0 U1170 ( .I(n1185), .Z(n1184) );
  BUFFD0 U1171 ( .I(n1186), .Z(n1185) );
  BUFFD0 U1172 ( .I(n1187), .Z(n1186) );
  BUFFD0 U1173 ( .I(n1188), .Z(n1187) );
  BUFFD0 U1174 ( .I(n1189), .Z(n1188) );
  BUFFD0 U1175 ( .I(n1190), .Z(n1189) );
  BUFFD0 U1176 ( .I(n1191), .Z(n1190) );
  BUFFD0 U1177 ( .I(n1192), .Z(n1191) );
  BUFFD0 U1178 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1179 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1180 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1181 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1182 ( .I(n1197), .Z(n1196) );
  BUFFD0 U1183 ( .I(DataOr[11]), .Z(n1197) );
  BUFFD0 U1184 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1185 ( .I(n1200), .Z(n1199) );
  BUFFD0 U1186 ( .I(n1201), .Z(n1200) );
  BUFFD0 U1187 ( .I(n1202), .Z(n1201) );
  BUFFD0 U1188 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1189 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1190 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1191 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1192 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1193 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1194 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1195 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1196 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1197 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1198 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1199 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1200 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1201 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1202 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1203 ( .I(n1218), .Z(n1217) );
  BUFFD0 U1204 ( .I(n1219), .Z(n1218) );
  BUFFD0 U1205 ( .I(n1220), .Z(n1219) );
  BUFFD0 U1206 ( .I(n1221), .Z(n1220) );
  BUFFD0 U1207 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1208 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1209 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1210 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1211 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1212 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1213 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1214 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1215 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1216 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1217 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1218 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1219 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1220 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1221 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1222 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1223 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1224 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1225 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1226 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1227 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1228 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1229 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1230 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1231 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1232 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1233 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1234 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1235 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1236 ( .I(n1251), .Z(n1250) );
  BUFFD0 U1237 ( .I(DataOr[10]), .Z(n1251) );
  BUFFD0 U1238 ( .I(n1253), .Z(n1252) );
  BUFFD0 U1239 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1240 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1241 ( .I(n1256), .Z(n1255) );
  BUFFD0 U1242 ( .I(n1257), .Z(n1256) );
  BUFFD0 U1243 ( .I(n1258), .Z(n1257) );
  BUFFD0 U1244 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1245 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1246 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1247 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1248 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1249 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1250 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1251 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1252 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1253 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1254 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1255 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1256 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1257 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1258 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1259 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1260 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1261 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1262 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1263 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1264 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1265 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1266 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1267 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1268 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1269 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1270 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1271 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1272 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1273 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1274 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1275 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1276 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1277 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1278 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1279 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1280 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1281 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1282 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1283 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1284 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1285 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1286 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1287 ( .I(n1302), .Z(n1301) );
  BUFFD0 U1288 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1289 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1290 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1291 ( .I(DataOr[9]), .Z(n1305) );
  BUFFD0 U1292 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1293 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1294 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1295 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1296 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1297 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1298 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1299 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1300 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1301 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1302 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1303 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1304 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1305 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1306 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1307 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1308 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1309 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1310 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1311 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1312 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1313 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1314 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1315 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1316 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1317 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1318 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1319 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1320 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1321 ( .I(n1336), .Z(n1335) );
  BUFFD0 U1322 ( .I(n1337), .Z(n1336) );
  BUFFD0 U1323 ( .I(n1338), .Z(n1337) );
  BUFFD0 U1324 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1325 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1326 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1327 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1328 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1329 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1330 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1331 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1332 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1333 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1334 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1335 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1336 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1337 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1338 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1339 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1340 ( .I(n1355), .Z(n1354) );
  BUFFD0 U1341 ( .I(n1356), .Z(n1355) );
  BUFFD0 U1342 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1343 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1344 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1345 ( .I(DataOr[8]), .Z(n1359) );
  BUFFD0 U1346 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1347 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1348 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1349 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1350 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1351 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1352 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1353 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1354 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1355 ( .I(n1370), .Z(n1369) );
  BUFFD0 U1356 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1357 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1358 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1359 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1360 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1361 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1362 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1363 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1364 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1365 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1366 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1367 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1368 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1369 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1370 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1371 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1372 ( .I(n1387), .Z(n1386) );
  BUFFD0 U1373 ( .I(n1388), .Z(n1387) );
  BUFFD0 U1374 ( .I(n1389), .Z(n1388) );
  BUFFD0 U1375 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1376 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1377 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1378 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1379 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1380 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1381 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1382 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1383 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1384 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1385 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1386 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1387 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1388 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1389 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1390 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1391 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1392 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1393 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1394 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1395 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1396 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1397 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1398 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1399 ( .I(DataOr[7]), .Z(n1413) );
  BUFFD0 U1400 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1401 ( .I(n1416), .Z(n1415) );
  BUFFD0 U1402 ( .I(n1417), .Z(n1416) );
  BUFFD0 U1403 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1404 ( .I(n1419), .Z(n1418) );
  BUFFD0 U1405 ( .I(n1420), .Z(n1419) );
  BUFFD0 U1406 ( .I(n1421), .Z(n1420) );
  BUFFD0 U1407 ( .I(n1422), .Z(n1421) );
  BUFFD0 U1408 ( .I(n1423), .Z(n1422) );
  BUFFD0 U1409 ( .I(n1424), .Z(n1423) );
  BUFFD0 U1410 ( .I(n1425), .Z(n1424) );
  BUFFD0 U1411 ( .I(n1426), .Z(n1425) );
  BUFFD0 U1412 ( .I(n1427), .Z(n1426) );
  BUFFD0 U1413 ( .I(n1428), .Z(n1427) );
  BUFFD0 U1414 ( .I(n1429), .Z(n1428) );
  BUFFD0 U1415 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1416 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1417 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1418 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1419 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1420 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1421 ( .I(n1436), .Z(n1435) );
  BUFFD0 U1422 ( .I(n1437), .Z(n1436) );
  BUFFD0 U1423 ( .I(n1438), .Z(n1437) );
  BUFFD0 U1424 ( .I(n1439), .Z(n1438) );
  BUFFD0 U1425 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1426 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1427 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1428 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1429 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1430 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1431 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1432 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1433 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1434 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1435 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1436 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1437 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1438 ( .I(n1453), .Z(n1452) );
  BUFFD0 U1439 ( .I(n1454), .Z(n1453) );
  BUFFD0 U1440 ( .I(n1455), .Z(n1454) );
  BUFFD0 U1441 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1442 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1443 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1444 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1445 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1446 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1447 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1448 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1449 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1450 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1451 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1452 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1453 ( .I(DataOr[6]), .Z(n1467) );
  BUFFD0 U1454 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1455 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1456 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1457 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1458 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1459 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1460 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1461 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1462 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1463 ( .I(n1478), .Z(n1477) );
  BUFFD0 U1464 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1465 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1466 ( .I(n1481), .Z(n1480) );
  BUFFD0 U1467 ( .I(n1482), .Z(n1481) );
  BUFFD0 U1468 ( .I(n1483), .Z(n1482) );
  BUFFD0 U1469 ( .I(n1484), .Z(n1483) );
  BUFFD0 U1470 ( .I(n1485), .Z(n1484) );
  BUFFD0 U1471 ( .I(n1486), .Z(n1485) );
  BUFFD0 U1472 ( .I(n1487), .Z(n1486) );
  BUFFD0 U1473 ( .I(n1488), .Z(n1487) );
  BUFFD0 U1474 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1475 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1476 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1477 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1478 ( .I(n1493), .Z(n1492) );
  BUFFD0 U1479 ( .I(n1494), .Z(n1493) );
  BUFFD0 U1480 ( .I(n1495), .Z(n1494) );
  BUFFD0 U1481 ( .I(n1496), .Z(n1495) );
  BUFFD0 U1482 ( .I(n1497), .Z(n1496) );
  BUFFD0 U1483 ( .I(n1498), .Z(n1497) );
  BUFFD0 U1484 ( .I(n1499), .Z(n1498) );
  BUFFD0 U1485 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1486 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1487 ( .I(n1502), .Z(n1501) );
  BUFFD0 U1488 ( .I(n1503), .Z(n1502) );
  BUFFD0 U1489 ( .I(n1504), .Z(n1503) );
  BUFFD0 U1490 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1491 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1492 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1493 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1494 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1495 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1496 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1497 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1498 ( .I(n1513), .Z(n1512) );
  BUFFD0 U1499 ( .I(n1514), .Z(n1513) );
  BUFFD0 U1500 ( .I(n1515), .Z(n1514) );
  BUFFD0 U1501 ( .I(n1516), .Z(n1515) );
  BUFFD0 U1502 ( .I(n1517), .Z(n1516) );
  BUFFD0 U1503 ( .I(n1518), .Z(n1517) );
  BUFFD0 U1504 ( .I(n1519), .Z(n1518) );
  BUFFD0 U1505 ( .I(n1520), .Z(n1519) );
  BUFFD0 U1506 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1507 ( .I(DataOr[5]), .Z(n1521) );
  BUFFD0 U1508 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1509 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1510 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1511 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1512 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1513 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1514 ( .I(n1529), .Z(n1528) );
  BUFFD0 U1515 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1516 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1517 ( .I(n1532), .Z(n1531) );
  BUFFD0 U1518 ( .I(n1533), .Z(n1532) );
  BUFFD0 U1519 ( .I(n1534), .Z(n1533) );
  BUFFD0 U1520 ( .I(n1535), .Z(n1534) );
  BUFFD0 U1521 ( .I(n1536), .Z(n1535) );
  BUFFD0 U1522 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1523 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1524 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1525 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1526 ( .I(n1541), .Z(n1540) );
  BUFFD0 U1527 ( .I(n1542), .Z(n1541) );
  BUFFD0 U1528 ( .I(n1543), .Z(n1542) );
  BUFFD0 U1529 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1530 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1531 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1532 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1533 ( .I(n1548), .Z(n1547) );
  BUFFD0 U1534 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1535 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1536 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1537 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1538 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1539 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1540 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1541 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1542 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1543 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1544 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1545 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1546 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1547 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1548 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1549 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1550 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1551 ( .I(n1566), .Z(n1565) );
  BUFFD0 U1552 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1553 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1554 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1555 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1556 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1557 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1558 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1559 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1560 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1561 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1562 ( .I(DataOr[4]), .Z(n1576) );
  BUFFD0 U1563 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1564 ( .I(n1579), .Z(n1578) );
  BUFFD0 U1565 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1566 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1567 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1568 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1569 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1570 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1571 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1572 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1573 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1574 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1575 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1576 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1577 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1578 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1579 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1580 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1581 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1582 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1583 ( .I(n1598), .Z(n1597) );
  BUFFD0 U1584 ( .I(n1599), .Z(n1598) );
  BUFFD0 U1585 ( .I(n1600), .Z(n1599) );
  BUFFD0 U1586 ( .I(n1601), .Z(n1600) );
  BUFFD0 U1587 ( .I(n1602), .Z(n1601) );
  BUFFD0 U1588 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1589 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1590 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1591 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1592 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1593 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1594 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1595 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1596 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1597 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1598 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1599 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1600 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1601 ( .I(n1616), .Z(n1615) );
  BUFFD0 U1602 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1603 ( .I(n1618), .Z(n1617) );
  BUFFD0 U1604 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1605 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1606 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1607 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1608 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1609 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1610 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1611 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1612 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1613 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1614 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1615 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1616 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1617 ( .I(DataOr[3]), .Z(n1631) );
  BUFFD0 U1618 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1619 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1620 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1621 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1622 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1623 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1624 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1625 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1626 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1627 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1628 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1629 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1630 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1631 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1632 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1633 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1634 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1635 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1636 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1637 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1638 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1639 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1640 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1641 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1642 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1643 ( .I(n1658), .Z(n1657) );
  BUFFD0 U1644 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1645 ( .I(n1660), .Z(n1659) );
  BUFFD0 U1646 ( .I(n1661), .Z(n1660) );
  BUFFD0 U1647 ( .I(n1662), .Z(n1661) );
  BUFFD0 U1648 ( .I(n1663), .Z(n1662) );
  BUFFD0 U1649 ( .I(n1664), .Z(n1663) );
  BUFFD0 U1650 ( .I(n1665), .Z(n1664) );
  BUFFD0 U1651 ( .I(n1666), .Z(n1665) );
  BUFFD0 U1652 ( .I(n1667), .Z(n1666) );
  BUFFD0 U1653 ( .I(n1668), .Z(n1667) );
  BUFFD0 U1654 ( .I(n1669), .Z(n1668) );
  BUFFD0 U1655 ( .I(n1670), .Z(n1669) );
  BUFFD0 U1656 ( .I(n1671), .Z(n1670) );
  BUFFD0 U1657 ( .I(n1672), .Z(n1671) );
  BUFFD0 U1658 ( .I(n1673), .Z(n1672) );
  BUFFD0 U1659 ( .I(n1674), .Z(n1673) );
  BUFFD0 U1660 ( .I(n1675), .Z(n1674) );
  BUFFD0 U1661 ( .I(n1676), .Z(n1675) );
  BUFFD0 U1662 ( .I(n1677), .Z(n1676) );
  BUFFD0 U1663 ( .I(n1678), .Z(n1677) );
  BUFFD0 U1664 ( .I(n1679), .Z(n1678) );
  BUFFD0 U1665 ( .I(n1680), .Z(n1679) );
  BUFFD0 U1666 ( .I(n1681), .Z(n1680) );
  BUFFD0 U1667 ( .I(n1682), .Z(n1681) );
  BUFFD0 U1668 ( .I(n1683), .Z(n1682) );
  BUFFD0 U1669 ( .I(n1684), .Z(n1683) );
  BUFFD0 U1670 ( .I(n1685), .Z(n1684) );
  BUFFD0 U1671 ( .I(n1686), .Z(n1685) );
  BUFFD0 U1672 ( .I(DataOr[2]), .Z(n1686) );
  BUFFD0 U1673 ( .I(n1688), .Z(n1687) );
  BUFFD0 U1674 ( .I(n1689), .Z(n1688) );
  BUFFD0 U1675 ( .I(n1690), .Z(n1689) );
  BUFFD0 U1676 ( .I(n1691), .Z(n1690) );
  BUFFD0 U1677 ( .I(n1692), .Z(n1691) );
  BUFFD0 U1678 ( .I(n1693), .Z(n1692) );
  BUFFD0 U1679 ( .I(n1694), .Z(n1693) );
  BUFFD0 U1680 ( .I(n1695), .Z(n1694) );
  BUFFD0 U1681 ( .I(n1696), .Z(n1695) );
  BUFFD0 U1682 ( .I(n1697), .Z(n1696) );
  BUFFD0 U1683 ( .I(n1698), .Z(n1697) );
  BUFFD0 U1684 ( .I(n1699), .Z(n1698) );
  BUFFD0 U1685 ( .I(n1700), .Z(n1699) );
  BUFFD0 U1686 ( .I(n1701), .Z(n1700) );
  BUFFD0 U1687 ( .I(n1702), .Z(n1701) );
  BUFFD0 U1688 ( .I(n1703), .Z(n1702) );
  BUFFD0 U1689 ( .I(n1704), .Z(n1703) );
  BUFFD0 U1690 ( .I(n1705), .Z(n1704) );
  BUFFD0 U1691 ( .I(n1706), .Z(n1705) );
  BUFFD0 U1692 ( .I(n1707), .Z(n1706) );
  BUFFD0 U1693 ( .I(n1708), .Z(n1707) );
  BUFFD0 U1694 ( .I(n1709), .Z(n1708) );
  BUFFD0 U1695 ( .I(n1710), .Z(n1709) );
  BUFFD0 U1696 ( .I(n1711), .Z(n1710) );
  BUFFD0 U1697 ( .I(n1712), .Z(n1711) );
  BUFFD0 U1698 ( .I(n1713), .Z(n1712) );
  BUFFD0 U1699 ( .I(n1714), .Z(n1713) );
  BUFFD0 U1700 ( .I(n1715), .Z(n1714) );
  BUFFD0 U1701 ( .I(n1716), .Z(n1715) );
  BUFFD0 U1702 ( .I(n1717), .Z(n1716) );
  BUFFD0 U1703 ( .I(n1718), .Z(n1717) );
  BUFFD0 U1704 ( .I(n1719), .Z(n1718) );
  BUFFD0 U1705 ( .I(n1720), .Z(n1719) );
  BUFFD0 U1706 ( .I(n1721), .Z(n1720) );
  BUFFD0 U1707 ( .I(n1722), .Z(n1721) );
  BUFFD0 U1708 ( .I(n1723), .Z(n1722) );
  BUFFD0 U1709 ( .I(n1724), .Z(n1723) );
  BUFFD0 U1710 ( .I(n1725), .Z(n1724) );
  BUFFD0 U1711 ( .I(n1726), .Z(n1725) );
  BUFFD0 U1712 ( .I(n1727), .Z(n1726) );
  BUFFD0 U1713 ( .I(n1728), .Z(n1727) );
  BUFFD0 U1714 ( .I(n1729), .Z(n1728) );
  BUFFD0 U1715 ( .I(n1730), .Z(n1729) );
  BUFFD0 U1716 ( .I(n1731), .Z(n1730) );
  BUFFD0 U1717 ( .I(n1732), .Z(n1731) );
  BUFFD0 U1718 ( .I(n1733), .Z(n1732) );
  BUFFD0 U1719 ( .I(n1734), .Z(n1733) );
  BUFFD0 U1720 ( .I(n1735), .Z(n1734) );
  BUFFD0 U1721 ( .I(n1736), .Z(n1735) );
  BUFFD0 U1722 ( .I(n1737), .Z(n1736) );
  BUFFD0 U1723 ( .I(n1738), .Z(n1737) );
  BUFFD0 U1724 ( .I(n1739), .Z(n1738) );
  BUFFD0 U1725 ( .I(n1740), .Z(n1739) );
  BUFFD0 U1726 ( .I(n1741), .Z(n1740) );
  BUFFD0 U1727 ( .I(DataOr[1]), .Z(n1741) );
  BUFFD0 U1728 ( .I(n1743), .Z(n1742) );
  BUFFD0 U1729 ( .I(n1744), .Z(n1743) );
  BUFFD0 U1730 ( .I(n1745), .Z(n1744) );
  BUFFD0 U1731 ( .I(n1746), .Z(n1745) );
  BUFFD0 U1732 ( .I(n1747), .Z(n1746) );
  BUFFD0 U1733 ( .I(n1748), .Z(n1747) );
  BUFFD0 U1734 ( .I(n1749), .Z(n1748) );
  BUFFD0 U1735 ( .I(n1750), .Z(n1749) );
  BUFFD0 U1736 ( .I(n1751), .Z(n1750) );
  BUFFD0 U1737 ( .I(n1752), .Z(n1751) );
  BUFFD0 U1738 ( .I(n1753), .Z(n1752) );
  BUFFD0 U1739 ( .I(n1754), .Z(n1753) );
  BUFFD0 U1740 ( .I(n1755), .Z(n1754) );
  BUFFD0 U1741 ( .I(n1756), .Z(n1755) );
  BUFFD0 U1742 ( .I(n1757), .Z(n1756) );
  BUFFD0 U1743 ( .I(n1758), .Z(n1757) );
  BUFFD0 U1744 ( .I(n1759), .Z(n1758) );
  BUFFD0 U1745 ( .I(n1760), .Z(n1759) );
  BUFFD0 U1746 ( .I(n1761), .Z(n1760) );
  BUFFD0 U1747 ( .I(n1762), .Z(n1761) );
  BUFFD0 U1748 ( .I(n1763), .Z(n1762) );
  BUFFD0 U1749 ( .I(n1764), .Z(n1763) );
  BUFFD0 U1750 ( .I(n1765), .Z(n1764) );
  BUFFD0 U1751 ( .I(n1766), .Z(n1765) );
  BUFFD0 U1752 ( .I(n1767), .Z(n1766) );
  BUFFD0 U1753 ( .I(n1768), .Z(n1767) );
  BUFFD0 U1754 ( .I(n1769), .Z(n1768) );
  BUFFD0 U1755 ( .I(n1770), .Z(n1769) );
  BUFFD0 U1756 ( .I(n1771), .Z(n1770) );
  BUFFD0 U1757 ( .I(n1772), .Z(n1771) );
  BUFFD0 U1758 ( .I(n1773), .Z(n1772) );
  BUFFD0 U1759 ( .I(n1774), .Z(n1773) );
  BUFFD0 U1760 ( .I(n1775), .Z(n1774) );
  BUFFD0 U1761 ( .I(n1776), .Z(n1775) );
  BUFFD0 U1762 ( .I(n1777), .Z(n1776) );
  BUFFD0 U1763 ( .I(n1778), .Z(n1777) );
  BUFFD0 U1764 ( .I(n1779), .Z(n1778) );
  BUFFD0 U1765 ( .I(n1780), .Z(n1779) );
  BUFFD0 U1766 ( .I(n1781), .Z(n1780) );
  BUFFD0 U1767 ( .I(n1782), .Z(n1781) );
  BUFFD0 U1768 ( .I(n1783), .Z(n1782) );
  BUFFD0 U1769 ( .I(n1784), .Z(n1783) );
  BUFFD0 U1770 ( .I(n1785), .Z(n1784) );
  BUFFD0 U1771 ( .I(n1786), .Z(n1785) );
  BUFFD0 U1772 ( .I(n1787), .Z(n1786) );
  BUFFD0 U1773 ( .I(n1788), .Z(n1787) );
  BUFFD0 U1774 ( .I(n1789), .Z(n1788) );
  BUFFD0 U1775 ( .I(n1790), .Z(n1789) );
  BUFFD0 U1776 ( .I(n1791), .Z(n1790) );
  BUFFD0 U1777 ( .I(n1792), .Z(n1791) );
  BUFFD0 U1778 ( .I(n1793), .Z(n1792) );
  BUFFD0 U1779 ( .I(n1794), .Z(n1793) );
  BUFFD0 U1780 ( .I(n1795), .Z(n1794) );
  BUFFD0 U1781 ( .I(n1796), .Z(n1795) );
  BUFFD0 U1782 ( .I(DataOr[0]), .Z(n1796) );
  BUFFD0 U1783 ( .I(n1801), .Z(n1797) );
  BUFFD0 U1784 ( .I(n103), .Z(n1798) );
  BUFFD0 U1785 ( .I(n1798), .Z(n1799) );
  BUFFD0 U1786 ( .I(n1799), .Z(n1800) );
  BUFFD0 U1787 ( .I(n1802), .Z(n1801) );
  BUFFD0 U1788 ( .I(n1803), .Z(n1802) );
  BUFFD0 U1789 ( .I(n1804), .Z(n1803) );
  BUFFD0 U1790 ( .I(n1805), .Z(n1804) );
  BUFFD0 U1791 ( .I(n1806), .Z(n1805) );
  BUFFD0 U1792 ( .I(n1807), .Z(n1806) );
  BUFFD0 U1793 ( .I(n1808), .Z(n1807) );
  BUFFD0 U1794 ( .I(n1809), .Z(n1808) );
  BUFFD0 U1795 ( .I(n1810), .Z(n1809) );
  BUFFD0 U1796 ( .I(n1811), .Z(n1810) );
  BUFFD0 U1797 ( .I(n1812), .Z(n1811) );
  BUFFD0 U1798 ( .I(n1813), .Z(n1812) );
  BUFFD0 U1799 ( .I(n1814), .Z(n1813) );
  BUFFD0 U1800 ( .I(n1815), .Z(n1814) );
  BUFFD0 U1801 ( .I(n1816), .Z(n1815) );
  BUFFD0 U1802 ( .I(n1817), .Z(n1816) );
  BUFFD0 U1803 ( .I(n1818), .Z(n1817) );
  BUFFD0 U1804 ( .I(n1819), .Z(n1818) );
  BUFFD0 U1805 ( .I(n1820), .Z(n1819) );
  BUFFD0 U1806 ( .I(n1821), .Z(n1820) );
  BUFFD0 U1807 ( .I(n1822), .Z(n1821) );
  BUFFD0 U1808 ( .I(n1823), .Z(n1822) );
  BUFFD0 U1809 ( .I(n1824), .Z(n1823) );
  BUFFD0 U1810 ( .I(n1825), .Z(n1824) );
  BUFFD0 U1811 ( .I(n1826), .Z(n1825) );
  BUFFD0 U1812 ( .I(n1827), .Z(n1826) );
  BUFFD0 U1813 ( .I(n1828), .Z(n1827) );
  BUFFD0 U1814 ( .I(n1829), .Z(n1828) );
  BUFFD0 U1815 ( .I(n1830), .Z(n1829) );
  BUFFD0 U1816 ( .I(n1831), .Z(n1830) );
  BUFFD0 U1817 ( .I(n1832), .Z(n1831) );
  BUFFD0 U1818 ( .I(n1833), .Z(n1832) );
  BUFFD0 U1819 ( .I(n1834), .Z(n1833) );
  BUFFD0 U1820 ( .I(n1835), .Z(n1834) );
  BUFFD0 U1821 ( .I(n1836), .Z(n1835) );
  BUFFD0 U1822 ( .I(n1837), .Z(n1836) );
  BUFFD0 U1823 ( .I(n1838), .Z(n1837) );
  BUFFD0 U1824 ( .I(n1839), .Z(n1838) );
  BUFFD0 U1825 ( .I(n1840), .Z(n1839) );
  BUFFD0 U1826 ( .I(n1841), .Z(n1840) );
  BUFFD0 U1827 ( .I(n1842), .Z(n1841) );
  BUFFD0 U1828 ( .I(n1843), .Z(n1842) );
  BUFFD0 U1829 ( .I(n1844), .Z(n1843) );
  BUFFD0 U1830 ( .I(n1845), .Z(n1844) );
  BUFFD0 U1831 ( .I(n1846), .Z(n1845) );
  BUFFD0 U1832 ( .I(n1847), .Z(n1846) );
  BUFFD0 U1833 ( .I(n1848), .Z(n1847) );
  BUFFD0 U1834 ( .I(n1849), .Z(n1848) );
  BUFFD0 U1835 ( .I(n1850), .Z(n1849) );
  BUFFD0 U1836 ( .I(n1851), .Z(n1850) );
  BUFFD0 U1837 ( .I(n1852), .Z(n1851) );
  BUFFD0 U1838 ( .I(n1853), .Z(n1852) );
  BUFFD0 U1839 ( .I(n1854), .Z(n1853) );
  BUFFD0 U1840 ( .I(n1855), .Z(n1854) );
  BUFFD0 U1841 ( .I(n1857), .Z(n1855) );
  BUFFD0 U1842 ( .I(n1859), .Z(n1856) );
  BUFFD0 U1843 ( .I(n1858), .Z(n1857) );
  BUFFD0 U1844 ( .I(n1800), .Z(n1858) );
  BUFFD0 U1845 ( .I(Dreadyr), .Z(n1859) );
  OR2D0 U1846 ( .A1(n4044), .A2(n1856), .Z(n103) );
  BUFFD0 U1847 ( .I(n1863), .Z(n1860) );
  BUFFD0 U1848 ( .I(n1861), .Z(n1862) );
  BUFFD0 U1849 ( .I(n1864), .Z(n1863) );
  BUFFD0 U1850 ( .I(n1865), .Z(n1864) );
  BUFFD0 U1851 ( .I(n1866), .Z(n1865) );
  BUFFD0 U1852 ( .I(n1867), .Z(n1866) );
  BUFFD0 U1853 ( .I(n1868), .Z(n1867) );
  BUFFD0 U1854 ( .I(n1869), .Z(n1868) );
  BUFFD0 U1855 ( .I(n1870), .Z(n1869) );
  BUFFD0 U1856 ( .I(n1871), .Z(n1870) );
  BUFFD0 U1857 ( .I(n1872), .Z(n1871) );
  BUFFD0 U1858 ( .I(n1873), .Z(n1872) );
  BUFFD0 U1859 ( .I(n1874), .Z(n1873) );
  BUFFD0 U1860 ( .I(n1875), .Z(n1874) );
  BUFFD0 U1861 ( .I(n1876), .Z(n1875) );
  BUFFD0 U1862 ( .I(n1877), .Z(n1876) );
  BUFFD0 U1863 ( .I(n1878), .Z(n1877) );
  BUFFD0 U1864 ( .I(n1879), .Z(n1878) );
  BUFFD0 U1865 ( .I(n1880), .Z(n1879) );
  BUFFD0 U1866 ( .I(n1881), .Z(n1880) );
  BUFFD0 U1867 ( .I(n1882), .Z(n1881) );
  BUFFD0 U1868 ( .I(n1883), .Z(n1882) );
  BUFFD0 U1869 ( .I(n1884), .Z(n1883) );
  BUFFD0 U1870 ( .I(n1885), .Z(n1884) );
  BUFFD0 U1871 ( .I(n1886), .Z(n1885) );
  BUFFD0 U1872 ( .I(n1887), .Z(n1886) );
  BUFFD0 U1873 ( .I(n1888), .Z(n1887) );
  BUFFD0 U1874 ( .I(n1889), .Z(n1888) );
  BUFFD0 U1875 ( .I(n1890), .Z(n1889) );
  BUFFD0 U1876 ( .I(n1891), .Z(n1890) );
  BUFFD0 U1877 ( .I(n1892), .Z(n1891) );
  BUFFD0 U1878 ( .I(n1893), .Z(n1892) );
  BUFFD0 U1879 ( .I(n1894), .Z(n1893) );
  BUFFD0 U1880 ( .I(n1895), .Z(n1894) );
  BUFFD0 U1881 ( .I(n1896), .Z(n1895) );
  BUFFD0 U1882 ( .I(n1897), .Z(n1896) );
  BUFFD0 U1883 ( .I(n1898), .Z(n1897) );
  BUFFD0 U1884 ( .I(n1899), .Z(n1898) );
  BUFFD0 U1885 ( .I(n1900), .Z(n1899) );
  BUFFD0 U1886 ( .I(n1901), .Z(n1900) );
  BUFFD0 U1887 ( .I(n1902), .Z(n1901) );
  BUFFD0 U1888 ( .I(n1903), .Z(n1902) );
  BUFFD0 U1889 ( .I(n1904), .Z(n1903) );
  BUFFD0 U1890 ( .I(n1905), .Z(n1904) );
  BUFFD0 U1891 ( .I(n1906), .Z(n1905) );
  BUFFD0 U1892 ( .I(n1907), .Z(n1906) );
  BUFFD0 U1893 ( .I(n1908), .Z(n1907) );
  BUFFD0 U1894 ( .I(n1909), .Z(n1908) );
  BUFFD0 U1895 ( .I(n1910), .Z(n1909) );
  BUFFD0 U1896 ( .I(n1911), .Z(n1910) );
  BUFFD0 U1897 ( .I(n1912), .Z(n1911) );
  BUFFD0 U1898 ( .I(n1913), .Z(n1912) );
  BUFFD0 U1899 ( .I(n1914), .Z(n1913) );
  BUFFD0 U1900 ( .I(n1915), .Z(n1914) );
  BUFFD0 U1901 ( .I(n1916), .Z(n1915) );
  BUFFD0 U1902 ( .I(n1917), .Z(n1916) );
  BUFFD0 U1903 ( .I(n1918), .Z(n1917) );
  BUFFD0 U1904 ( .I(n1919), .Z(n1918) );
  BUFFD0 U1905 ( .I(n1920), .Z(n1919) );
  BUFFD0 U1906 ( .I(n1921), .Z(n1920) );
  BUFFD0 U1907 ( .I(n1922), .Z(n1921) );
  BUFFD0 U1908 ( .I(n1923), .Z(n1922) );
  BUFFD0 U1909 ( .I(n1924), .Z(n1923) );
  BUFFD0 U1910 ( .I(n1925), .Z(n1924) );
  BUFFD0 U1911 ( .I(n1862), .Z(n1925) );
  BUFFD0 U1912 ( .I(n1929), .Z(n1926) );
  BUFFD0 U1913 ( .I(N51), .Z(n1927) );
  BUFFD0 U1914 ( .I(n1927), .Z(n1928) );
  BUFFD0 U1915 ( .I(n1930), .Z(n1929) );
  BUFFD0 U1916 ( .I(n1931), .Z(n1930) );
  BUFFD0 U1917 ( .I(n1932), .Z(n1931) );
  BUFFD0 U1918 ( .I(n1933), .Z(n1932) );
  BUFFD0 U1919 ( .I(n1934), .Z(n1933) );
  BUFFD0 U1920 ( .I(n1935), .Z(n1934) );
  BUFFD0 U1921 ( .I(n1936), .Z(n1935) );
  BUFFD0 U1922 ( .I(n1937), .Z(n1936) );
  BUFFD0 U1923 ( .I(n1938), .Z(n1937) );
  BUFFD0 U1924 ( .I(n1939), .Z(n1938) );
  BUFFD0 U1925 ( .I(n1940), .Z(n1939) );
  BUFFD0 U1926 ( .I(n1941), .Z(n1940) );
  BUFFD0 U1927 ( .I(n1942), .Z(n1941) );
  BUFFD0 U1928 ( .I(n1943), .Z(n1942) );
  BUFFD0 U1929 ( .I(n1944), .Z(n1943) );
  BUFFD0 U1930 ( .I(n1945), .Z(n1944) );
  BUFFD0 U1931 ( .I(n1946), .Z(n1945) );
  BUFFD0 U1932 ( .I(n1947), .Z(n1946) );
  BUFFD0 U1933 ( .I(n1948), .Z(n1947) );
  BUFFD0 U1934 ( .I(n1949), .Z(n1948) );
  BUFFD0 U1935 ( .I(n1950), .Z(n1949) );
  BUFFD0 U1936 ( .I(n1951), .Z(n1950) );
  BUFFD0 U1937 ( .I(n1952), .Z(n1951) );
  BUFFD0 U1938 ( .I(n1953), .Z(n1952) );
  BUFFD0 U1939 ( .I(n1954), .Z(n1953) );
  BUFFD0 U1940 ( .I(n1955), .Z(n1954) );
  BUFFD0 U1941 ( .I(n1956), .Z(n1955) );
  BUFFD0 U1942 ( .I(n1957), .Z(n1956) );
  BUFFD0 U1943 ( .I(n1958), .Z(n1957) );
  BUFFD0 U1944 ( .I(n1959), .Z(n1958) );
  BUFFD0 U1945 ( .I(n1960), .Z(n1959) );
  BUFFD0 U1946 ( .I(n1961), .Z(n1960) );
  BUFFD0 U1947 ( .I(n1962), .Z(n1961) );
  BUFFD0 U1948 ( .I(n1963), .Z(n1962) );
  BUFFD0 U1949 ( .I(n1964), .Z(n1963) );
  BUFFD0 U1950 ( .I(n1965), .Z(n1964) );
  BUFFD0 U1951 ( .I(n1966), .Z(n1965) );
  BUFFD0 U1952 ( .I(n1967), .Z(n1966) );
  BUFFD0 U1953 ( .I(n1968), .Z(n1967) );
  BUFFD0 U1954 ( .I(n1969), .Z(n1968) );
  BUFFD0 U1955 ( .I(n1970), .Z(n1969) );
  BUFFD0 U1956 ( .I(n1971), .Z(n1970) );
  BUFFD0 U1957 ( .I(n1972), .Z(n1971) );
  BUFFD0 U1958 ( .I(n1973), .Z(n1972) );
  BUFFD0 U1959 ( .I(n1974), .Z(n1973) );
  BUFFD0 U1960 ( .I(n1975), .Z(n1974) );
  BUFFD0 U1961 ( .I(n1976), .Z(n1975) );
  BUFFD0 U1962 ( .I(n1977), .Z(n1976) );
  BUFFD0 U1963 ( .I(n1978), .Z(n1977) );
  BUFFD0 U1964 ( .I(n1979), .Z(n1978) );
  BUFFD0 U1965 ( .I(n1980), .Z(n1979) );
  BUFFD0 U1966 ( .I(n1981), .Z(n1980) );
  BUFFD0 U1967 ( .I(n1982), .Z(n1981) );
  BUFFD0 U1968 ( .I(n1983), .Z(n1982) );
  BUFFD0 U1969 ( .I(n1984), .Z(n1983) );
  BUFFD0 U1970 ( .I(n1985), .Z(n1984) );
  BUFFD0 U1971 ( .I(n1986), .Z(n1985) );
  BUFFD0 U1972 ( .I(n1987), .Z(n1986) );
  BUFFD0 U1973 ( .I(n1988), .Z(n1987) );
  BUFFD0 U1974 ( .I(n1989), .Z(n1988) );
  BUFFD0 U1975 ( .I(n1990), .Z(n1989) );
  BUFFD0 U1976 ( .I(n1991), .Z(n1990) );
  BUFFD0 U1977 ( .I(n1928), .Z(n1991) );
  CKBD0 U1978 ( .CLK(N52), .C(n1993) );
  BUFFD0 U1979 ( .I(n1995), .Z(n1992) );
  BUFFD0 U1980 ( .I(n1993), .Z(n1994) );
  BUFFD0 U1981 ( .I(n1996), .Z(n1995) );
  BUFFD0 U1982 ( .I(n1997), .Z(n1996) );
  BUFFD0 U1983 ( .I(n1998), .Z(n1997) );
  BUFFD0 U1984 ( .I(n1999), .Z(n1998) );
  BUFFD0 U1985 ( .I(n2000), .Z(n1999) );
  BUFFD0 U1986 ( .I(n2001), .Z(n2000) );
  BUFFD0 U1987 ( .I(n2002), .Z(n2001) );
  BUFFD0 U1988 ( .I(n2003), .Z(n2002) );
  BUFFD0 U1989 ( .I(n2004), .Z(n2003) );
  BUFFD0 U1990 ( .I(n2005), .Z(n2004) );
  BUFFD0 U1991 ( .I(n2006), .Z(n2005) );
  BUFFD0 U1992 ( .I(n2007), .Z(n2006) );
  BUFFD0 U1993 ( .I(n2008), .Z(n2007) );
  BUFFD0 U1994 ( .I(n2009), .Z(n2008) );
  BUFFD0 U1995 ( .I(n2010), .Z(n2009) );
  BUFFD0 U1996 ( .I(n2011), .Z(n2010) );
  BUFFD0 U1997 ( .I(n2012), .Z(n2011) );
  BUFFD0 U1998 ( .I(n2013), .Z(n2012) );
  BUFFD0 U1999 ( .I(n2014), .Z(n2013) );
  BUFFD0 U2000 ( .I(n2015), .Z(n2014) );
  BUFFD0 U2001 ( .I(n2016), .Z(n2015) );
  BUFFD0 U2002 ( .I(n2017), .Z(n2016) );
  BUFFD0 U2003 ( .I(n2018), .Z(n2017) );
  BUFFD0 U2004 ( .I(n2019), .Z(n2018) );
  BUFFD0 U2005 ( .I(n2020), .Z(n2019) );
  BUFFD0 U2006 ( .I(n2021), .Z(n2020) );
  BUFFD0 U2007 ( .I(n2022), .Z(n2021) );
  BUFFD0 U2008 ( .I(n2023), .Z(n2022) );
  BUFFD0 U2009 ( .I(n2024), .Z(n2023) );
  BUFFD0 U2010 ( .I(n2025), .Z(n2024) );
  BUFFD0 U2011 ( .I(n2026), .Z(n2025) );
  BUFFD0 U2012 ( .I(n2027), .Z(n2026) );
  BUFFD0 U2013 ( .I(n2028), .Z(n2027) );
  BUFFD0 U2014 ( .I(n2029), .Z(n2028) );
  BUFFD0 U2015 ( .I(n2030), .Z(n2029) );
  BUFFD0 U2016 ( .I(n2031), .Z(n2030) );
  BUFFD0 U2017 ( .I(n2032), .Z(n2031) );
  BUFFD0 U2018 ( .I(n2033), .Z(n2032) );
  BUFFD0 U2019 ( .I(n2034), .Z(n2033) );
  BUFFD0 U2020 ( .I(n2035), .Z(n2034) );
  BUFFD0 U2021 ( .I(n2036), .Z(n2035) );
  BUFFD0 U2022 ( .I(n2037), .Z(n2036) );
  BUFFD0 U2023 ( .I(n2038), .Z(n2037) );
  BUFFD0 U2024 ( .I(n2039), .Z(n2038) );
  BUFFD0 U2025 ( .I(n2040), .Z(n2039) );
  BUFFD0 U2026 ( .I(n2041), .Z(n2040) );
  BUFFD0 U2027 ( .I(n2042), .Z(n2041) );
  BUFFD0 U2028 ( .I(n2043), .Z(n2042) );
  BUFFD0 U2029 ( .I(n2044), .Z(n2043) );
  BUFFD0 U2030 ( .I(n2045), .Z(n2044) );
  BUFFD0 U2031 ( .I(n2046), .Z(n2045) );
  BUFFD0 U2032 ( .I(n2047), .Z(n2046) );
  BUFFD0 U2033 ( .I(n2048), .Z(n2047) );
  BUFFD0 U2034 ( .I(n2049), .Z(n2048) );
  BUFFD0 U2035 ( .I(n2050), .Z(n2049) );
  BUFFD0 U2036 ( .I(n2051), .Z(n2050) );
  BUFFD0 U2037 ( .I(n2052), .Z(n2051) );
  BUFFD0 U2038 ( .I(n2053), .Z(n2052) );
  BUFFD0 U2039 ( .I(n2054), .Z(n2053) );
  BUFFD0 U2040 ( .I(n2055), .Z(n2054) );
  BUFFD0 U2041 ( .I(n2056), .Z(n2055) );
  BUFFD0 U2042 ( .I(n2057), .Z(n2056) );
  BUFFD0 U2043 ( .I(n1994), .Z(n2057) );
  CKBD0 U2044 ( .CLK(N53), .C(n2059) );
  BUFFD0 U2045 ( .I(n2061), .Z(n2058) );
  BUFFD0 U2046 ( .I(n2059), .Z(n2060) );
  BUFFD0 U2047 ( .I(n2062), .Z(n2061) );
  BUFFD0 U2048 ( .I(n2063), .Z(n2062) );
  BUFFD0 U2049 ( .I(n2064), .Z(n2063) );
  BUFFD0 U2050 ( .I(n2065), .Z(n2064) );
  BUFFD0 U2051 ( .I(n2066), .Z(n2065) );
  BUFFD0 U2052 ( .I(n2067), .Z(n2066) );
  BUFFD0 U2053 ( .I(n2068), .Z(n2067) );
  BUFFD0 U2054 ( .I(n2069), .Z(n2068) );
  BUFFD0 U2055 ( .I(n2070), .Z(n2069) );
  BUFFD0 U2056 ( .I(n2071), .Z(n2070) );
  BUFFD0 U2057 ( .I(n2072), .Z(n2071) );
  BUFFD0 U2058 ( .I(n2073), .Z(n2072) );
  BUFFD0 U2059 ( .I(n2074), .Z(n2073) );
  BUFFD0 U2060 ( .I(n2075), .Z(n2074) );
  BUFFD0 U2061 ( .I(n2076), .Z(n2075) );
  BUFFD0 U2062 ( .I(n2077), .Z(n2076) );
  BUFFD0 U2063 ( .I(n2078), .Z(n2077) );
  BUFFD0 U2064 ( .I(n2079), .Z(n2078) );
  BUFFD0 U2065 ( .I(n2080), .Z(n2079) );
  BUFFD0 U2066 ( .I(n2081), .Z(n2080) );
  BUFFD0 U2067 ( .I(n2082), .Z(n2081) );
  BUFFD0 U2068 ( .I(n2083), .Z(n2082) );
  BUFFD0 U2069 ( .I(n2084), .Z(n2083) );
  BUFFD0 U2070 ( .I(n2085), .Z(n2084) );
  BUFFD0 U2071 ( .I(n2086), .Z(n2085) );
  BUFFD0 U2072 ( .I(n2087), .Z(n2086) );
  BUFFD0 U2073 ( .I(n2088), .Z(n2087) );
  BUFFD0 U2074 ( .I(n2089), .Z(n2088) );
  BUFFD0 U2075 ( .I(n2090), .Z(n2089) );
  BUFFD0 U2076 ( .I(n2091), .Z(n2090) );
  BUFFD0 U2077 ( .I(n2092), .Z(n2091) );
  BUFFD0 U2078 ( .I(n2093), .Z(n2092) );
  BUFFD0 U2079 ( .I(n2094), .Z(n2093) );
  BUFFD0 U2080 ( .I(n2095), .Z(n2094) );
  BUFFD0 U2081 ( .I(n2096), .Z(n2095) );
  BUFFD0 U2082 ( .I(n2097), .Z(n2096) );
  BUFFD0 U2083 ( .I(n2098), .Z(n2097) );
  BUFFD0 U2084 ( .I(n2099), .Z(n2098) );
  BUFFD0 U2085 ( .I(n2100), .Z(n2099) );
  BUFFD0 U2086 ( .I(n2101), .Z(n2100) );
  BUFFD0 U2087 ( .I(n2102), .Z(n2101) );
  BUFFD0 U2088 ( .I(n2103), .Z(n2102) );
  BUFFD0 U2089 ( .I(n2104), .Z(n2103) );
  BUFFD0 U2090 ( .I(n2105), .Z(n2104) );
  BUFFD0 U2091 ( .I(n2106), .Z(n2105) );
  BUFFD0 U2092 ( .I(n2107), .Z(n2106) );
  BUFFD0 U2093 ( .I(n2108), .Z(n2107) );
  BUFFD0 U2094 ( .I(n2109), .Z(n2108) );
  BUFFD0 U2095 ( .I(n2110), .Z(n2109) );
  BUFFD0 U2096 ( .I(n2111), .Z(n2110) );
  BUFFD0 U2097 ( .I(n2112), .Z(n2111) );
  BUFFD0 U2098 ( .I(n2113), .Z(n2112) );
  BUFFD0 U2099 ( .I(n2114), .Z(n2113) );
  BUFFD0 U2100 ( .I(n2115), .Z(n2114) );
  BUFFD0 U2101 ( .I(n2116), .Z(n2115) );
  BUFFD0 U2102 ( .I(n2117), .Z(n2116) );
  BUFFD0 U2103 ( .I(n2118), .Z(n2117) );
  BUFFD0 U2104 ( .I(n2119), .Z(n2118) );
  BUFFD0 U2105 ( .I(n2120), .Z(n2119) );
  BUFFD0 U2106 ( .I(n2121), .Z(n2120) );
  BUFFD0 U2107 ( .I(n2122), .Z(n2121) );
  BUFFD0 U2108 ( .I(n2123), .Z(n2122) );
  BUFFD0 U2109 ( .I(n2060), .Z(n2123) );
  BUFFD0 U2110 ( .I(n2127), .Z(n2124) );
  BUFFD0 U2111 ( .I(n2125), .Z(n2126) );
  BUFFD0 U2112 ( .I(n2128), .Z(n2127) );
  BUFFD0 U2113 ( .I(n2129), .Z(n2128) );
  BUFFD0 U2114 ( .I(n2130), .Z(n2129) );
  BUFFD0 U2115 ( .I(n2131), .Z(n2130) );
  BUFFD0 U2116 ( .I(n2132), .Z(n2131) );
  BUFFD0 U2117 ( .I(n2133), .Z(n2132) );
  BUFFD0 U2118 ( .I(n2134), .Z(n2133) );
  BUFFD0 U2119 ( .I(n2135), .Z(n2134) );
  BUFFD0 U2120 ( .I(n2136), .Z(n2135) );
  BUFFD0 U2121 ( .I(n2137), .Z(n2136) );
  BUFFD0 U2122 ( .I(n2138), .Z(n2137) );
  BUFFD0 U2123 ( .I(n2139), .Z(n2138) );
  BUFFD0 U2124 ( .I(n2140), .Z(n2139) );
  BUFFD0 U2125 ( .I(n2141), .Z(n2140) );
  BUFFD0 U2126 ( .I(n2142), .Z(n2141) );
  BUFFD0 U2127 ( .I(n2143), .Z(n2142) );
  BUFFD0 U2128 ( .I(n2144), .Z(n2143) );
  BUFFD0 U2129 ( .I(n2145), .Z(n2144) );
  BUFFD0 U2130 ( .I(n2146), .Z(n2145) );
  BUFFD0 U2131 ( .I(n2147), .Z(n2146) );
  BUFFD0 U2132 ( .I(n2148), .Z(n2147) );
  BUFFD0 U2133 ( .I(n2149), .Z(n2148) );
  BUFFD0 U2134 ( .I(n2150), .Z(n2149) );
  BUFFD0 U2135 ( .I(n2151), .Z(n2150) );
  BUFFD0 U2136 ( .I(n2152), .Z(n2151) );
  BUFFD0 U2137 ( .I(n2153), .Z(n2152) );
  BUFFD0 U2138 ( .I(n2154), .Z(n2153) );
  BUFFD0 U2139 ( .I(n2155), .Z(n2154) );
  BUFFD0 U2140 ( .I(n2156), .Z(n2155) );
  BUFFD0 U2141 ( .I(n2157), .Z(n2156) );
  BUFFD0 U2142 ( .I(n2158), .Z(n2157) );
  BUFFD0 U2143 ( .I(n2159), .Z(n2158) );
  BUFFD0 U2144 ( .I(n2160), .Z(n2159) );
  BUFFD0 U2145 ( .I(n2161), .Z(n2160) );
  BUFFD0 U2146 ( .I(n2162), .Z(n2161) );
  BUFFD0 U2147 ( .I(n2163), .Z(n2162) );
  BUFFD0 U2148 ( .I(n2164), .Z(n2163) );
  BUFFD0 U2149 ( .I(n2165), .Z(n2164) );
  BUFFD0 U2150 ( .I(n2166), .Z(n2165) );
  BUFFD0 U2151 ( .I(n2167), .Z(n2166) );
  BUFFD0 U2152 ( .I(n2168), .Z(n2167) );
  BUFFD0 U2153 ( .I(n2169), .Z(n2168) );
  BUFFD0 U2154 ( .I(n2170), .Z(n2169) );
  BUFFD0 U2155 ( .I(n2171), .Z(n2170) );
  BUFFD0 U2156 ( .I(n2172), .Z(n2171) );
  BUFFD0 U2157 ( .I(n2173), .Z(n2172) );
  BUFFD0 U2158 ( .I(n2174), .Z(n2173) );
  BUFFD0 U2159 ( .I(n2175), .Z(n2174) );
  BUFFD0 U2160 ( .I(n2176), .Z(n2175) );
  BUFFD0 U2161 ( .I(n2177), .Z(n2176) );
  BUFFD0 U2162 ( .I(n2178), .Z(n2177) );
  BUFFD0 U2163 ( .I(n2179), .Z(n2178) );
  BUFFD0 U2164 ( .I(n2180), .Z(n2179) );
  BUFFD0 U2165 ( .I(n2181), .Z(n2180) );
  BUFFD0 U2166 ( .I(n2182), .Z(n2181) );
  BUFFD0 U2167 ( .I(n2183), .Z(n2182) );
  BUFFD0 U2168 ( .I(n2184), .Z(n2183) );
  BUFFD0 U2169 ( .I(n2185), .Z(n2184) );
  BUFFD0 U2170 ( .I(n2186), .Z(n2185) );
  BUFFD0 U2171 ( .I(n2187), .Z(n2186) );
  BUFFD0 U2172 ( .I(n2188), .Z(n2187) );
  BUFFD0 U2173 ( .I(n2189), .Z(n2188) );
  BUFFD0 U2174 ( .I(n2126), .Z(n2189) );
  BUFFD0 U2175 ( .I(n2193), .Z(n2190) );
  BUFFD0 U2176 ( .I(N55), .Z(n2191) );
  BUFFD0 U2177 ( .I(n2191), .Z(n2192) );
  BUFFD0 U2178 ( .I(n2194), .Z(n2193) );
  BUFFD0 U2179 ( .I(n2195), .Z(n2194) );
  BUFFD0 U2180 ( .I(n2196), .Z(n2195) );
  BUFFD0 U2181 ( .I(n2197), .Z(n2196) );
  BUFFD0 U2182 ( .I(n2198), .Z(n2197) );
  BUFFD0 U2183 ( .I(n2199), .Z(n2198) );
  BUFFD0 U2184 ( .I(n2200), .Z(n2199) );
  BUFFD0 U2185 ( .I(n2201), .Z(n2200) );
  BUFFD0 U2186 ( .I(n2202), .Z(n2201) );
  BUFFD0 U2187 ( .I(n2203), .Z(n2202) );
  BUFFD0 U2188 ( .I(n2204), .Z(n2203) );
  BUFFD0 U2189 ( .I(n2205), .Z(n2204) );
  BUFFD0 U2190 ( .I(n2206), .Z(n2205) );
  BUFFD0 U2191 ( .I(n2207), .Z(n2206) );
  BUFFD0 U2192 ( .I(n2208), .Z(n2207) );
  BUFFD0 U2193 ( .I(n2209), .Z(n2208) );
  BUFFD0 U2194 ( .I(n2210), .Z(n2209) );
  BUFFD0 U2195 ( .I(n2211), .Z(n2210) );
  BUFFD0 U2196 ( .I(n2212), .Z(n2211) );
  BUFFD0 U2197 ( .I(n2213), .Z(n2212) );
  BUFFD0 U2198 ( .I(n2214), .Z(n2213) );
  BUFFD0 U2199 ( .I(n2215), .Z(n2214) );
  BUFFD0 U2200 ( .I(n2216), .Z(n2215) );
  BUFFD0 U2201 ( .I(n2217), .Z(n2216) );
  BUFFD0 U2202 ( .I(n2218), .Z(n2217) );
  BUFFD0 U2203 ( .I(n2219), .Z(n2218) );
  BUFFD0 U2204 ( .I(n2220), .Z(n2219) );
  BUFFD0 U2205 ( .I(n2221), .Z(n2220) );
  BUFFD0 U2206 ( .I(n2222), .Z(n2221) );
  BUFFD0 U2207 ( .I(n2223), .Z(n2222) );
  BUFFD0 U2208 ( .I(n2224), .Z(n2223) );
  BUFFD0 U2209 ( .I(n2225), .Z(n2224) );
  BUFFD0 U2210 ( .I(n2226), .Z(n2225) );
  BUFFD0 U2211 ( .I(n2227), .Z(n2226) );
  BUFFD0 U2212 ( .I(n2228), .Z(n2227) );
  BUFFD0 U2213 ( .I(n2229), .Z(n2228) );
  BUFFD0 U2214 ( .I(n2230), .Z(n2229) );
  BUFFD0 U2215 ( .I(n2231), .Z(n2230) );
  BUFFD0 U2216 ( .I(n2232), .Z(n2231) );
  BUFFD0 U2217 ( .I(n2233), .Z(n2232) );
  BUFFD0 U2218 ( .I(n2234), .Z(n2233) );
  BUFFD0 U2219 ( .I(n2235), .Z(n2234) );
  BUFFD0 U2220 ( .I(n2236), .Z(n2235) );
  BUFFD0 U2221 ( .I(n2237), .Z(n2236) );
  BUFFD0 U2222 ( .I(n2238), .Z(n2237) );
  BUFFD0 U2223 ( .I(n2239), .Z(n2238) );
  BUFFD0 U2224 ( .I(n2240), .Z(n2239) );
  BUFFD0 U2225 ( .I(n2241), .Z(n2240) );
  BUFFD0 U2226 ( .I(n2242), .Z(n2241) );
  BUFFD0 U2227 ( .I(n2243), .Z(n2242) );
  BUFFD0 U2228 ( .I(n2244), .Z(n2243) );
  BUFFD0 U2229 ( .I(n2245), .Z(n2244) );
  BUFFD0 U2230 ( .I(n2246), .Z(n2245) );
  BUFFD0 U2231 ( .I(n2247), .Z(n2246) );
  BUFFD0 U2232 ( .I(n2248), .Z(n2247) );
  BUFFD0 U2233 ( .I(n2249), .Z(n2248) );
  BUFFD0 U2234 ( .I(n2250), .Z(n2249) );
  BUFFD0 U2235 ( .I(n2251), .Z(n2250) );
  BUFFD0 U2236 ( .I(n2252), .Z(n2251) );
  BUFFD0 U2237 ( .I(n2253), .Z(n2252) );
  BUFFD0 U2238 ( .I(n2254), .Z(n2253) );
  BUFFD0 U2239 ( .I(n2255), .Z(n2254) );
  BUFFD0 U2240 ( .I(n2192), .Z(n2255) );
  CKBD0 U2241 ( .CLK(N56), .C(n2257) );
  BUFFD0 U2242 ( .I(n2259), .Z(n2256) );
  BUFFD0 U2243 ( .I(n2257), .Z(n2258) );
  BUFFD0 U2244 ( .I(n2260), .Z(n2259) );
  BUFFD0 U2245 ( .I(n2261), .Z(n2260) );
  BUFFD0 U2246 ( .I(n2262), .Z(n2261) );
  BUFFD0 U2247 ( .I(n2263), .Z(n2262) );
  BUFFD0 U2248 ( .I(n2264), .Z(n2263) );
  BUFFD0 U2249 ( .I(n2265), .Z(n2264) );
  BUFFD0 U2250 ( .I(n2266), .Z(n2265) );
  BUFFD0 U2251 ( .I(n2267), .Z(n2266) );
  BUFFD0 U2252 ( .I(n2268), .Z(n2267) );
  BUFFD0 U2253 ( .I(n2269), .Z(n2268) );
  BUFFD0 U2254 ( .I(n2270), .Z(n2269) );
  BUFFD0 U2255 ( .I(n2271), .Z(n2270) );
  BUFFD0 U2256 ( .I(n2272), .Z(n2271) );
  BUFFD0 U2257 ( .I(n2273), .Z(n2272) );
  BUFFD0 U2258 ( .I(n2274), .Z(n2273) );
  BUFFD0 U2259 ( .I(n2275), .Z(n2274) );
  BUFFD0 U2260 ( .I(n2276), .Z(n2275) );
  BUFFD0 U2261 ( .I(n2277), .Z(n2276) );
  BUFFD0 U2262 ( .I(n2278), .Z(n2277) );
  BUFFD0 U2263 ( .I(n2279), .Z(n2278) );
  BUFFD0 U2264 ( .I(n2280), .Z(n2279) );
  BUFFD0 U2265 ( .I(n2281), .Z(n2280) );
  BUFFD0 U2266 ( .I(n2282), .Z(n2281) );
  BUFFD0 U2267 ( .I(n2283), .Z(n2282) );
  BUFFD0 U2268 ( .I(n2284), .Z(n2283) );
  BUFFD0 U2269 ( .I(n2285), .Z(n2284) );
  BUFFD0 U2270 ( .I(n2286), .Z(n2285) );
  BUFFD0 U2271 ( .I(n2287), .Z(n2286) );
  BUFFD0 U2272 ( .I(n2288), .Z(n2287) );
  BUFFD0 U2273 ( .I(n2289), .Z(n2288) );
  BUFFD0 U2274 ( .I(n2290), .Z(n2289) );
  BUFFD0 U2275 ( .I(n2291), .Z(n2290) );
  BUFFD0 U2276 ( .I(n2292), .Z(n2291) );
  BUFFD0 U2277 ( .I(n2293), .Z(n2292) );
  BUFFD0 U2278 ( .I(n2294), .Z(n2293) );
  BUFFD0 U2279 ( .I(n2295), .Z(n2294) );
  BUFFD0 U2280 ( .I(n2296), .Z(n2295) );
  BUFFD0 U2281 ( .I(n2297), .Z(n2296) );
  BUFFD0 U2282 ( .I(n2298), .Z(n2297) );
  BUFFD0 U2283 ( .I(n2299), .Z(n2298) );
  BUFFD0 U2284 ( .I(n2300), .Z(n2299) );
  BUFFD0 U2285 ( .I(n2301), .Z(n2300) );
  BUFFD0 U2286 ( .I(n2302), .Z(n2301) );
  BUFFD0 U2287 ( .I(n2303), .Z(n2302) );
  BUFFD0 U2288 ( .I(n2304), .Z(n2303) );
  BUFFD0 U2289 ( .I(n2305), .Z(n2304) );
  BUFFD0 U2290 ( .I(n2306), .Z(n2305) );
  BUFFD0 U2291 ( .I(n2307), .Z(n2306) );
  BUFFD0 U2292 ( .I(n2308), .Z(n2307) );
  BUFFD0 U2293 ( .I(n2309), .Z(n2308) );
  BUFFD0 U2294 ( .I(n2310), .Z(n2309) );
  BUFFD0 U2295 ( .I(n2311), .Z(n2310) );
  BUFFD0 U2296 ( .I(n2312), .Z(n2311) );
  BUFFD0 U2297 ( .I(n2313), .Z(n2312) );
  BUFFD0 U2298 ( .I(n2314), .Z(n2313) );
  BUFFD0 U2299 ( .I(n2315), .Z(n2314) );
  BUFFD0 U2300 ( .I(n2316), .Z(n2315) );
  BUFFD0 U2301 ( .I(n2317), .Z(n2316) );
  BUFFD0 U2302 ( .I(n2318), .Z(n2317) );
  BUFFD0 U2303 ( .I(n2319), .Z(n2318) );
  BUFFD0 U2304 ( .I(n2320), .Z(n2319) );
  BUFFD0 U2305 ( .I(n2321), .Z(n2320) );
  BUFFD0 U2306 ( .I(n2258), .Z(n2321) );
  BUFFD0 U2307 ( .I(n2325), .Z(n2322) );
  BUFFD0 U2308 ( .I(n2323), .Z(n2324) );
  BUFFD0 U2309 ( .I(n2326), .Z(n2325) );
  BUFFD0 U2310 ( .I(n2327), .Z(n2326) );
  BUFFD0 U2311 ( .I(n2328), .Z(n2327) );
  BUFFD0 U2312 ( .I(n2329), .Z(n2328) );
  BUFFD0 U2313 ( .I(n2330), .Z(n2329) );
  BUFFD0 U2314 ( .I(n2331), .Z(n2330) );
  BUFFD0 U2315 ( .I(n2332), .Z(n2331) );
  BUFFD0 U2316 ( .I(n2333), .Z(n2332) );
  BUFFD0 U2317 ( .I(n2334), .Z(n2333) );
  BUFFD0 U2318 ( .I(n2335), .Z(n2334) );
  BUFFD0 U2319 ( .I(n2336), .Z(n2335) );
  BUFFD0 U2320 ( .I(n2337), .Z(n2336) );
  BUFFD0 U2321 ( .I(n2338), .Z(n2337) );
  BUFFD0 U2322 ( .I(n2339), .Z(n2338) );
  BUFFD0 U2323 ( .I(n2340), .Z(n2339) );
  BUFFD0 U2324 ( .I(n2341), .Z(n2340) );
  BUFFD0 U2325 ( .I(n2342), .Z(n2341) );
  BUFFD0 U2326 ( .I(n2343), .Z(n2342) );
  BUFFD0 U2327 ( .I(n2344), .Z(n2343) );
  BUFFD0 U2328 ( .I(n2345), .Z(n2344) );
  BUFFD0 U2329 ( .I(n2346), .Z(n2345) );
  BUFFD0 U2330 ( .I(n2347), .Z(n2346) );
  BUFFD0 U2331 ( .I(n2348), .Z(n2347) );
  BUFFD0 U2332 ( .I(n2349), .Z(n2348) );
  BUFFD0 U2333 ( .I(n2350), .Z(n2349) );
  BUFFD0 U2334 ( .I(n2351), .Z(n2350) );
  BUFFD0 U2335 ( .I(n2352), .Z(n2351) );
  BUFFD0 U2336 ( .I(n2353), .Z(n2352) );
  BUFFD0 U2337 ( .I(n2354), .Z(n2353) );
  BUFFD0 U2338 ( .I(n2355), .Z(n2354) );
  BUFFD0 U2339 ( .I(n2356), .Z(n2355) );
  BUFFD0 U2340 ( .I(n2357), .Z(n2356) );
  BUFFD0 U2341 ( .I(n2358), .Z(n2357) );
  BUFFD0 U2342 ( .I(n2359), .Z(n2358) );
  BUFFD0 U2343 ( .I(n2360), .Z(n2359) );
  BUFFD0 U2344 ( .I(n2361), .Z(n2360) );
  BUFFD0 U2345 ( .I(n2362), .Z(n2361) );
  BUFFD0 U2346 ( .I(n2363), .Z(n2362) );
  BUFFD0 U2347 ( .I(n2364), .Z(n2363) );
  BUFFD0 U2348 ( .I(n2365), .Z(n2364) );
  BUFFD0 U2349 ( .I(n2366), .Z(n2365) );
  BUFFD0 U2350 ( .I(n2367), .Z(n2366) );
  BUFFD0 U2351 ( .I(n2368), .Z(n2367) );
  BUFFD0 U2352 ( .I(n2369), .Z(n2368) );
  BUFFD0 U2353 ( .I(n2370), .Z(n2369) );
  BUFFD0 U2354 ( .I(n2371), .Z(n2370) );
  BUFFD0 U2355 ( .I(n2372), .Z(n2371) );
  BUFFD0 U2356 ( .I(n2373), .Z(n2372) );
  BUFFD0 U2357 ( .I(n2374), .Z(n2373) );
  BUFFD0 U2358 ( .I(n2375), .Z(n2374) );
  BUFFD0 U2359 ( .I(n2376), .Z(n2375) );
  BUFFD0 U2360 ( .I(n2377), .Z(n2376) );
  BUFFD0 U2361 ( .I(n2378), .Z(n2377) );
  BUFFD0 U2362 ( .I(n2379), .Z(n2378) );
  BUFFD0 U2363 ( .I(n2380), .Z(n2379) );
  BUFFD0 U2364 ( .I(n2381), .Z(n2380) );
  BUFFD0 U2365 ( .I(n2382), .Z(n2381) );
  BUFFD0 U2366 ( .I(n2383), .Z(n2382) );
  BUFFD0 U2367 ( .I(n2384), .Z(n2383) );
  BUFFD0 U2368 ( .I(n2385), .Z(n2384) );
  BUFFD0 U2369 ( .I(n2386), .Z(n2385) );
  BUFFD0 U2370 ( .I(n2387), .Z(n2386) );
  BUFFD0 U2371 ( .I(n2324), .Z(n2387) );
  BUFFD0 U2372 ( .I(n2392), .Z(n2388) );
  BUFFD0 U2373 ( .I(n3943), .Z(n2389) );
  BUFFD0 U2374 ( .I(n2389), .Z(n2390) );
  BUFFD0 U2375 ( .I(n2390), .Z(n2391) );
  BUFFD0 U2376 ( .I(n2393), .Z(n2392) );
  BUFFD0 U2377 ( .I(n2394), .Z(n2393) );
  BUFFD0 U2378 ( .I(n2395), .Z(n2394) );
  BUFFD0 U2379 ( .I(n2396), .Z(n2395) );
  BUFFD0 U2380 ( .I(n2397), .Z(n2396) );
  BUFFD0 U2381 ( .I(n2398), .Z(n2397) );
  BUFFD0 U2382 ( .I(n2399), .Z(n2398) );
  BUFFD0 U2383 ( .I(n2400), .Z(n2399) );
  BUFFD0 U2384 ( .I(n2401), .Z(n2400) );
  BUFFD0 U2385 ( .I(n2402), .Z(n2401) );
  BUFFD0 U2386 ( .I(n2403), .Z(n2402) );
  BUFFD0 U2387 ( .I(n2404), .Z(n2403) );
  BUFFD0 U2388 ( .I(n2405), .Z(n2404) );
  BUFFD0 U2389 ( .I(n2406), .Z(n2405) );
  BUFFD0 U2390 ( .I(n2407), .Z(n2406) );
  BUFFD0 U2391 ( .I(n2408), .Z(n2407) );
  BUFFD0 U2392 ( .I(n2409), .Z(n2408) );
  BUFFD0 U2393 ( .I(n2410), .Z(n2409) );
  BUFFD0 U2394 ( .I(n2411), .Z(n2410) );
  BUFFD0 U2395 ( .I(n2412), .Z(n2411) );
  BUFFD0 U2396 ( .I(n2413), .Z(n2412) );
  BUFFD0 U2397 ( .I(n2414), .Z(n2413) );
  BUFFD0 U2398 ( .I(n2415), .Z(n2414) );
  BUFFD0 U2399 ( .I(n2416), .Z(n2415) );
  BUFFD0 U2400 ( .I(n2417), .Z(n2416) );
  BUFFD0 U2401 ( .I(n2418), .Z(n2417) );
  BUFFD0 U2402 ( .I(n2419), .Z(n2418) );
  BUFFD0 U2403 ( .I(n2420), .Z(n2419) );
  BUFFD0 U2404 ( .I(n2421), .Z(n2420) );
  BUFFD0 U2405 ( .I(n2422), .Z(n2421) );
  BUFFD0 U2406 ( .I(n2423), .Z(n2422) );
  BUFFD0 U2407 ( .I(n2424), .Z(n2423) );
  BUFFD0 U2408 ( .I(n2425), .Z(n2424) );
  BUFFD0 U2409 ( .I(n2426), .Z(n2425) );
  BUFFD0 U2410 ( .I(n2427), .Z(n2426) );
  BUFFD0 U2411 ( .I(n2428), .Z(n2427) );
  BUFFD0 U2412 ( .I(n2429), .Z(n2428) );
  BUFFD0 U2413 ( .I(n2430), .Z(n2429) );
  BUFFD0 U2414 ( .I(n2431), .Z(n2430) );
  BUFFD0 U2415 ( .I(n2432), .Z(n2431) );
  BUFFD0 U2416 ( .I(n2433), .Z(n2432) );
  BUFFD0 U2417 ( .I(n2434), .Z(n2433) );
  BUFFD0 U2418 ( .I(n2435), .Z(n2434) );
  BUFFD0 U2419 ( .I(n2436), .Z(n2435) );
  BUFFD0 U2420 ( .I(n2437), .Z(n2436) );
  BUFFD0 U2421 ( .I(n2438), .Z(n2437) );
  BUFFD0 U2422 ( .I(n2439), .Z(n2438) );
  BUFFD0 U2423 ( .I(n2440), .Z(n2439) );
  BUFFD0 U2424 ( .I(n2441), .Z(n2440) );
  BUFFD0 U2425 ( .I(n2442), .Z(n2441) );
  BUFFD0 U2426 ( .I(n2443), .Z(n2442) );
  BUFFD0 U2427 ( .I(n2444), .Z(n2443) );
  BUFFD0 U2428 ( .I(n2445), .Z(n2444) );
  BUFFD0 U2429 ( .I(n2446), .Z(n2445) );
  BUFFD0 U2430 ( .I(n2447), .Z(n2446) );
  BUFFD0 U2431 ( .I(n2448), .Z(n2447) );
  BUFFD0 U2432 ( .I(n2449), .Z(n2448) );
  BUFFD0 U2433 ( .I(n2450), .Z(n2449) );
  BUFFD0 U2434 ( .I(n2391), .Z(n2450) );
  BUFFD0 U2435 ( .I(N58), .Z(n2451) );
  BUFFD0 U2436 ( .I(n2451), .Z(n2452) );
  BUFFD0 U2437 ( .I(n2452), .Z(n2453) );
  BUFFD0 U2438 ( .I(n2458), .Z(n2454) );
  BUFFD0 U2439 ( .I(N59), .Z(n2455) );
  BUFFD0 U2440 ( .I(n2455), .Z(n2456) );
  BUFFD0 U2441 ( .I(n2456), .Z(n2457) );
  BUFFD0 U2442 ( .I(n2459), .Z(n2458) );
  BUFFD0 U2443 ( .I(n2460), .Z(n2459) );
  BUFFD0 U2444 ( .I(n2461), .Z(n2460) );
  BUFFD0 U2445 ( .I(n2462), .Z(n2461) );
  BUFFD0 U2446 ( .I(n2463), .Z(n2462) );
  BUFFD0 U2447 ( .I(n2464), .Z(n2463) );
  BUFFD0 U2448 ( .I(n2465), .Z(n2464) );
  BUFFD0 U2449 ( .I(n2466), .Z(n2465) );
  BUFFD0 U2450 ( .I(n2467), .Z(n2466) );
  BUFFD0 U2451 ( .I(n2468), .Z(n2467) );
  BUFFD0 U2452 ( .I(n2469), .Z(n2468) );
  BUFFD0 U2453 ( .I(n2470), .Z(n2469) );
  BUFFD0 U2454 ( .I(n2471), .Z(n2470) );
  BUFFD0 U2455 ( .I(n2472), .Z(n2471) );
  BUFFD0 U2456 ( .I(n2473), .Z(n2472) );
  BUFFD0 U2457 ( .I(n2474), .Z(n2473) );
  BUFFD0 U2458 ( .I(n2475), .Z(n2474) );
  BUFFD0 U2459 ( .I(n2476), .Z(n2475) );
  BUFFD0 U2460 ( .I(n2477), .Z(n2476) );
  BUFFD0 U2461 ( .I(n2478), .Z(n2477) );
  BUFFD0 U2462 ( .I(n2479), .Z(n2478) );
  BUFFD0 U2463 ( .I(n2480), .Z(n2479) );
  BUFFD0 U2464 ( .I(n2481), .Z(n2480) );
  BUFFD0 U2465 ( .I(n2482), .Z(n2481) );
  BUFFD0 U2466 ( .I(n2483), .Z(n2482) );
  BUFFD0 U2467 ( .I(n2484), .Z(n2483) );
  BUFFD0 U2468 ( .I(n2485), .Z(n2484) );
  BUFFD0 U2469 ( .I(n2486), .Z(n2485) );
  BUFFD0 U2470 ( .I(n2487), .Z(n2486) );
  BUFFD0 U2471 ( .I(n2488), .Z(n2487) );
  BUFFD0 U2472 ( .I(n2489), .Z(n2488) );
  BUFFD0 U2473 ( .I(n2490), .Z(n2489) );
  BUFFD0 U2474 ( .I(n2491), .Z(n2490) );
  BUFFD0 U2475 ( .I(n2492), .Z(n2491) );
  BUFFD0 U2476 ( .I(n2493), .Z(n2492) );
  BUFFD0 U2477 ( .I(n2494), .Z(n2493) );
  BUFFD0 U2478 ( .I(n2495), .Z(n2494) );
  BUFFD0 U2479 ( .I(n2496), .Z(n2495) );
  BUFFD0 U2480 ( .I(n2497), .Z(n2496) );
  BUFFD0 U2481 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2482 ( .I(n2499), .Z(n2498) );
  BUFFD0 U2483 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2484 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2485 ( .I(n2502), .Z(n2501) );
  BUFFD0 U2486 ( .I(n2503), .Z(n2502) );
  BUFFD0 U2487 ( .I(n2504), .Z(n2503) );
  BUFFD0 U2488 ( .I(n2505), .Z(n2504) );
  BUFFD0 U2489 ( .I(n2506), .Z(n2505) );
  BUFFD0 U2490 ( .I(n2507), .Z(n2506) );
  BUFFD0 U2491 ( .I(n2508), .Z(n2507) );
  BUFFD0 U2492 ( .I(n2509), .Z(n2508) );
  BUFFD0 U2493 ( .I(n2510), .Z(n2509) );
  BUFFD0 U2494 ( .I(n2511), .Z(n2510) );
  BUFFD0 U2495 ( .I(n2512), .Z(n2511) );
  BUFFD0 U2496 ( .I(n2513), .Z(n2512) );
  BUFFD0 U2497 ( .I(n2514), .Z(n2513) );
  BUFFD0 U2498 ( .I(n2515), .Z(n2514) );
  BUFFD0 U2499 ( .I(n3925), .Z(n2515) );
  BUFFD0 U2500 ( .I(n2457), .Z(n2516) );
  BUFFD0 U2501 ( .I(n2516), .Z(n2517) );
  BUFFD0 U2502 ( .I(n2517), .Z(n2518) );
  BUFFD0 U2503 ( .I(n2523), .Z(n2519) );
  BUFFD0 U2504 ( .I(N60), .Z(n2520) );
  BUFFD0 U2505 ( .I(n2520), .Z(n2521) );
  BUFFD0 U2506 ( .I(n2521), .Z(n2522) );
  BUFFD0 U2507 ( .I(n2524), .Z(n2523) );
  BUFFD0 U2508 ( .I(n2525), .Z(n2524) );
  BUFFD0 U2509 ( .I(n2526), .Z(n2525) );
  BUFFD0 U2510 ( .I(n2527), .Z(n2526) );
  BUFFD0 U2511 ( .I(n2528), .Z(n2527) );
  BUFFD0 U2512 ( .I(n2529), .Z(n2528) );
  BUFFD0 U2513 ( .I(n2530), .Z(n2529) );
  BUFFD0 U2514 ( .I(n2531), .Z(n2530) );
  BUFFD0 U2515 ( .I(n2532), .Z(n2531) );
  BUFFD0 U2516 ( .I(n2533), .Z(n2532) );
  BUFFD0 U2517 ( .I(n2534), .Z(n2533) );
  BUFFD0 U2518 ( .I(n2535), .Z(n2534) );
  BUFFD0 U2519 ( .I(n2536), .Z(n2535) );
  BUFFD0 U2520 ( .I(n2537), .Z(n2536) );
  BUFFD0 U2521 ( .I(n2538), .Z(n2537) );
  BUFFD0 U2522 ( .I(n2539), .Z(n2538) );
  BUFFD0 U2523 ( .I(n2540), .Z(n2539) );
  BUFFD0 U2524 ( .I(n2541), .Z(n2540) );
  BUFFD0 U2525 ( .I(n2542), .Z(n2541) );
  BUFFD0 U2526 ( .I(n2543), .Z(n2542) );
  BUFFD0 U2527 ( .I(n2544), .Z(n2543) );
  BUFFD0 U2528 ( .I(n2545), .Z(n2544) );
  BUFFD0 U2529 ( .I(n2546), .Z(n2545) );
  BUFFD0 U2530 ( .I(n2547), .Z(n2546) );
  BUFFD0 U2531 ( .I(n2548), .Z(n2547) );
  BUFFD0 U2532 ( .I(n2549), .Z(n2548) );
  BUFFD0 U2533 ( .I(n2550), .Z(n2549) );
  BUFFD0 U2534 ( .I(n2551), .Z(n2550) );
  BUFFD0 U2535 ( .I(n2552), .Z(n2551) );
  BUFFD0 U2536 ( .I(n2553), .Z(n2552) );
  BUFFD0 U2537 ( .I(n2554), .Z(n2553) );
  BUFFD0 U2538 ( .I(n2555), .Z(n2554) );
  BUFFD0 U2539 ( .I(n2556), .Z(n2555) );
  BUFFD0 U2540 ( .I(n2557), .Z(n2556) );
  BUFFD0 U2541 ( .I(n2558), .Z(n2557) );
  BUFFD0 U2542 ( .I(n2559), .Z(n2558) );
  BUFFD0 U2543 ( .I(n2560), .Z(n2559) );
  BUFFD0 U2544 ( .I(n2561), .Z(n2560) );
  BUFFD0 U2545 ( .I(n2562), .Z(n2561) );
  BUFFD0 U2546 ( .I(n2563), .Z(n2562) );
  BUFFD0 U2547 ( .I(n2564), .Z(n2563) );
  BUFFD0 U2548 ( .I(n2565), .Z(n2564) );
  BUFFD0 U2549 ( .I(n2566), .Z(n2565) );
  BUFFD0 U2550 ( .I(n2567), .Z(n2566) );
  BUFFD0 U2551 ( .I(n2568), .Z(n2567) );
  BUFFD0 U2552 ( .I(n2569), .Z(n2568) );
  BUFFD0 U2553 ( .I(n2570), .Z(n2569) );
  BUFFD0 U2554 ( .I(n2571), .Z(n2570) );
  BUFFD0 U2555 ( .I(n2572), .Z(n2571) );
  BUFFD0 U2556 ( .I(n2573), .Z(n2572) );
  BUFFD0 U2557 ( .I(n2574), .Z(n2573) );
  BUFFD0 U2558 ( .I(n2575), .Z(n2574) );
  BUFFD0 U2559 ( .I(n2576), .Z(n2575) );
  BUFFD0 U2560 ( .I(n2577), .Z(n2576) );
  BUFFD0 U2561 ( .I(n2578), .Z(n2577) );
  BUFFD0 U2562 ( .I(n2579), .Z(n2578) );
  BUFFD0 U2563 ( .I(n2580), .Z(n2579) );
  BUFFD0 U2564 ( .I(n3932), .Z(n2580) );
  BUFFD0 U2565 ( .I(n2522), .Z(n2581) );
  BUFFD0 U2566 ( .I(n2581), .Z(n2582) );
  BUFFD0 U2567 ( .I(n2582), .Z(n2583) );
  BUFFD0 U2568 ( .I(n2583), .Z(n2584) );
  BUFFD0 U2569 ( .I(n2589), .Z(n2585) );
  BUFFD0 U2570 ( .I(n3924), .Z(n2586) );
  BUFFD0 U2571 ( .I(n2586), .Z(n2587) );
  BUFFD0 U2572 ( .I(n2587), .Z(n2588) );
  BUFFD0 U2573 ( .I(n2590), .Z(n2589) );
  BUFFD0 U2574 ( .I(n2591), .Z(n2590) );
  BUFFD0 U2575 ( .I(n2592), .Z(n2591) );
  BUFFD0 U2576 ( .I(n2593), .Z(n2592) );
  BUFFD0 U2577 ( .I(n2594), .Z(n2593) );
  BUFFD0 U2578 ( .I(n2595), .Z(n2594) );
  BUFFD0 U2579 ( .I(n2596), .Z(n2595) );
  BUFFD0 U2580 ( .I(n2597), .Z(n2596) );
  BUFFD0 U2581 ( .I(n2598), .Z(n2597) );
  BUFFD0 U2582 ( .I(n2599), .Z(n2598) );
  BUFFD0 U2583 ( .I(n2600), .Z(n2599) );
  BUFFD0 U2584 ( .I(n2601), .Z(n2600) );
  BUFFD0 U2585 ( .I(n2602), .Z(n2601) );
  BUFFD0 U2586 ( .I(n2603), .Z(n2602) );
  BUFFD0 U2587 ( .I(n2604), .Z(n2603) );
  BUFFD0 U2588 ( .I(n2605), .Z(n2604) );
  BUFFD0 U2589 ( .I(n2606), .Z(n2605) );
  BUFFD0 U2590 ( .I(n2607), .Z(n2606) );
  BUFFD0 U2591 ( .I(n2608), .Z(n2607) );
  BUFFD0 U2592 ( .I(n2609), .Z(n2608) );
  BUFFD0 U2593 ( .I(n2610), .Z(n2609) );
  BUFFD0 U2594 ( .I(n2611), .Z(n2610) );
  BUFFD0 U2595 ( .I(n2612), .Z(n2611) );
  BUFFD0 U2596 ( .I(n2613), .Z(n2612) );
  BUFFD0 U2597 ( .I(n2614), .Z(n2613) );
  BUFFD0 U2598 ( .I(n2615), .Z(n2614) );
  BUFFD0 U2599 ( .I(n2616), .Z(n2615) );
  BUFFD0 U2600 ( .I(n2617), .Z(n2616) );
  BUFFD0 U2601 ( .I(n2618), .Z(n2617) );
  BUFFD0 U2602 ( .I(n2619), .Z(n2618) );
  BUFFD0 U2603 ( .I(n2620), .Z(n2619) );
  BUFFD0 U2604 ( .I(n2621), .Z(n2620) );
  BUFFD0 U2605 ( .I(n2622), .Z(n2621) );
  BUFFD0 U2606 ( .I(n2623), .Z(n2622) );
  BUFFD0 U2607 ( .I(n2624), .Z(n2623) );
  BUFFD0 U2608 ( .I(n2625), .Z(n2624) );
  BUFFD0 U2609 ( .I(n2626), .Z(n2625) );
  BUFFD0 U2610 ( .I(n2627), .Z(n2626) );
  BUFFD0 U2611 ( .I(n2628), .Z(n2627) );
  BUFFD0 U2612 ( .I(n2629), .Z(n2628) );
  BUFFD0 U2613 ( .I(n2630), .Z(n2629) );
  BUFFD0 U2614 ( .I(n2631), .Z(n2630) );
  BUFFD0 U2615 ( .I(n2632), .Z(n2631) );
  BUFFD0 U2616 ( .I(n2633), .Z(n2632) );
  BUFFD0 U2617 ( .I(n2634), .Z(n2633) );
  BUFFD0 U2618 ( .I(n2635), .Z(n2634) );
  BUFFD0 U2619 ( .I(n2636), .Z(n2635) );
  BUFFD0 U2620 ( .I(n2637), .Z(n2636) );
  BUFFD0 U2621 ( .I(n2638), .Z(n2637) );
  BUFFD0 U2622 ( .I(n2639), .Z(n2638) );
  BUFFD0 U2623 ( .I(n2640), .Z(n2639) );
  BUFFD0 U2624 ( .I(n2641), .Z(n2640) );
  BUFFD0 U2625 ( .I(n2642), .Z(n2641) );
  BUFFD0 U2626 ( .I(n2643), .Z(n2642) );
  BUFFD0 U2627 ( .I(n2644), .Z(n2643) );
  BUFFD0 U2628 ( .I(n2645), .Z(n2644) );
  BUFFD0 U2629 ( .I(n2646), .Z(n2645) );
  BUFFD0 U2630 ( .I(n2647), .Z(n2646) );
  BUFFD0 U2631 ( .I(n2588), .Z(n2647) );
  BUFFD0 U2632 ( .I(N61), .Z(n2648) );
  BUFFD0 U2633 ( .I(n2648), .Z(n2649) );
  BUFFD0 U2634 ( .I(n2649), .Z(n2650) );
  BUFFD0 U2635 ( .I(n2655), .Z(n2651) );
  BUFFD0 U2636 ( .I(n3931), .Z(n2652) );
  BUFFD0 U2637 ( .I(n2652), .Z(n2653) );
  BUFFD0 U2638 ( .I(n2653), .Z(n2654) );
  BUFFD0 U2639 ( .I(n2656), .Z(n2655) );
  BUFFD0 U2640 ( .I(n2657), .Z(n2656) );
  BUFFD0 U2641 ( .I(n2658), .Z(n2657) );
  BUFFD0 U2642 ( .I(n2659), .Z(n2658) );
  BUFFD0 U2643 ( .I(n2660), .Z(n2659) );
  BUFFD0 U2644 ( .I(n2661), .Z(n2660) );
  BUFFD0 U2645 ( .I(n2662), .Z(n2661) );
  BUFFD0 U2646 ( .I(n2663), .Z(n2662) );
  BUFFD0 U2647 ( .I(n2664), .Z(n2663) );
  BUFFD0 U2648 ( .I(n2665), .Z(n2664) );
  BUFFD0 U2649 ( .I(n2666), .Z(n2665) );
  BUFFD0 U2650 ( .I(n2667), .Z(n2666) );
  BUFFD0 U2651 ( .I(n2668), .Z(n2667) );
  BUFFD0 U2652 ( .I(n2669), .Z(n2668) );
  BUFFD0 U2653 ( .I(n2670), .Z(n2669) );
  BUFFD0 U2654 ( .I(n2671), .Z(n2670) );
  BUFFD0 U2655 ( .I(n2672), .Z(n2671) );
  BUFFD0 U2656 ( .I(n2673), .Z(n2672) );
  BUFFD0 U2657 ( .I(n2674), .Z(n2673) );
  BUFFD0 U2658 ( .I(n2675), .Z(n2674) );
  BUFFD0 U2659 ( .I(n2676), .Z(n2675) );
  BUFFD0 U2660 ( .I(n2677), .Z(n2676) );
  BUFFD0 U2661 ( .I(n2678), .Z(n2677) );
  BUFFD0 U2662 ( .I(n2679), .Z(n2678) );
  BUFFD0 U2663 ( .I(n2680), .Z(n2679) );
  BUFFD0 U2664 ( .I(n2681), .Z(n2680) );
  BUFFD0 U2665 ( .I(n2682), .Z(n2681) );
  BUFFD0 U2666 ( .I(n2683), .Z(n2682) );
  BUFFD0 U2667 ( .I(n2684), .Z(n2683) );
  BUFFD0 U2668 ( .I(n2685), .Z(n2684) );
  BUFFD0 U2669 ( .I(n2686), .Z(n2685) );
  BUFFD0 U2670 ( .I(n2687), .Z(n2686) );
  BUFFD0 U2671 ( .I(n2688), .Z(n2687) );
  BUFFD0 U2672 ( .I(n2689), .Z(n2688) );
  BUFFD0 U2673 ( .I(n2690), .Z(n2689) );
  BUFFD0 U2674 ( .I(n2691), .Z(n2690) );
  BUFFD0 U2675 ( .I(n2692), .Z(n2691) );
  BUFFD0 U2676 ( .I(n2693), .Z(n2692) );
  BUFFD0 U2677 ( .I(n2694), .Z(n2693) );
  BUFFD0 U2678 ( .I(n2695), .Z(n2694) );
  BUFFD0 U2679 ( .I(n2696), .Z(n2695) );
  BUFFD0 U2680 ( .I(n2697), .Z(n2696) );
  BUFFD0 U2681 ( .I(n2698), .Z(n2697) );
  BUFFD0 U2682 ( .I(n2699), .Z(n2698) );
  BUFFD0 U2683 ( .I(n2700), .Z(n2699) );
  BUFFD0 U2684 ( .I(n2701), .Z(n2700) );
  BUFFD0 U2685 ( .I(n2702), .Z(n2701) );
  BUFFD0 U2686 ( .I(n2703), .Z(n2702) );
  BUFFD0 U2687 ( .I(n2704), .Z(n2703) );
  BUFFD0 U2688 ( .I(n2705), .Z(n2704) );
  BUFFD0 U2689 ( .I(n2706), .Z(n2705) );
  BUFFD0 U2690 ( .I(n2707), .Z(n2706) );
  BUFFD0 U2691 ( .I(n2708), .Z(n2707) );
  BUFFD0 U2692 ( .I(n2709), .Z(n2708) );
  BUFFD0 U2693 ( .I(n2710), .Z(n2709) );
  BUFFD0 U2694 ( .I(n2711), .Z(n2710) );
  BUFFD0 U2695 ( .I(n2712), .Z(n2711) );
  BUFFD0 U2696 ( .I(n2713), .Z(n2712) );
  BUFFD0 U2697 ( .I(n2654), .Z(n2713) );
  BUFFD0 U2698 ( .I(N62), .Z(n2714) );
  BUFFD0 U2699 ( .I(n2714), .Z(n2715) );
  BUFFD0 U2700 ( .I(n2715), .Z(n2716) );
  BUFFD0 U2701 ( .I(n2721), .Z(n2717) );
  BUFFD0 U2702 ( .I(N63), .Z(n2718) );
  BUFFD0 U2703 ( .I(n2718), .Z(n2719) );
  BUFFD0 U2704 ( .I(n2719), .Z(n2720) );
  BUFFD0 U2705 ( .I(n2722), .Z(n2721) );
  BUFFD0 U2706 ( .I(n2723), .Z(n2722) );
  BUFFD0 U2707 ( .I(n2724), .Z(n2723) );
  BUFFD0 U2708 ( .I(n2725), .Z(n2724) );
  BUFFD0 U2709 ( .I(n2726), .Z(n2725) );
  BUFFD0 U2710 ( .I(n2727), .Z(n2726) );
  BUFFD0 U2711 ( .I(n2728), .Z(n2727) );
  BUFFD0 U2712 ( .I(n2729), .Z(n2728) );
  BUFFD0 U2713 ( .I(n2730), .Z(n2729) );
  BUFFD0 U2714 ( .I(n2731), .Z(n2730) );
  BUFFD0 U2715 ( .I(n2732), .Z(n2731) );
  BUFFD0 U2716 ( .I(n2733), .Z(n2732) );
  BUFFD0 U2717 ( .I(n2734), .Z(n2733) );
  BUFFD0 U2718 ( .I(n2735), .Z(n2734) );
  BUFFD0 U2719 ( .I(n2736), .Z(n2735) );
  BUFFD0 U2720 ( .I(n2737), .Z(n2736) );
  BUFFD0 U2721 ( .I(n2738), .Z(n2737) );
  BUFFD0 U2722 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2723 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2724 ( .I(n2741), .Z(n2740) );
  BUFFD0 U2725 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2726 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2727 ( .I(n2744), .Z(n2743) );
  BUFFD0 U2728 ( .I(n2745), .Z(n2744) );
  BUFFD0 U2729 ( .I(n2746), .Z(n2745) );
  BUFFD0 U2730 ( .I(n2747), .Z(n2746) );
  BUFFD0 U2731 ( .I(n2748), .Z(n2747) );
  BUFFD0 U2732 ( .I(n2749), .Z(n2748) );
  BUFFD0 U2733 ( .I(n2750), .Z(n2749) );
  BUFFD0 U2734 ( .I(n2751), .Z(n2750) );
  BUFFD0 U2735 ( .I(n2752), .Z(n2751) );
  BUFFD0 U2736 ( .I(n2753), .Z(n2752) );
  BUFFD0 U2737 ( .I(n2754), .Z(n2753) );
  BUFFD0 U2738 ( .I(n2755), .Z(n2754) );
  BUFFD0 U2739 ( .I(n2756), .Z(n2755) );
  BUFFD0 U2740 ( .I(n2757), .Z(n2756) );
  BUFFD0 U2741 ( .I(n2758), .Z(n2757) );
  BUFFD0 U2742 ( .I(n2759), .Z(n2758) );
  BUFFD0 U2743 ( .I(n2760), .Z(n2759) );
  BUFFD0 U2744 ( .I(n2761), .Z(n2760) );
  BUFFD0 U2745 ( .I(n2762), .Z(n2761) );
  BUFFD0 U2746 ( .I(n2763), .Z(n2762) );
  BUFFD0 U2747 ( .I(n2764), .Z(n2763) );
  BUFFD0 U2748 ( .I(n2765), .Z(n2764) );
  BUFFD0 U2749 ( .I(n2766), .Z(n2765) );
  BUFFD0 U2750 ( .I(n2767), .Z(n2766) );
  BUFFD0 U2751 ( .I(n2768), .Z(n2767) );
  BUFFD0 U2752 ( .I(n2769), .Z(n2768) );
  BUFFD0 U2753 ( .I(n2770), .Z(n2769) );
  BUFFD0 U2754 ( .I(n2771), .Z(n2770) );
  BUFFD0 U2755 ( .I(n2772), .Z(n2771) );
  BUFFD0 U2756 ( .I(n2773), .Z(n2772) );
  BUFFD0 U2757 ( .I(n2774), .Z(n2773) );
  BUFFD0 U2758 ( .I(n2775), .Z(n2774) );
  BUFFD0 U2759 ( .I(n2776), .Z(n2775) );
  BUFFD0 U2760 ( .I(n2777), .Z(n2776) );
  BUFFD0 U2761 ( .I(n2778), .Z(n2777) );
  BUFFD0 U2762 ( .I(n3935), .Z(n2778) );
  BUFFD0 U2763 ( .I(n2720), .Z(n2779) );
  BUFFD0 U2764 ( .I(n2779), .Z(n2780) );
  BUFFD0 U2765 ( .I(n2780), .Z(n2781) );
  BUFFD0 U2766 ( .I(n2781), .Z(n2782) );
  BUFFD0 U2767 ( .I(n2787), .Z(n2783) );
  BUFFD0 U2768 ( .I(n3933), .Z(n2784) );
  BUFFD0 U2769 ( .I(n2784), .Z(n2785) );
  BUFFD0 U2770 ( .I(n2785), .Z(n2786) );
  BUFFD0 U2771 ( .I(n2788), .Z(n2787) );
  BUFFD0 U2772 ( .I(n2789), .Z(n2788) );
  BUFFD0 U2773 ( .I(n2790), .Z(n2789) );
  BUFFD0 U2774 ( .I(n2791), .Z(n2790) );
  BUFFD0 U2775 ( .I(n2792), .Z(n2791) );
  BUFFD0 U2776 ( .I(n2793), .Z(n2792) );
  BUFFD0 U2777 ( .I(n2794), .Z(n2793) );
  BUFFD0 U2778 ( .I(n2795), .Z(n2794) );
  BUFFD0 U2779 ( .I(n2796), .Z(n2795) );
  BUFFD0 U2780 ( .I(n2797), .Z(n2796) );
  BUFFD0 U2781 ( .I(n2798), .Z(n2797) );
  BUFFD0 U2782 ( .I(n2799), .Z(n2798) );
  BUFFD0 U2783 ( .I(n2800), .Z(n2799) );
  BUFFD0 U2784 ( .I(n2801), .Z(n2800) );
  BUFFD0 U2785 ( .I(n2802), .Z(n2801) );
  BUFFD0 U2786 ( .I(n2803), .Z(n2802) );
  BUFFD0 U2787 ( .I(n2804), .Z(n2803) );
  BUFFD0 U2788 ( .I(n2805), .Z(n2804) );
  BUFFD0 U2789 ( .I(n2806), .Z(n2805) );
  BUFFD0 U2790 ( .I(n2807), .Z(n2806) );
  BUFFD0 U2791 ( .I(n2808), .Z(n2807) );
  BUFFD0 U2792 ( .I(n2809), .Z(n2808) );
  BUFFD0 U2793 ( .I(n2810), .Z(n2809) );
  BUFFD0 U2794 ( .I(n2811), .Z(n2810) );
  BUFFD0 U2795 ( .I(n2812), .Z(n2811) );
  BUFFD0 U2796 ( .I(n2813), .Z(n2812) );
  BUFFD0 U2797 ( .I(n2814), .Z(n2813) );
  BUFFD0 U2798 ( .I(n2815), .Z(n2814) );
  BUFFD0 U2799 ( .I(n2816), .Z(n2815) );
  BUFFD0 U2800 ( .I(n2817), .Z(n2816) );
  BUFFD0 U2801 ( .I(n2818), .Z(n2817) );
  BUFFD0 U2802 ( .I(n2819), .Z(n2818) );
  BUFFD0 U2803 ( .I(n2820), .Z(n2819) );
  BUFFD0 U2804 ( .I(n2821), .Z(n2820) );
  BUFFD0 U2805 ( .I(n2822), .Z(n2821) );
  BUFFD0 U2806 ( .I(n2823), .Z(n2822) );
  BUFFD0 U2807 ( .I(n2824), .Z(n2823) );
  BUFFD0 U2808 ( .I(n2825), .Z(n2824) );
  BUFFD0 U2809 ( .I(n2826), .Z(n2825) );
  BUFFD0 U2810 ( .I(n2827), .Z(n2826) );
  BUFFD0 U2811 ( .I(n2828), .Z(n2827) );
  BUFFD0 U2812 ( .I(n2829), .Z(n2828) );
  BUFFD0 U2813 ( .I(n2830), .Z(n2829) );
  BUFFD0 U2814 ( .I(n2831), .Z(n2830) );
  BUFFD0 U2815 ( .I(n2832), .Z(n2831) );
  BUFFD0 U2816 ( .I(n2833), .Z(n2832) );
  BUFFD0 U2817 ( .I(n2834), .Z(n2833) );
  BUFFD0 U2818 ( .I(n2835), .Z(n2834) );
  BUFFD0 U2819 ( .I(n2836), .Z(n2835) );
  BUFFD0 U2820 ( .I(n2837), .Z(n2836) );
  BUFFD0 U2821 ( .I(n2838), .Z(n2837) );
  BUFFD0 U2822 ( .I(n2839), .Z(n2838) );
  BUFFD0 U2823 ( .I(n2840), .Z(n2839) );
  BUFFD0 U2824 ( .I(n2841), .Z(n2840) );
  BUFFD0 U2825 ( .I(n2842), .Z(n2841) );
  BUFFD0 U2826 ( .I(n2843), .Z(n2842) );
  BUFFD0 U2827 ( .I(n2844), .Z(n2843) );
  BUFFD0 U2828 ( .I(n2845), .Z(n2844) );
  BUFFD0 U2829 ( .I(n2786), .Z(n2845) );
  BUFFD0 U2830 ( .I(n2850), .Z(n2846) );
  BUFFD0 U2831 ( .I(n3956), .Z(n2847) );
  BUFFD0 U2832 ( .I(n2847), .Z(n2848) );
  BUFFD0 U2833 ( .I(n2848), .Z(n2849) );
  BUFFD0 U2834 ( .I(n2851), .Z(n2850) );
  BUFFD0 U2835 ( .I(n2852), .Z(n2851) );
  BUFFD0 U2836 ( .I(n2853), .Z(n2852) );
  BUFFD0 U2837 ( .I(n2854), .Z(n2853) );
  BUFFD0 U2838 ( .I(n2855), .Z(n2854) );
  BUFFD0 U2839 ( .I(n2856), .Z(n2855) );
  BUFFD0 U2840 ( .I(n2857), .Z(n2856) );
  BUFFD0 U2841 ( .I(n2858), .Z(n2857) );
  BUFFD0 U2842 ( .I(n2859), .Z(n2858) );
  BUFFD0 U2843 ( .I(n2860), .Z(n2859) );
  BUFFD0 U2844 ( .I(n2861), .Z(n2860) );
  BUFFD0 U2845 ( .I(n2862), .Z(n2861) );
  BUFFD0 U2846 ( .I(n2863), .Z(n2862) );
  BUFFD0 U2847 ( .I(n2864), .Z(n2863) );
  BUFFD0 U2848 ( .I(n2865), .Z(n2864) );
  BUFFD0 U2849 ( .I(n2866), .Z(n2865) );
  BUFFD0 U2850 ( .I(n2867), .Z(n2866) );
  BUFFD0 U2851 ( .I(n2868), .Z(n2867) );
  BUFFD0 U2852 ( .I(n2869), .Z(n2868) );
  BUFFD0 U2853 ( .I(n2870), .Z(n2869) );
  BUFFD0 U2854 ( .I(n2871), .Z(n2870) );
  BUFFD0 U2855 ( .I(n2872), .Z(n2871) );
  BUFFD0 U2856 ( .I(n2873), .Z(n2872) );
  BUFFD0 U2857 ( .I(n2874), .Z(n2873) );
  BUFFD0 U2858 ( .I(n2875), .Z(n2874) );
  BUFFD0 U2859 ( .I(n2876), .Z(n2875) );
  BUFFD0 U2860 ( .I(n2877), .Z(n2876) );
  BUFFD0 U2861 ( .I(n2878), .Z(n2877) );
  BUFFD0 U2862 ( .I(n2879), .Z(n2878) );
  BUFFD0 U2863 ( .I(n2880), .Z(n2879) );
  BUFFD0 U2864 ( .I(n2881), .Z(n2880) );
  BUFFD0 U2865 ( .I(n2882), .Z(n2881) );
  BUFFD0 U2866 ( .I(n2883), .Z(n2882) );
  BUFFD0 U2867 ( .I(n2884), .Z(n2883) );
  BUFFD0 U2868 ( .I(n2885), .Z(n2884) );
  BUFFD0 U2869 ( .I(n2886), .Z(n2885) );
  BUFFD0 U2870 ( .I(n2887), .Z(n2886) );
  BUFFD0 U2871 ( .I(n2888), .Z(n2887) );
  BUFFD0 U2872 ( .I(n2889), .Z(n2888) );
  BUFFD0 U2873 ( .I(n2890), .Z(n2889) );
  BUFFD0 U2874 ( .I(n2891), .Z(n2890) );
  BUFFD0 U2875 ( .I(n2892), .Z(n2891) );
  BUFFD0 U2876 ( .I(n2893), .Z(n2892) );
  BUFFD0 U2877 ( .I(n2894), .Z(n2893) );
  BUFFD0 U2878 ( .I(n2895), .Z(n2894) );
  BUFFD0 U2879 ( .I(n2896), .Z(n2895) );
  BUFFD0 U2880 ( .I(n2897), .Z(n2896) );
  BUFFD0 U2881 ( .I(n2898), .Z(n2897) );
  BUFFD0 U2882 ( .I(n2899), .Z(n2898) );
  BUFFD0 U2883 ( .I(n2900), .Z(n2899) );
  BUFFD0 U2884 ( .I(n2901), .Z(n2900) );
  BUFFD0 U2885 ( .I(n2902), .Z(n2901) );
  BUFFD0 U2886 ( .I(n2903), .Z(n2902) );
  BUFFD0 U2887 ( .I(n2904), .Z(n2903) );
  BUFFD0 U2888 ( .I(n2905), .Z(n2904) );
  BUFFD0 U2889 ( .I(n2906), .Z(n2905) );
  BUFFD0 U2890 ( .I(n2907), .Z(n2906) );
  BUFFD0 U2891 ( .I(n2908), .Z(n2907) );
  BUFFD0 U2892 ( .I(n2849), .Z(n2908) );
  BUFFD0 U2893 ( .I(n2913), .Z(n2909) );
  BUFFD0 U2894 ( .I(N66), .Z(n2910) );
  BUFFD0 U2895 ( .I(n2910), .Z(n2911) );
  BUFFD0 U2896 ( .I(n2911), .Z(n2912) );
  BUFFD0 U2897 ( .I(n2914), .Z(n2913) );
  BUFFD0 U2898 ( .I(n2915), .Z(n2914) );
  BUFFD0 U2899 ( .I(n2916), .Z(n2915) );
  BUFFD0 U2900 ( .I(n2917), .Z(n2916) );
  BUFFD0 U2901 ( .I(n2918), .Z(n2917) );
  BUFFD0 U2902 ( .I(n2919), .Z(n2918) );
  BUFFD0 U2903 ( .I(n2920), .Z(n2919) );
  BUFFD0 U2904 ( .I(n2921), .Z(n2920) );
  BUFFD0 U2905 ( .I(n2922), .Z(n2921) );
  BUFFD0 U2906 ( .I(n2923), .Z(n2922) );
  BUFFD0 U2907 ( .I(n2924), .Z(n2923) );
  BUFFD0 U2908 ( .I(n2925), .Z(n2924) );
  BUFFD0 U2909 ( .I(n2926), .Z(n2925) );
  BUFFD0 U2910 ( .I(n2927), .Z(n2926) );
  BUFFD0 U2911 ( .I(n2928), .Z(n2927) );
  BUFFD0 U2912 ( .I(n2929), .Z(n2928) );
  BUFFD0 U2913 ( .I(n2930), .Z(n2929) );
  BUFFD0 U2914 ( .I(n2931), .Z(n2930) );
  BUFFD0 U2915 ( .I(n2932), .Z(n2931) );
  BUFFD0 U2916 ( .I(n2933), .Z(n2932) );
  BUFFD0 U2917 ( .I(n2934), .Z(n2933) );
  BUFFD0 U2918 ( .I(n2935), .Z(n2934) );
  BUFFD0 U2919 ( .I(n2936), .Z(n2935) );
  BUFFD0 U2920 ( .I(n2937), .Z(n2936) );
  BUFFD0 U2921 ( .I(n2938), .Z(n2937) );
  BUFFD0 U2922 ( .I(n2939), .Z(n2938) );
  BUFFD0 U2923 ( .I(n2940), .Z(n2939) );
  BUFFD0 U2924 ( .I(n2941), .Z(n2940) );
  BUFFD0 U2925 ( .I(n2942), .Z(n2941) );
  BUFFD0 U2926 ( .I(n2943), .Z(n2942) );
  BUFFD0 U2927 ( .I(n2944), .Z(n2943) );
  BUFFD0 U2928 ( .I(n2945), .Z(n2944) );
  BUFFD0 U2929 ( .I(n2946), .Z(n2945) );
  BUFFD0 U2930 ( .I(n2947), .Z(n2946) );
  BUFFD0 U2931 ( .I(n2948), .Z(n2947) );
  BUFFD0 U2932 ( .I(n2949), .Z(n2948) );
  BUFFD0 U2933 ( .I(n2950), .Z(n2949) );
  BUFFD0 U2934 ( .I(n2951), .Z(n2950) );
  BUFFD0 U2935 ( .I(n2952), .Z(n2951) );
  BUFFD0 U2936 ( .I(n2953), .Z(n2952) );
  BUFFD0 U2937 ( .I(n2954), .Z(n2953) );
  BUFFD0 U2938 ( .I(n2955), .Z(n2954) );
  BUFFD0 U2939 ( .I(n2956), .Z(n2955) );
  BUFFD0 U2940 ( .I(n2957), .Z(n2956) );
  BUFFD0 U2941 ( .I(n2958), .Z(n2957) );
  BUFFD0 U2942 ( .I(n2959), .Z(n2958) );
  BUFFD0 U2943 ( .I(n2960), .Z(n2959) );
  BUFFD0 U2944 ( .I(n2961), .Z(n2960) );
  BUFFD0 U2945 ( .I(n2962), .Z(n2961) );
  BUFFD0 U2946 ( .I(n2963), .Z(n2962) );
  BUFFD0 U2947 ( .I(n2964), .Z(n2963) );
  BUFFD0 U2948 ( .I(n2965), .Z(n2964) );
  BUFFD0 U2949 ( .I(n2966), .Z(n2965) );
  BUFFD0 U2950 ( .I(n2967), .Z(n2966) );
  BUFFD0 U2951 ( .I(n2968), .Z(n2967) );
  BUFFD0 U2952 ( .I(n2969), .Z(n2968) );
  BUFFD0 U2953 ( .I(n2970), .Z(n2969) );
  BUFFD0 U2954 ( .I(n3960), .Z(n2970) );
  BUFFD0 U2955 ( .I(n2912), .Z(n2971) );
  BUFFD0 U2956 ( .I(n2976), .Z(n2972) );
  BUFFD0 U2957 ( .I(N67), .Z(n2973) );
  BUFFD0 U2958 ( .I(n2973), .Z(n2974) );
  BUFFD0 U2959 ( .I(n2974), .Z(n2975) );
  BUFFD0 U2960 ( .I(n2977), .Z(n2976) );
  BUFFD0 U2961 ( .I(n2978), .Z(n2977) );
  BUFFD0 U2962 ( .I(n2979), .Z(n2978) );
  BUFFD0 U2963 ( .I(n2980), .Z(n2979) );
  BUFFD0 U2964 ( .I(n2981), .Z(n2980) );
  BUFFD0 U2965 ( .I(n2982), .Z(n2981) );
  BUFFD0 U2966 ( .I(n2983), .Z(n2982) );
  BUFFD0 U2967 ( .I(n2984), .Z(n2983) );
  BUFFD0 U2968 ( .I(n2985), .Z(n2984) );
  BUFFD0 U2969 ( .I(n2986), .Z(n2985) );
  BUFFD0 U2970 ( .I(n2987), .Z(n2986) );
  BUFFD0 U2971 ( .I(n2988), .Z(n2987) );
  BUFFD0 U2972 ( .I(n2989), .Z(n2988) );
  BUFFD0 U2973 ( .I(n2990), .Z(n2989) );
  BUFFD0 U2974 ( .I(n2991), .Z(n2990) );
  BUFFD0 U2975 ( .I(n2992), .Z(n2991) );
  BUFFD0 U2976 ( .I(n2993), .Z(n2992) );
  BUFFD0 U2977 ( .I(n2994), .Z(n2993) );
  BUFFD0 U2978 ( .I(n2995), .Z(n2994) );
  BUFFD0 U2979 ( .I(n2996), .Z(n2995) );
  BUFFD0 U2980 ( .I(n2997), .Z(n2996) );
  BUFFD0 U2981 ( .I(n2998), .Z(n2997) );
  BUFFD0 U2982 ( .I(n2999), .Z(n2998) );
  BUFFD0 U2983 ( .I(n3000), .Z(n2999) );
  BUFFD0 U2984 ( .I(n3001), .Z(n3000) );
  BUFFD0 U2985 ( .I(n3002), .Z(n3001) );
  BUFFD0 U2986 ( .I(n3003), .Z(n3002) );
  BUFFD0 U2987 ( .I(n3004), .Z(n3003) );
  BUFFD0 U2988 ( .I(n3005), .Z(n3004) );
  BUFFD0 U2989 ( .I(n3006), .Z(n3005) );
  BUFFD0 U2990 ( .I(n3007), .Z(n3006) );
  BUFFD0 U2991 ( .I(n3008), .Z(n3007) );
  BUFFD0 U2992 ( .I(n3009), .Z(n3008) );
  BUFFD0 U2993 ( .I(n3010), .Z(n3009) );
  BUFFD0 U2994 ( .I(n3011), .Z(n3010) );
  BUFFD0 U2995 ( .I(n3012), .Z(n3011) );
  BUFFD0 U2996 ( .I(n3013), .Z(n3012) );
  BUFFD0 U2997 ( .I(n3014), .Z(n3013) );
  BUFFD0 U2998 ( .I(n3015), .Z(n3014) );
  BUFFD0 U2999 ( .I(n3016), .Z(n3015) );
  BUFFD0 U3000 ( .I(n3017), .Z(n3016) );
  BUFFD0 U3001 ( .I(n3018), .Z(n3017) );
  BUFFD0 U3002 ( .I(n3019), .Z(n3018) );
  BUFFD0 U3003 ( .I(n3020), .Z(n3019) );
  BUFFD0 U3004 ( .I(n3021), .Z(n3020) );
  BUFFD0 U3005 ( .I(n3022), .Z(n3021) );
  BUFFD0 U3006 ( .I(n3023), .Z(n3022) );
  BUFFD0 U3007 ( .I(n3024), .Z(n3023) );
  BUFFD0 U3008 ( .I(n3025), .Z(n3024) );
  BUFFD0 U3009 ( .I(n3026), .Z(n3025) );
  BUFFD0 U3010 ( .I(n3027), .Z(n3026) );
  BUFFD0 U3011 ( .I(n3028), .Z(n3027) );
  BUFFD0 U3012 ( .I(n3029), .Z(n3028) );
  BUFFD0 U3013 ( .I(n3030), .Z(n3029) );
  BUFFD0 U3014 ( .I(n3031), .Z(n3030) );
  BUFFD0 U3015 ( .I(n3032), .Z(n3031) );
  BUFFD0 U3016 ( .I(n3033), .Z(n3032) );
  BUFFD0 U3017 ( .I(n3971), .Z(n3033) );
  BUFFD0 U3018 ( .I(n3038), .Z(n3034) );
  BUFFD0 U3019 ( .I(n3965), .Z(n3035) );
  BUFFD0 U3020 ( .I(n3035), .Z(n3036) );
  BUFFD0 U3021 ( .I(n3036), .Z(n3037) );
  BUFFD0 U3022 ( .I(n3039), .Z(n3038) );
  BUFFD0 U3023 ( .I(n3040), .Z(n3039) );
  BUFFD0 U3024 ( .I(n3041), .Z(n3040) );
  BUFFD0 U3025 ( .I(n3042), .Z(n3041) );
  BUFFD0 U3026 ( .I(n3043), .Z(n3042) );
  BUFFD0 U3027 ( .I(n3044), .Z(n3043) );
  BUFFD0 U3028 ( .I(n3045), .Z(n3044) );
  BUFFD0 U3029 ( .I(n3046), .Z(n3045) );
  BUFFD0 U3030 ( .I(n3047), .Z(n3046) );
  BUFFD0 U3031 ( .I(n3048), .Z(n3047) );
  BUFFD0 U3032 ( .I(n3049), .Z(n3048) );
  BUFFD0 U3033 ( .I(n3050), .Z(n3049) );
  BUFFD0 U3034 ( .I(n3051), .Z(n3050) );
  BUFFD0 U3035 ( .I(n3052), .Z(n3051) );
  BUFFD0 U3036 ( .I(n3053), .Z(n3052) );
  BUFFD0 U3037 ( .I(n3054), .Z(n3053) );
  BUFFD0 U3038 ( .I(n3055), .Z(n3054) );
  BUFFD0 U3039 ( .I(n3056), .Z(n3055) );
  BUFFD0 U3040 ( .I(n3057), .Z(n3056) );
  BUFFD0 U3041 ( .I(n3058), .Z(n3057) );
  BUFFD0 U3042 ( .I(n3059), .Z(n3058) );
  BUFFD0 U3043 ( .I(n3060), .Z(n3059) );
  BUFFD0 U3044 ( .I(n3061), .Z(n3060) );
  BUFFD0 U3045 ( .I(n3062), .Z(n3061) );
  BUFFD0 U3046 ( .I(n3063), .Z(n3062) );
  BUFFD0 U3047 ( .I(n3064), .Z(n3063) );
  BUFFD0 U3048 ( .I(n3065), .Z(n3064) );
  BUFFD0 U3049 ( .I(n3066), .Z(n3065) );
  BUFFD0 U3050 ( .I(n3067), .Z(n3066) );
  BUFFD0 U3051 ( .I(n3068), .Z(n3067) );
  BUFFD0 U3052 ( .I(n3069), .Z(n3068) );
  BUFFD0 U3053 ( .I(n3070), .Z(n3069) );
  BUFFD0 U3054 ( .I(n3071), .Z(n3070) );
  BUFFD0 U3055 ( .I(n3072), .Z(n3071) );
  BUFFD0 U3056 ( .I(n3073), .Z(n3072) );
  BUFFD0 U3057 ( .I(n3074), .Z(n3073) );
  BUFFD0 U3058 ( .I(n3075), .Z(n3074) );
  BUFFD0 U3059 ( .I(n3076), .Z(n3075) );
  BUFFD0 U3060 ( .I(n3077), .Z(n3076) );
  BUFFD0 U3061 ( .I(n3078), .Z(n3077) );
  BUFFD0 U3062 ( .I(n3079), .Z(n3078) );
  BUFFD0 U3063 ( .I(n3080), .Z(n3079) );
  BUFFD0 U3064 ( .I(n3081), .Z(n3080) );
  BUFFD0 U3065 ( .I(n3082), .Z(n3081) );
  BUFFD0 U3066 ( .I(n3083), .Z(n3082) );
  BUFFD0 U3067 ( .I(n3084), .Z(n3083) );
  BUFFD0 U3068 ( .I(n3085), .Z(n3084) );
  BUFFD0 U3069 ( .I(n3086), .Z(n3085) );
  BUFFD0 U3070 ( .I(n3087), .Z(n3086) );
  BUFFD0 U3071 ( .I(n3088), .Z(n3087) );
  BUFFD0 U3072 ( .I(n3089), .Z(n3088) );
  BUFFD0 U3073 ( .I(n3090), .Z(n3089) );
  BUFFD0 U3074 ( .I(n3091), .Z(n3090) );
  BUFFD0 U3075 ( .I(n3092), .Z(n3091) );
  BUFFD0 U3076 ( .I(n3093), .Z(n3092) );
  BUFFD0 U3077 ( .I(n3094), .Z(n3093) );
  BUFFD0 U3078 ( .I(n3095), .Z(n3094) );
  BUFFD0 U3079 ( .I(n3037), .Z(n3095) );
  BUFFD0 U3080 ( .I(n3100), .Z(n3096) );
  BUFFD0 U3081 ( .I(n3961), .Z(n3097) );
  BUFFD0 U3082 ( .I(n3097), .Z(n3098) );
  BUFFD0 U3083 ( .I(n3098), .Z(n3099) );
  BUFFD0 U3084 ( .I(n3101), .Z(n3100) );
  BUFFD0 U3085 ( .I(n3102), .Z(n3101) );
  BUFFD0 U3086 ( .I(n3103), .Z(n3102) );
  BUFFD0 U3087 ( .I(n3104), .Z(n3103) );
  BUFFD0 U3088 ( .I(n3105), .Z(n3104) );
  BUFFD0 U3089 ( .I(n3106), .Z(n3105) );
  BUFFD0 U3090 ( .I(n3107), .Z(n3106) );
  BUFFD0 U3091 ( .I(n3108), .Z(n3107) );
  BUFFD0 U3092 ( .I(n3109), .Z(n3108) );
  BUFFD0 U3093 ( .I(n3110), .Z(n3109) );
  BUFFD0 U3094 ( .I(n3111), .Z(n3110) );
  BUFFD0 U3095 ( .I(n3112), .Z(n3111) );
  BUFFD0 U3096 ( .I(n3113), .Z(n3112) );
  BUFFD0 U3097 ( .I(n3114), .Z(n3113) );
  BUFFD0 U3098 ( .I(n3115), .Z(n3114) );
  BUFFD0 U3099 ( .I(n3116), .Z(n3115) );
  BUFFD0 U3100 ( .I(n3117), .Z(n3116) );
  BUFFD0 U3101 ( .I(n3118), .Z(n3117) );
  BUFFD0 U3102 ( .I(n3119), .Z(n3118) );
  BUFFD0 U3103 ( .I(n3120), .Z(n3119) );
  BUFFD0 U3104 ( .I(n3121), .Z(n3120) );
  BUFFD0 U3105 ( .I(n3122), .Z(n3121) );
  BUFFD0 U3106 ( .I(n3123), .Z(n3122) );
  BUFFD0 U3107 ( .I(n3124), .Z(n3123) );
  BUFFD0 U3108 ( .I(n3125), .Z(n3124) );
  BUFFD0 U3109 ( .I(n3126), .Z(n3125) );
  BUFFD0 U3110 ( .I(n3127), .Z(n3126) );
  BUFFD0 U3111 ( .I(n3128), .Z(n3127) );
  BUFFD0 U3112 ( .I(n3129), .Z(n3128) );
  BUFFD0 U3113 ( .I(n3130), .Z(n3129) );
  BUFFD0 U3114 ( .I(n3131), .Z(n3130) );
  BUFFD0 U3115 ( .I(n3132), .Z(n3131) );
  BUFFD0 U3116 ( .I(n3133), .Z(n3132) );
  BUFFD0 U3117 ( .I(n3134), .Z(n3133) );
  BUFFD0 U3118 ( .I(n3135), .Z(n3134) );
  BUFFD0 U3119 ( .I(n3136), .Z(n3135) );
  BUFFD0 U3120 ( .I(n3137), .Z(n3136) );
  BUFFD0 U3121 ( .I(n3138), .Z(n3137) );
  BUFFD0 U3122 ( .I(n3139), .Z(n3138) );
  BUFFD0 U3123 ( .I(n3140), .Z(n3139) );
  BUFFD0 U3124 ( .I(n3141), .Z(n3140) );
  BUFFD0 U3125 ( .I(n3142), .Z(n3141) );
  BUFFD0 U3126 ( .I(n3143), .Z(n3142) );
  BUFFD0 U3127 ( .I(n3144), .Z(n3143) );
  BUFFD0 U3128 ( .I(n3145), .Z(n3144) );
  BUFFD0 U3129 ( .I(n3146), .Z(n3145) );
  BUFFD0 U3130 ( .I(n3147), .Z(n3146) );
  BUFFD0 U3131 ( .I(n3148), .Z(n3147) );
  BUFFD0 U3132 ( .I(n3149), .Z(n3148) );
  BUFFD0 U3133 ( .I(n3150), .Z(n3149) );
  BUFFD0 U3134 ( .I(n3151), .Z(n3150) );
  BUFFD0 U3135 ( .I(n3152), .Z(n3151) );
  BUFFD0 U3136 ( .I(n3153), .Z(n3152) );
  BUFFD0 U3137 ( .I(n3154), .Z(n3153) );
  BUFFD0 U3138 ( .I(n3155), .Z(n3154) );
  BUFFD0 U3139 ( .I(n3156), .Z(n3155) );
  BUFFD0 U3140 ( .I(n3157), .Z(n3156) );
  BUFFD0 U3141 ( .I(n3158), .Z(n3157) );
  BUFFD0 U3142 ( .I(n3099), .Z(n3158) );
  BUFFD0 U3143 ( .I(n3163), .Z(n3159) );
  BUFFD0 U3144 ( .I(N70), .Z(n3160) );
  BUFFD0 U3145 ( .I(n3160), .Z(n3161) );
  BUFFD0 U3146 ( .I(n3161), .Z(n3162) );
  BUFFD0 U3147 ( .I(n3164), .Z(n3163) );
  BUFFD0 U3148 ( .I(n3165), .Z(n3164) );
  BUFFD0 U3149 ( .I(n3166), .Z(n3165) );
  BUFFD0 U3150 ( .I(n3167), .Z(n3166) );
  BUFFD0 U3151 ( .I(n3168), .Z(n3167) );
  BUFFD0 U3152 ( .I(n3169), .Z(n3168) );
  BUFFD0 U3153 ( .I(n3170), .Z(n3169) );
  BUFFD0 U3154 ( .I(n3171), .Z(n3170) );
  BUFFD0 U3155 ( .I(n3172), .Z(n3171) );
  BUFFD0 U3156 ( .I(n3173), .Z(n3172) );
  BUFFD0 U3157 ( .I(n3174), .Z(n3173) );
  BUFFD0 U3158 ( .I(n3175), .Z(n3174) );
  BUFFD0 U3159 ( .I(n3176), .Z(n3175) );
  BUFFD0 U3160 ( .I(n3177), .Z(n3176) );
  BUFFD0 U3161 ( .I(n3178), .Z(n3177) );
  BUFFD0 U3162 ( .I(n3179), .Z(n3178) );
  BUFFD0 U3163 ( .I(n3180), .Z(n3179) );
  BUFFD0 U3164 ( .I(n3181), .Z(n3180) );
  BUFFD0 U3165 ( .I(n3182), .Z(n3181) );
  BUFFD0 U3166 ( .I(n3183), .Z(n3182) );
  BUFFD0 U3167 ( .I(n3184), .Z(n3183) );
  BUFFD0 U3168 ( .I(n3185), .Z(n3184) );
  BUFFD0 U3169 ( .I(n3186), .Z(n3185) );
  BUFFD0 U3170 ( .I(n3187), .Z(n3186) );
  BUFFD0 U3171 ( .I(n3188), .Z(n3187) );
  BUFFD0 U3172 ( .I(n3189), .Z(n3188) );
  BUFFD0 U3173 ( .I(n3190), .Z(n3189) );
  BUFFD0 U3174 ( .I(n3191), .Z(n3190) );
  BUFFD0 U3175 ( .I(n3192), .Z(n3191) );
  BUFFD0 U3176 ( .I(n3193), .Z(n3192) );
  BUFFD0 U3177 ( .I(n3194), .Z(n3193) );
  BUFFD0 U3178 ( .I(n3195), .Z(n3194) );
  BUFFD0 U3179 ( .I(n3196), .Z(n3195) );
  BUFFD0 U3180 ( .I(n3197), .Z(n3196) );
  BUFFD0 U3181 ( .I(n3198), .Z(n3197) );
  BUFFD0 U3182 ( .I(n3199), .Z(n3198) );
  BUFFD0 U3183 ( .I(n3200), .Z(n3199) );
  BUFFD0 U3184 ( .I(n3201), .Z(n3200) );
  BUFFD0 U3185 ( .I(n3202), .Z(n3201) );
  BUFFD0 U3186 ( .I(n3203), .Z(n3202) );
  BUFFD0 U3187 ( .I(n3204), .Z(n3203) );
  BUFFD0 U3188 ( .I(n3205), .Z(n3204) );
  BUFFD0 U3189 ( .I(n3206), .Z(n3205) );
  BUFFD0 U3190 ( .I(n3207), .Z(n3206) );
  BUFFD0 U3191 ( .I(n3208), .Z(n3207) );
  BUFFD0 U3192 ( .I(n3209), .Z(n3208) );
  BUFFD0 U3193 ( .I(n3210), .Z(n3209) );
  BUFFD0 U3194 ( .I(n3211), .Z(n3210) );
  BUFFD0 U3195 ( .I(n3212), .Z(n3211) );
  BUFFD0 U3196 ( .I(n3213), .Z(n3212) );
  BUFFD0 U3197 ( .I(n3214), .Z(n3213) );
  BUFFD0 U3198 ( .I(n3215), .Z(n3214) );
  BUFFD0 U3199 ( .I(n3216), .Z(n3215) );
  BUFFD0 U3200 ( .I(n3217), .Z(n3216) );
  BUFFD0 U3201 ( .I(n3218), .Z(n3217) );
  BUFFD0 U3202 ( .I(n3219), .Z(n3218) );
  BUFFD0 U3203 ( .I(n3220), .Z(n3219) );
  BUFFD0 U3204 ( .I(n3963), .Z(n3220) );
  BUFFD0 U3205 ( .I(n3162), .Z(n3221) );
  BUFFD0 U3206 ( .I(n3226), .Z(n3222) );
  BUFFD0 U3207 ( .I(N71), .Z(n3223) );
  BUFFD0 U3208 ( .I(n3223), .Z(n3224) );
  BUFFD0 U3209 ( .I(n3224), .Z(n3225) );
  BUFFD0 U3210 ( .I(n3227), .Z(n3226) );
  BUFFD0 U3211 ( .I(n3228), .Z(n3227) );
  BUFFD0 U3212 ( .I(n3229), .Z(n3228) );
  BUFFD0 U3213 ( .I(n3230), .Z(n3229) );
  BUFFD0 U3214 ( .I(n3231), .Z(n3230) );
  BUFFD0 U3215 ( .I(n3232), .Z(n3231) );
  BUFFD0 U3216 ( .I(n3233), .Z(n3232) );
  BUFFD0 U3217 ( .I(n3234), .Z(n3233) );
  BUFFD0 U3218 ( .I(n3235), .Z(n3234) );
  BUFFD0 U3219 ( .I(n3236), .Z(n3235) );
  BUFFD0 U3220 ( .I(n3237), .Z(n3236) );
  BUFFD0 U3221 ( .I(n3238), .Z(n3237) );
  BUFFD0 U3222 ( .I(n3239), .Z(n3238) );
  BUFFD0 U3223 ( .I(n3240), .Z(n3239) );
  BUFFD0 U3224 ( .I(n3241), .Z(n3240) );
  BUFFD0 U3225 ( .I(n3242), .Z(n3241) );
  BUFFD0 U3226 ( .I(n3243), .Z(n3242) );
  BUFFD0 U3227 ( .I(n3244), .Z(n3243) );
  BUFFD0 U3228 ( .I(n3245), .Z(n3244) );
  BUFFD0 U3229 ( .I(n3246), .Z(n3245) );
  BUFFD0 U3230 ( .I(n3247), .Z(n3246) );
  BUFFD0 U3231 ( .I(n3248), .Z(n3247) );
  BUFFD0 U3232 ( .I(n3249), .Z(n3248) );
  BUFFD0 U3233 ( .I(n3250), .Z(n3249) );
  BUFFD0 U3234 ( .I(n3251), .Z(n3250) );
  BUFFD0 U3235 ( .I(n3252), .Z(n3251) );
  BUFFD0 U3236 ( .I(n3253), .Z(n3252) );
  BUFFD0 U3237 ( .I(n3254), .Z(n3253) );
  BUFFD0 U3238 ( .I(n3255), .Z(n3254) );
  BUFFD0 U3239 ( .I(n3256), .Z(n3255) );
  BUFFD0 U3240 ( .I(n3257), .Z(n3256) );
  BUFFD0 U3241 ( .I(n3258), .Z(n3257) );
  BUFFD0 U3242 ( .I(n3259), .Z(n3258) );
  BUFFD0 U3243 ( .I(n3260), .Z(n3259) );
  BUFFD0 U3244 ( .I(n3261), .Z(n3260) );
  BUFFD0 U3245 ( .I(n3262), .Z(n3261) );
  BUFFD0 U3246 ( .I(n3263), .Z(n3262) );
  BUFFD0 U3247 ( .I(n3264), .Z(n3263) );
  BUFFD0 U3248 ( .I(n3265), .Z(n3264) );
  BUFFD0 U3249 ( .I(n3266), .Z(n3265) );
  BUFFD0 U3250 ( .I(n3267), .Z(n3266) );
  BUFFD0 U3251 ( .I(n3268), .Z(n3267) );
  BUFFD0 U3252 ( .I(n3269), .Z(n3268) );
  BUFFD0 U3253 ( .I(n3270), .Z(n3269) );
  BUFFD0 U3254 ( .I(n3271), .Z(n3270) );
  BUFFD0 U3255 ( .I(n3272), .Z(n3271) );
  BUFFD0 U3256 ( .I(n3273), .Z(n3272) );
  BUFFD0 U3257 ( .I(n3274), .Z(n3273) );
  BUFFD0 U3258 ( .I(n3275), .Z(n3274) );
  BUFFD0 U3259 ( .I(n3276), .Z(n3275) );
  BUFFD0 U3260 ( .I(n3277), .Z(n3276) );
  BUFFD0 U3261 ( .I(n3278), .Z(n3277) );
  BUFFD0 U3262 ( .I(n3279), .Z(n3278) );
  BUFFD0 U3263 ( .I(n3280), .Z(n3279) );
  BUFFD0 U3264 ( .I(n3281), .Z(n3280) );
  BUFFD0 U3265 ( .I(n3282), .Z(n3281) );
  BUFFD0 U3266 ( .I(n4002), .Z(n3282) );
  BUFFD0 U3267 ( .I(n3287), .Z(n3283) );
  BUFFD0 U3268 ( .I(N72), .Z(n3284) );
  BUFFD0 U3269 ( .I(n3284), .Z(n3285) );
  BUFFD0 U3270 ( .I(n3285), .Z(n3286) );
  BUFFD0 U3271 ( .I(n3288), .Z(n3287) );
  BUFFD0 U3272 ( .I(n3289), .Z(n3288) );
  BUFFD0 U3273 ( .I(n3290), .Z(n3289) );
  BUFFD0 U3274 ( .I(n3291), .Z(n3290) );
  BUFFD0 U3275 ( .I(n3292), .Z(n3291) );
  BUFFD0 U3276 ( .I(n3293), .Z(n3292) );
  BUFFD0 U3277 ( .I(n3294), .Z(n3293) );
  BUFFD0 U3278 ( .I(n3295), .Z(n3294) );
  BUFFD0 U3279 ( .I(n3296), .Z(n3295) );
  BUFFD0 U3280 ( .I(n3297), .Z(n3296) );
  BUFFD0 U3281 ( .I(n3298), .Z(n3297) );
  BUFFD0 U3282 ( .I(n3299), .Z(n3298) );
  BUFFD0 U3283 ( .I(n3300), .Z(n3299) );
  BUFFD0 U3284 ( .I(n3301), .Z(n3300) );
  BUFFD0 U3285 ( .I(n3302), .Z(n3301) );
  BUFFD0 U3286 ( .I(n3303), .Z(n3302) );
  BUFFD0 U3287 ( .I(n3304), .Z(n3303) );
  BUFFD0 U3288 ( .I(n3305), .Z(n3304) );
  BUFFD0 U3289 ( .I(n3306), .Z(n3305) );
  BUFFD0 U3290 ( .I(n3307), .Z(n3306) );
  BUFFD0 U3291 ( .I(n3308), .Z(n3307) );
  BUFFD0 U3292 ( .I(n3309), .Z(n3308) );
  BUFFD0 U3293 ( .I(n3310), .Z(n3309) );
  BUFFD0 U3294 ( .I(n3311), .Z(n3310) );
  BUFFD0 U3295 ( .I(n3312), .Z(n3311) );
  BUFFD0 U3296 ( .I(n3313), .Z(n3312) );
  BUFFD0 U3297 ( .I(n3314), .Z(n3313) );
  BUFFD0 U3298 ( .I(n3315), .Z(n3314) );
  BUFFD0 U3299 ( .I(n3316), .Z(n3315) );
  BUFFD0 U3300 ( .I(n3317), .Z(n3316) );
  BUFFD0 U3301 ( .I(n3318), .Z(n3317) );
  BUFFD0 U3302 ( .I(n3319), .Z(n3318) );
  BUFFD0 U3303 ( .I(n3320), .Z(n3319) );
  BUFFD0 U3304 ( .I(n3321), .Z(n3320) );
  BUFFD0 U3305 ( .I(n3322), .Z(n3321) );
  BUFFD0 U3306 ( .I(n3323), .Z(n3322) );
  BUFFD0 U3307 ( .I(n3324), .Z(n3323) );
  BUFFD0 U3308 ( .I(n3325), .Z(n3324) );
  BUFFD0 U3309 ( .I(n3326), .Z(n3325) );
  BUFFD0 U3310 ( .I(n3327), .Z(n3326) );
  BUFFD0 U3311 ( .I(n3328), .Z(n3327) );
  BUFFD0 U3312 ( .I(n3329), .Z(n3328) );
  BUFFD0 U3313 ( .I(n3330), .Z(n3329) );
  BUFFD0 U3314 ( .I(n3331), .Z(n3330) );
  BUFFD0 U3315 ( .I(n3332), .Z(n3331) );
  BUFFD0 U3316 ( .I(n3333), .Z(n3332) );
  BUFFD0 U3317 ( .I(n3334), .Z(n3333) );
  BUFFD0 U3318 ( .I(n3335), .Z(n3334) );
  BUFFD0 U3319 ( .I(n3336), .Z(n3335) );
  BUFFD0 U3320 ( .I(n3337), .Z(n3336) );
  BUFFD0 U3321 ( .I(n3338), .Z(n3337) );
  BUFFD0 U3322 ( .I(n3339), .Z(n3338) );
  BUFFD0 U3323 ( .I(n3340), .Z(n3339) );
  BUFFD0 U3324 ( .I(n4031), .Z(n3340) );
  BUFFD0 U3325 ( .I(n3345), .Z(n3341) );
  BUFFD0 U3326 ( .I(n4037), .Z(n3342) );
  BUFFD0 U3327 ( .I(n3342), .Z(n3343) );
  BUFFD0 U3328 ( .I(n3343), .Z(n3344) );
  BUFFD0 U3329 ( .I(n3346), .Z(n3345) );
  BUFFD0 U3330 ( .I(n3347), .Z(n3346) );
  BUFFD0 U3331 ( .I(n3348), .Z(n3347) );
  BUFFD0 U3332 ( .I(n3349), .Z(n3348) );
  BUFFD0 U3333 ( .I(n3350), .Z(n3349) );
  BUFFD0 U3334 ( .I(n3351), .Z(n3350) );
  BUFFD0 U3335 ( .I(n3352), .Z(n3351) );
  BUFFD0 U3336 ( .I(n3353), .Z(n3352) );
  BUFFD0 U3337 ( .I(n3354), .Z(n3353) );
  BUFFD0 U3338 ( .I(n3355), .Z(n3354) );
  BUFFD0 U3339 ( .I(n3356), .Z(n3355) );
  BUFFD0 U3340 ( .I(n3357), .Z(n3356) );
  BUFFD0 U3341 ( .I(n3358), .Z(n3357) );
  BUFFD0 U3342 ( .I(n3359), .Z(n3358) );
  BUFFD0 U3343 ( .I(n3360), .Z(n3359) );
  BUFFD0 U3344 ( .I(n3361), .Z(n3360) );
  BUFFD0 U3345 ( .I(n3362), .Z(n3361) );
  BUFFD0 U3346 ( .I(n3363), .Z(n3362) );
  BUFFD0 U3347 ( .I(n3364), .Z(n3363) );
  BUFFD0 U3348 ( .I(n3365), .Z(n3364) );
  BUFFD0 U3349 ( .I(n3366), .Z(n3365) );
  BUFFD0 U3350 ( .I(n3367), .Z(n3366) );
  BUFFD0 U3351 ( .I(n3368), .Z(n3367) );
  BUFFD0 U3352 ( .I(n3369), .Z(n3368) );
  BUFFD0 U3353 ( .I(n3370), .Z(n3369) );
  BUFFD0 U3354 ( .I(n3371), .Z(n3370) );
  BUFFD0 U3355 ( .I(n3372), .Z(n3371) );
  BUFFD0 U3356 ( .I(n3373), .Z(n3372) );
  BUFFD0 U3357 ( .I(n3374), .Z(n3373) );
  BUFFD0 U3358 ( .I(n3375), .Z(n3374) );
  BUFFD0 U3359 ( .I(n3376), .Z(n3375) );
  BUFFD0 U3360 ( .I(n3377), .Z(n3376) );
  BUFFD0 U3361 ( .I(n3378), .Z(n3377) );
  BUFFD0 U3362 ( .I(n3379), .Z(n3378) );
  BUFFD0 U3363 ( .I(n3380), .Z(n3379) );
  BUFFD0 U3364 ( .I(n3381), .Z(n3380) );
  BUFFD0 U3365 ( .I(n3382), .Z(n3381) );
  BUFFD0 U3366 ( .I(n3383), .Z(n3382) );
  BUFFD0 U3367 ( .I(n3384), .Z(n3383) );
  BUFFD0 U3368 ( .I(n3385), .Z(n3384) );
  BUFFD0 U3369 ( .I(n3386), .Z(n3385) );
  BUFFD0 U3370 ( .I(n3387), .Z(n3386) );
  BUFFD0 U3371 ( .I(n3388), .Z(n3387) );
  BUFFD0 U3372 ( .I(n3389), .Z(n3388) );
  BUFFD0 U3373 ( .I(n3390), .Z(n3389) );
  BUFFD0 U3374 ( .I(n3391), .Z(n3390) );
  BUFFD0 U3375 ( .I(n3392), .Z(n3391) );
  BUFFD0 U3376 ( .I(n3393), .Z(n3392) );
  BUFFD0 U3377 ( .I(n3394), .Z(n3393) );
  BUFFD0 U3378 ( .I(n3395), .Z(n3394) );
  BUFFD0 U3379 ( .I(n3396), .Z(n3395) );
  BUFFD0 U3380 ( .I(n3397), .Z(n3396) );
  BUFFD0 U3381 ( .I(n3344), .Z(n3397) );
  BUFFD0 U3382 ( .I(n3402), .Z(n3398) );
  BUFFD0 U3383 ( .I(n4001), .Z(n3399) );
  BUFFD0 U3384 ( .I(n3399), .Z(n3400) );
  BUFFD0 U3385 ( .I(n3400), .Z(n3401) );
  BUFFD0 U3386 ( .I(n3403), .Z(n3402) );
  BUFFD0 U3387 ( .I(n3404), .Z(n3403) );
  BUFFD0 U3388 ( .I(n3405), .Z(n3404) );
  BUFFD0 U3389 ( .I(n3406), .Z(n3405) );
  BUFFD0 U3390 ( .I(n3407), .Z(n3406) );
  BUFFD0 U3391 ( .I(n3408), .Z(n3407) );
  BUFFD0 U3392 ( .I(n3409), .Z(n3408) );
  BUFFD0 U3393 ( .I(n3410), .Z(n3409) );
  BUFFD0 U3394 ( .I(n3411), .Z(n3410) );
  BUFFD0 U3395 ( .I(n3412), .Z(n3411) );
  BUFFD0 U3396 ( .I(n3413), .Z(n3412) );
  BUFFD0 U3397 ( .I(n3414), .Z(n3413) );
  BUFFD0 U3398 ( .I(n3415), .Z(n3414) );
  BUFFD0 U3399 ( .I(n3416), .Z(n3415) );
  BUFFD0 U3400 ( .I(n3417), .Z(n3416) );
  BUFFD0 U3401 ( .I(n3418), .Z(n3417) );
  BUFFD0 U3402 ( .I(n3419), .Z(n3418) );
  BUFFD0 U3403 ( .I(n3420), .Z(n3419) );
  BUFFD0 U3404 ( .I(n3421), .Z(n3420) );
  BUFFD0 U3405 ( .I(n3422), .Z(n3421) );
  BUFFD0 U3406 ( .I(n3423), .Z(n3422) );
  BUFFD0 U3407 ( .I(n3424), .Z(n3423) );
  BUFFD0 U3408 ( .I(n3425), .Z(n3424) );
  BUFFD0 U3409 ( .I(n3426), .Z(n3425) );
  BUFFD0 U3410 ( .I(n3427), .Z(n3426) );
  BUFFD0 U3411 ( .I(n3428), .Z(n3427) );
  BUFFD0 U3412 ( .I(n3429), .Z(n3428) );
  BUFFD0 U3413 ( .I(n3430), .Z(n3429) );
  BUFFD0 U3414 ( .I(n3431), .Z(n3430) );
  BUFFD0 U3415 ( .I(n3432), .Z(n3431) );
  BUFFD0 U3416 ( .I(n3433), .Z(n3432) );
  BUFFD0 U3417 ( .I(n3434), .Z(n3433) );
  BUFFD0 U3418 ( .I(n3435), .Z(n3434) );
  BUFFD0 U3419 ( .I(n3436), .Z(n3435) );
  BUFFD0 U3420 ( .I(n3437), .Z(n3436) );
  BUFFD0 U3421 ( .I(n3438), .Z(n3437) );
  BUFFD0 U3422 ( .I(n3439), .Z(n3438) );
  BUFFD0 U3423 ( .I(n3440), .Z(n3439) );
  BUFFD0 U3424 ( .I(n3441), .Z(n3440) );
  BUFFD0 U3425 ( .I(n3442), .Z(n3441) );
  BUFFD0 U3426 ( .I(n3443), .Z(n3442) );
  BUFFD0 U3427 ( .I(n3444), .Z(n3443) );
  BUFFD0 U3428 ( .I(n3445), .Z(n3444) );
  BUFFD0 U3429 ( .I(n3446), .Z(n3445) );
  BUFFD0 U3430 ( .I(n3447), .Z(n3446) );
  BUFFD0 U3431 ( .I(n3448), .Z(n3447) );
  BUFFD0 U3432 ( .I(n3449), .Z(n3448) );
  BUFFD0 U3433 ( .I(n3450), .Z(n3449) );
  BUFFD0 U3434 ( .I(n3451), .Z(n3450) );
  BUFFD0 U3435 ( .I(n3452), .Z(n3451) );
  BUFFD0 U3436 ( .I(n3453), .Z(n3452) );
  BUFFD0 U3437 ( .I(n3454), .Z(n3453) );
  BUFFD0 U3438 ( .I(n3455), .Z(n3454) );
  BUFFD0 U3439 ( .I(n3456), .Z(n3455) );
  BUFFD0 U3440 ( .I(n3457), .Z(n3456) );
  BUFFD0 U3441 ( .I(n3401), .Z(n3457) );
  BUFFD0 U3442 ( .I(n3462), .Z(n3458) );
  BUFFD0 U3443 ( .I(n4012), .Z(n3459) );
  BUFFD0 U3444 ( .I(n3459), .Z(n3460) );
  BUFFD0 U3445 ( .I(n3460), .Z(n3461) );
  BUFFD0 U3446 ( .I(n3463), .Z(n3462) );
  BUFFD0 U3447 ( .I(n3464), .Z(n3463) );
  BUFFD0 U3448 ( .I(n3465), .Z(n3464) );
  BUFFD0 U3449 ( .I(n3466), .Z(n3465) );
  BUFFD0 U3450 ( .I(n3467), .Z(n3466) );
  BUFFD0 U3451 ( .I(n3468), .Z(n3467) );
  BUFFD0 U3452 ( .I(n3469), .Z(n3468) );
  BUFFD0 U3453 ( .I(n3470), .Z(n3469) );
  BUFFD0 U3454 ( .I(n3471), .Z(n3470) );
  BUFFD0 U3455 ( .I(n3472), .Z(n3471) );
  BUFFD0 U3456 ( .I(n3473), .Z(n3472) );
  BUFFD0 U3457 ( .I(n3474), .Z(n3473) );
  BUFFD0 U3458 ( .I(n3475), .Z(n3474) );
  BUFFD0 U3459 ( .I(n3476), .Z(n3475) );
  BUFFD0 U3460 ( .I(n3477), .Z(n3476) );
  BUFFD0 U3461 ( .I(n3478), .Z(n3477) );
  BUFFD0 U3462 ( .I(n3479), .Z(n3478) );
  BUFFD0 U3463 ( .I(n3480), .Z(n3479) );
  BUFFD0 U3464 ( .I(n3481), .Z(n3480) );
  BUFFD0 U3465 ( .I(n3482), .Z(n3481) );
  BUFFD0 U3466 ( .I(n3483), .Z(n3482) );
  BUFFD0 U3467 ( .I(n3484), .Z(n3483) );
  BUFFD0 U3468 ( .I(n3485), .Z(n3484) );
  BUFFD0 U3469 ( .I(n3486), .Z(n3485) );
  BUFFD0 U3470 ( .I(n3487), .Z(n3486) );
  BUFFD0 U3471 ( .I(n3488), .Z(n3487) );
  BUFFD0 U3472 ( .I(n3489), .Z(n3488) );
  BUFFD0 U3473 ( .I(n3490), .Z(n3489) );
  BUFFD0 U3474 ( .I(n3491), .Z(n3490) );
  BUFFD0 U3475 ( .I(n3492), .Z(n3491) );
  BUFFD0 U3476 ( .I(n3493), .Z(n3492) );
  BUFFD0 U3477 ( .I(n3494), .Z(n3493) );
  BUFFD0 U3478 ( .I(n3495), .Z(n3494) );
  BUFFD0 U3479 ( .I(n3496), .Z(n3495) );
  BUFFD0 U3480 ( .I(n3497), .Z(n3496) );
  BUFFD0 U3481 ( .I(n3498), .Z(n3497) );
  BUFFD0 U3482 ( .I(n3499), .Z(n3498) );
  BUFFD0 U3483 ( .I(n3500), .Z(n3499) );
  BUFFD0 U3484 ( .I(n3501), .Z(n3500) );
  BUFFD0 U3485 ( .I(n3502), .Z(n3501) );
  BUFFD0 U3486 ( .I(n3503), .Z(n3502) );
  BUFFD0 U3487 ( .I(n3504), .Z(n3503) );
  BUFFD0 U3488 ( .I(n3505), .Z(n3504) );
  BUFFD0 U3489 ( .I(n3506), .Z(n3505) );
  BUFFD0 U3490 ( .I(n3507), .Z(n3506) );
  BUFFD0 U3491 ( .I(n3508), .Z(n3507) );
  BUFFD0 U3492 ( .I(n3509), .Z(n3508) );
  BUFFD0 U3493 ( .I(n3510), .Z(n3509) );
  BUFFD0 U3494 ( .I(n3511), .Z(n3510) );
  BUFFD0 U3495 ( .I(n3512), .Z(n3511) );
  BUFFD0 U3496 ( .I(n3513), .Z(n3512) );
  BUFFD0 U3497 ( .I(n3514), .Z(n3513) );
  BUFFD0 U3498 ( .I(n3515), .Z(n3514) );
  BUFFD0 U3499 ( .I(n3516), .Z(n3515) );
  BUFFD0 U3500 ( .I(n3461), .Z(n3516) );
  BUFFD0 U3501 ( .I(n3521), .Z(n3517) );
  BUFFD0 U3502 ( .I(N76), .Z(n3518) );
  BUFFD0 U3503 ( .I(n3518), .Z(n3519) );
  BUFFD0 U3504 ( .I(n3519), .Z(n3520) );
  BUFFD0 U3505 ( .I(n3522), .Z(n3521) );
  BUFFD0 U3506 ( .I(n3523), .Z(n3522) );
  BUFFD0 U3507 ( .I(n3524), .Z(n3523) );
  BUFFD0 U3508 ( .I(n3525), .Z(n3524) );
  BUFFD0 U3509 ( .I(n3526), .Z(n3525) );
  BUFFD0 U3510 ( .I(n3527), .Z(n3526) );
  BUFFD0 U3511 ( .I(n3528), .Z(n3527) );
  BUFFD0 U3512 ( .I(n3529), .Z(n3528) );
  BUFFD0 U3513 ( .I(n3530), .Z(n3529) );
  BUFFD0 U3514 ( .I(n3531), .Z(n3530) );
  BUFFD0 U3515 ( .I(n3532), .Z(n3531) );
  BUFFD0 U3516 ( .I(n3533), .Z(n3532) );
  BUFFD0 U3517 ( .I(n3534), .Z(n3533) );
  BUFFD0 U3518 ( .I(n3535), .Z(n3534) );
  BUFFD0 U3519 ( .I(n3536), .Z(n3535) );
  BUFFD0 U3520 ( .I(n3537), .Z(n3536) );
  BUFFD0 U3521 ( .I(n3538), .Z(n3537) );
  BUFFD0 U3522 ( .I(n3539), .Z(n3538) );
  BUFFD0 U3523 ( .I(n3540), .Z(n3539) );
  BUFFD0 U3524 ( .I(n3541), .Z(n3540) );
  BUFFD0 U3525 ( .I(n3542), .Z(n3541) );
  BUFFD0 U3526 ( .I(n3543), .Z(n3542) );
  BUFFD0 U3527 ( .I(n3544), .Z(n3543) );
  BUFFD0 U3528 ( .I(n3545), .Z(n3544) );
  BUFFD0 U3529 ( .I(n3546), .Z(n3545) );
  BUFFD0 U3530 ( .I(n3547), .Z(n3546) );
  BUFFD0 U3531 ( .I(n3548), .Z(n3547) );
  BUFFD0 U3532 ( .I(n3549), .Z(n3548) );
  BUFFD0 U3533 ( .I(n3550), .Z(n3549) );
  BUFFD0 U3534 ( .I(n3551), .Z(n3550) );
  BUFFD0 U3535 ( .I(n3552), .Z(n3551) );
  BUFFD0 U3536 ( .I(n3553), .Z(n3552) );
  BUFFD0 U3537 ( .I(n3554), .Z(n3553) );
  BUFFD0 U3538 ( .I(n3555), .Z(n3554) );
  BUFFD0 U3539 ( .I(n3556), .Z(n3555) );
  BUFFD0 U3540 ( .I(n3557), .Z(n3556) );
  BUFFD0 U3541 ( .I(n3558), .Z(n3557) );
  BUFFD0 U3542 ( .I(n3559), .Z(n3558) );
  BUFFD0 U3543 ( .I(n3560), .Z(n3559) );
  BUFFD0 U3544 ( .I(n3561), .Z(n3560) );
  BUFFD0 U3545 ( .I(n3562), .Z(n3561) );
  BUFFD0 U3546 ( .I(n3563), .Z(n3562) );
  BUFFD0 U3547 ( .I(n3564), .Z(n3563) );
  BUFFD0 U3548 ( .I(n3565), .Z(n3564) );
  BUFFD0 U3549 ( .I(n3566), .Z(n3565) );
  BUFFD0 U3550 ( .I(n3567), .Z(n3566) );
  BUFFD0 U3551 ( .I(n3568), .Z(n3567) );
  BUFFD0 U3552 ( .I(n3569), .Z(n3568) );
  BUFFD0 U3553 ( .I(n3570), .Z(n3569) );
  BUFFD0 U3554 ( .I(n3571), .Z(n3570) );
  BUFFD0 U3555 ( .I(n3572), .Z(n3571) );
  BUFFD0 U3556 ( .I(n3573), .Z(n3572) );
  BUFFD0 U3557 ( .I(n3574), .Z(n3573) );
  BUFFD0 U3558 ( .I(n3575), .Z(n3574) );
  BUFFD0 U3559 ( .I(n4015), .Z(n3575) );
  BUFFD0 U3560 ( .I(n3580), .Z(n3576) );
  BUFFD0 U3561 ( .I(N77), .Z(n3577) );
  BUFFD0 U3562 ( .I(n3577), .Z(n3578) );
  BUFFD0 U3563 ( .I(n3578), .Z(n3579) );
  BUFFD0 U3564 ( .I(n3581), .Z(n3580) );
  BUFFD0 U3565 ( .I(n3582), .Z(n3581) );
  BUFFD0 U3566 ( .I(n3583), .Z(n3582) );
  BUFFD0 U3567 ( .I(n3584), .Z(n3583) );
  BUFFD0 U3568 ( .I(n3585), .Z(n3584) );
  BUFFD0 U3569 ( .I(n3586), .Z(n3585) );
  BUFFD0 U3570 ( .I(n3587), .Z(n3586) );
  BUFFD0 U3571 ( .I(n3588), .Z(n3587) );
  BUFFD0 U3572 ( .I(n3589), .Z(n3588) );
  BUFFD0 U3573 ( .I(n3590), .Z(n3589) );
  BUFFD0 U3574 ( .I(n3591), .Z(n3590) );
  BUFFD0 U3575 ( .I(n3592), .Z(n3591) );
  BUFFD0 U3576 ( .I(n3593), .Z(n3592) );
  BUFFD0 U3577 ( .I(n3594), .Z(n3593) );
  BUFFD0 U3578 ( .I(n3595), .Z(n3594) );
  BUFFD0 U3579 ( .I(n3596), .Z(n3595) );
  BUFFD0 U3580 ( .I(n3597), .Z(n3596) );
  BUFFD0 U3581 ( .I(n3598), .Z(n3597) );
  BUFFD0 U3582 ( .I(n3599), .Z(n3598) );
  BUFFD0 U3583 ( .I(n3600), .Z(n3599) );
  BUFFD0 U3584 ( .I(n3601), .Z(n3600) );
  BUFFD0 U3585 ( .I(n3602), .Z(n3601) );
  BUFFD0 U3586 ( .I(n3603), .Z(n3602) );
  BUFFD0 U3587 ( .I(n3604), .Z(n3603) );
  BUFFD0 U3588 ( .I(n3605), .Z(n3604) );
  BUFFD0 U3589 ( .I(n3606), .Z(n3605) );
  BUFFD0 U3590 ( .I(n3607), .Z(n3606) );
  BUFFD0 U3591 ( .I(n3608), .Z(n3607) );
  BUFFD0 U3592 ( .I(n3609), .Z(n3608) );
  BUFFD0 U3593 ( .I(n3610), .Z(n3609) );
  BUFFD0 U3594 ( .I(n3611), .Z(n3610) );
  BUFFD0 U3595 ( .I(n3612), .Z(n3611) );
  BUFFD0 U3596 ( .I(n3613), .Z(n3612) );
  BUFFD0 U3597 ( .I(n3614), .Z(n3613) );
  BUFFD0 U3598 ( .I(n3615), .Z(n3614) );
  BUFFD0 U3599 ( .I(n3616), .Z(n3615) );
  BUFFD0 U3600 ( .I(n3617), .Z(n3616) );
  BUFFD0 U3601 ( .I(n3618), .Z(n3617) );
  BUFFD0 U3602 ( .I(n3619), .Z(n3618) );
  BUFFD0 U3603 ( .I(n3620), .Z(n3619) );
  BUFFD0 U3604 ( .I(n3621), .Z(n3620) );
  BUFFD0 U3605 ( .I(n3622), .Z(n3621) );
  BUFFD0 U3606 ( .I(n3623), .Z(n3622) );
  BUFFD0 U3607 ( .I(n3624), .Z(n3623) );
  BUFFD0 U3608 ( .I(n3625), .Z(n3624) );
  BUFFD0 U3609 ( .I(n3626), .Z(n3625) );
  BUFFD0 U3610 ( .I(n3627), .Z(n3626) );
  BUFFD0 U3611 ( .I(n3628), .Z(n3627) );
  BUFFD0 U3612 ( .I(n3629), .Z(n3628) );
  BUFFD0 U3613 ( .I(n3630), .Z(n3629) );
  BUFFD0 U3614 ( .I(n3631), .Z(n3630) );
  BUFFD0 U3615 ( .I(n3632), .Z(n3631) );
  BUFFD0 U3616 ( .I(n3633), .Z(n3632) );
  BUFFD0 U3617 ( .I(n3634), .Z(n3633) );
  BUFFD0 U3618 ( .I(n4008), .Z(n3634) );
  BUFFD0 U3619 ( .I(n3639), .Z(n3635) );
  BUFFD0 U3620 ( .I(N78), .Z(n3636) );
  BUFFD0 U3621 ( .I(n3636), .Z(n3637) );
  BUFFD0 U3622 ( .I(n3637), .Z(n3638) );
  BUFFD0 U3623 ( .I(n3640), .Z(n3639) );
  BUFFD0 U3624 ( .I(n3641), .Z(n3640) );
  BUFFD0 U3625 ( .I(n3642), .Z(n3641) );
  BUFFD0 U3626 ( .I(n3643), .Z(n3642) );
  BUFFD0 U3627 ( .I(n3644), .Z(n3643) );
  BUFFD0 U3628 ( .I(n3645), .Z(n3644) );
  BUFFD0 U3629 ( .I(n3646), .Z(n3645) );
  BUFFD0 U3630 ( .I(n3647), .Z(n3646) );
  BUFFD0 U3631 ( .I(n3648), .Z(n3647) );
  BUFFD0 U3632 ( .I(n3649), .Z(n3648) );
  BUFFD0 U3633 ( .I(n3650), .Z(n3649) );
  BUFFD0 U3634 ( .I(n3651), .Z(n3650) );
  BUFFD0 U3635 ( .I(n3652), .Z(n3651) );
  BUFFD0 U3636 ( .I(n3653), .Z(n3652) );
  BUFFD0 U3637 ( .I(n3654), .Z(n3653) );
  BUFFD0 U3638 ( .I(n3655), .Z(n3654) );
  BUFFD0 U3639 ( .I(n3656), .Z(n3655) );
  BUFFD0 U3640 ( .I(n3657), .Z(n3656) );
  BUFFD0 U3641 ( .I(n3658), .Z(n3657) );
  BUFFD0 U3642 ( .I(n3659), .Z(n3658) );
  BUFFD0 U3643 ( .I(n3660), .Z(n3659) );
  BUFFD0 U3644 ( .I(n3661), .Z(n3660) );
  BUFFD0 U3645 ( .I(n3662), .Z(n3661) );
  BUFFD0 U3646 ( .I(n3663), .Z(n3662) );
  BUFFD0 U3647 ( .I(n3664), .Z(n3663) );
  BUFFD0 U3648 ( .I(n3665), .Z(n3664) );
  BUFFD0 U3649 ( .I(n3666), .Z(n3665) );
  BUFFD0 U3650 ( .I(n3667), .Z(n3666) );
  BUFFD0 U3651 ( .I(n3668), .Z(n3667) );
  BUFFD0 U3652 ( .I(n3669), .Z(n3668) );
  BUFFD0 U3653 ( .I(n3670), .Z(n3669) );
  BUFFD0 U3654 ( .I(n3671), .Z(n3670) );
  BUFFD0 U3655 ( .I(n3672), .Z(n3671) );
  BUFFD0 U3656 ( .I(n3673), .Z(n3672) );
  BUFFD0 U3657 ( .I(n3674), .Z(n3673) );
  BUFFD0 U3658 ( .I(n3675), .Z(n3674) );
  BUFFD0 U3659 ( .I(n3676), .Z(n3675) );
  BUFFD0 U3660 ( .I(n3677), .Z(n3676) );
  BUFFD0 U3661 ( .I(n3678), .Z(n3677) );
  BUFFD0 U3662 ( .I(n3679), .Z(n3678) );
  BUFFD0 U3663 ( .I(n3680), .Z(n3679) );
  BUFFD0 U3664 ( .I(n3681), .Z(n3680) );
  BUFFD0 U3665 ( .I(n3682), .Z(n3681) );
  BUFFD0 U3666 ( .I(n3683), .Z(n3682) );
  BUFFD0 U3667 ( .I(n3684), .Z(n3683) );
  BUFFD0 U3668 ( .I(n3685), .Z(n3684) );
  BUFFD0 U3669 ( .I(n3686), .Z(n3685) );
  BUFFD0 U3670 ( .I(n3687), .Z(n3686) );
  BUFFD0 U3671 ( .I(n3688), .Z(n3687) );
  BUFFD0 U3672 ( .I(n3689), .Z(n3688) );
  BUFFD0 U3673 ( .I(n3690), .Z(n3689) );
  BUFFD0 U3674 ( .I(n4038), .Z(n3690) );
  BUFFD0 U3675 ( .I(n3695), .Z(n3691) );
  BUFFD0 U3676 ( .I(n4006), .Z(n3692) );
  BUFFD0 U3677 ( .I(n3692), .Z(n3693) );
  BUFFD0 U3678 ( .I(n3693), .Z(n3694) );
  BUFFD0 U3679 ( .I(n3696), .Z(n3695) );
  BUFFD0 U3680 ( .I(n3697), .Z(n3696) );
  BUFFD0 U3681 ( .I(n3698), .Z(n3697) );
  BUFFD0 U3682 ( .I(n3699), .Z(n3698) );
  BUFFD0 U3683 ( .I(n3700), .Z(n3699) );
  BUFFD0 U3684 ( .I(n3701), .Z(n3700) );
  BUFFD0 U3685 ( .I(n3702), .Z(n3701) );
  BUFFD0 U3686 ( .I(n3703), .Z(n3702) );
  BUFFD0 U3687 ( .I(n3704), .Z(n3703) );
  BUFFD0 U3688 ( .I(n3705), .Z(n3704) );
  BUFFD0 U3689 ( .I(n3706), .Z(n3705) );
  BUFFD0 U3690 ( .I(n3707), .Z(n3706) );
  BUFFD0 U3691 ( .I(n3708), .Z(n3707) );
  BUFFD0 U3692 ( .I(n3709), .Z(n3708) );
  BUFFD0 U3693 ( .I(n3710), .Z(n3709) );
  BUFFD0 U3694 ( .I(n3711), .Z(n3710) );
  BUFFD0 U3695 ( .I(n3712), .Z(n3711) );
  BUFFD0 U3696 ( .I(n3713), .Z(n3712) );
  BUFFD0 U3697 ( .I(n3714), .Z(n3713) );
  BUFFD0 U3698 ( .I(n3715), .Z(n3714) );
  BUFFD0 U3699 ( .I(n3716), .Z(n3715) );
  BUFFD0 U3700 ( .I(n3717), .Z(n3716) );
  BUFFD0 U3701 ( .I(n3718), .Z(n3717) );
  BUFFD0 U3702 ( .I(n3719), .Z(n3718) );
  BUFFD0 U3703 ( .I(n3720), .Z(n3719) );
  BUFFD0 U3704 ( .I(n3721), .Z(n3720) );
  BUFFD0 U3705 ( .I(n3722), .Z(n3721) );
  BUFFD0 U3706 ( .I(n3723), .Z(n3722) );
  BUFFD0 U3707 ( .I(n3724), .Z(n3723) );
  BUFFD0 U3708 ( .I(n3725), .Z(n3724) );
  BUFFD0 U3709 ( .I(n3726), .Z(n3725) );
  BUFFD0 U3710 ( .I(n3727), .Z(n3726) );
  BUFFD0 U3711 ( .I(n3728), .Z(n3727) );
  BUFFD0 U3712 ( .I(n3729), .Z(n3728) );
  BUFFD0 U3713 ( .I(n3730), .Z(n3729) );
  BUFFD0 U3714 ( .I(n3731), .Z(n3730) );
  BUFFD0 U3715 ( .I(n3732), .Z(n3731) );
  BUFFD0 U3716 ( .I(n3733), .Z(n3732) );
  BUFFD0 U3717 ( .I(n3734), .Z(n3733) );
  BUFFD0 U3718 ( .I(n3735), .Z(n3734) );
  BUFFD0 U3719 ( .I(n3736), .Z(n3735) );
  BUFFD0 U3720 ( .I(n3737), .Z(n3736) );
  BUFFD0 U3721 ( .I(n3738), .Z(n3737) );
  BUFFD0 U3722 ( .I(n3739), .Z(n3738) );
  BUFFD0 U3723 ( .I(n3740), .Z(n3739) );
  BUFFD0 U3724 ( .I(n3741), .Z(n3740) );
  BUFFD0 U3725 ( .I(n3742), .Z(n3741) );
  BUFFD0 U3726 ( .I(n3743), .Z(n3742) );
  BUFFD0 U3727 ( .I(n3744), .Z(n3743) );
  BUFFD0 U3728 ( .I(n3745), .Z(n3744) );
  BUFFD0 U3729 ( .I(n3746), .Z(n3745) );
  BUFFD0 U3730 ( .I(n3747), .Z(n3746) );
  BUFFD0 U3731 ( .I(n3748), .Z(n3747) );
  BUFFD0 U3732 ( .I(n3749), .Z(n3748) );
  BUFFD0 U3733 ( .I(n3694), .Z(n3749) );
  BUFFD0 U3734 ( .I(n3754), .Z(n3750) );
  BUFFD0 U3735 ( .I(n4004), .Z(n3751) );
  BUFFD0 U3736 ( .I(n3751), .Z(n3752) );
  BUFFD0 U3737 ( .I(n3752), .Z(n3753) );
  BUFFD0 U3738 ( .I(n3755), .Z(n3754) );
  BUFFD0 U3739 ( .I(n3756), .Z(n3755) );
  BUFFD0 U3740 ( .I(n3757), .Z(n3756) );
  BUFFD0 U3741 ( .I(n3758), .Z(n3757) );
  BUFFD0 U3742 ( .I(n3759), .Z(n3758) );
  BUFFD0 U3743 ( .I(n3760), .Z(n3759) );
  BUFFD0 U3744 ( .I(n3761), .Z(n3760) );
  BUFFD0 U3745 ( .I(n3762), .Z(n3761) );
  BUFFD0 U3746 ( .I(n3763), .Z(n3762) );
  BUFFD0 U3747 ( .I(n3764), .Z(n3763) );
  BUFFD0 U3748 ( .I(n3765), .Z(n3764) );
  BUFFD0 U3749 ( .I(n3766), .Z(n3765) );
  BUFFD0 U3750 ( .I(n3767), .Z(n3766) );
  BUFFD0 U3751 ( .I(n3768), .Z(n3767) );
  BUFFD0 U3752 ( .I(n3769), .Z(n3768) );
  BUFFD0 U3753 ( .I(n3770), .Z(n3769) );
  BUFFD0 U3754 ( .I(n3771), .Z(n3770) );
  BUFFD0 U3755 ( .I(n3772), .Z(n3771) );
  BUFFD0 U3756 ( .I(n3773), .Z(n3772) );
  BUFFD0 U3757 ( .I(n3774), .Z(n3773) );
  BUFFD0 U3758 ( .I(n3775), .Z(n3774) );
  BUFFD0 U3759 ( .I(n3776), .Z(n3775) );
  BUFFD0 U3760 ( .I(n3777), .Z(n3776) );
  BUFFD0 U3761 ( .I(n3778), .Z(n3777) );
  BUFFD0 U3762 ( .I(n3779), .Z(n3778) );
  BUFFD0 U3763 ( .I(n3780), .Z(n3779) );
  BUFFD0 U3764 ( .I(n3781), .Z(n3780) );
  BUFFD0 U3765 ( .I(n3782), .Z(n3781) );
  BUFFD0 U3766 ( .I(n3783), .Z(n3782) );
  BUFFD0 U3767 ( .I(n3784), .Z(n3783) );
  BUFFD0 U3768 ( .I(n3785), .Z(n3784) );
  BUFFD0 U3769 ( .I(n3786), .Z(n3785) );
  BUFFD0 U3770 ( .I(n3787), .Z(n3786) );
  BUFFD0 U3771 ( .I(n3788), .Z(n3787) );
  BUFFD0 U3772 ( .I(n3789), .Z(n3788) );
  BUFFD0 U3773 ( .I(n3790), .Z(n3789) );
  BUFFD0 U3774 ( .I(n3791), .Z(n3790) );
  BUFFD0 U3775 ( .I(n3792), .Z(n3791) );
  BUFFD0 U3776 ( .I(n3793), .Z(n3792) );
  BUFFD0 U3777 ( .I(n3794), .Z(n3793) );
  BUFFD0 U3778 ( .I(n3795), .Z(n3794) );
  BUFFD0 U3779 ( .I(n3796), .Z(n3795) );
  BUFFD0 U3780 ( .I(n3797), .Z(n3796) );
  BUFFD0 U3781 ( .I(n3798), .Z(n3797) );
  BUFFD0 U3782 ( .I(n3799), .Z(n3798) );
  BUFFD0 U3783 ( .I(n3800), .Z(n3799) );
  BUFFD0 U3784 ( .I(n3801), .Z(n3800) );
  BUFFD0 U3785 ( .I(n3802), .Z(n3801) );
  BUFFD0 U3786 ( .I(n3803), .Z(n3802) );
  BUFFD0 U3787 ( .I(n3804), .Z(n3803) );
  BUFFD0 U3788 ( .I(n3805), .Z(n3804) );
  BUFFD0 U3789 ( .I(n3806), .Z(n3805) );
  BUFFD0 U3790 ( .I(n3807), .Z(n3806) );
  BUFFD0 U3791 ( .I(n3808), .Z(n3807) );
  BUFFD0 U3792 ( .I(n3753), .Z(n3808) );
  BUFFD0 U3793 ( .I(n3813), .Z(n3809) );
  BUFFD0 U3794 ( .I(N81), .Z(n3810) );
  BUFFD0 U3795 ( .I(n3810), .Z(n3811) );
  BUFFD0 U3796 ( .I(n3811), .Z(n3812) );
  BUFFD0 U3797 ( .I(n3814), .Z(n3813) );
  BUFFD0 U3798 ( .I(n3815), .Z(n3814) );
  BUFFD0 U3799 ( .I(n3816), .Z(n3815) );
  BUFFD0 U3800 ( .I(n3817), .Z(n3816) );
  BUFFD0 U3801 ( .I(n3818), .Z(n3817) );
  BUFFD0 U3802 ( .I(n3819), .Z(n3818) );
  BUFFD0 U3803 ( .I(n3820), .Z(n3819) );
  BUFFD0 U3804 ( .I(n3821), .Z(n3820) );
  BUFFD0 U3805 ( .I(n3822), .Z(n3821) );
  BUFFD0 U3806 ( .I(n3823), .Z(n3822) );
  BUFFD0 U3807 ( .I(n3824), .Z(n3823) );
  BUFFD0 U3808 ( .I(n3825), .Z(n3824) );
  BUFFD0 U3809 ( .I(n3826), .Z(n3825) );
  BUFFD0 U3810 ( .I(n3827), .Z(n3826) );
  BUFFD0 U3811 ( .I(n3828), .Z(n3827) );
  BUFFD0 U3812 ( .I(n3829), .Z(n3828) );
  BUFFD0 U3813 ( .I(n3830), .Z(n3829) );
  BUFFD0 U3814 ( .I(n3831), .Z(n3830) );
  BUFFD0 U3815 ( .I(n3832), .Z(n3831) );
  BUFFD0 U3816 ( .I(n3833), .Z(n3832) );
  BUFFD0 U3817 ( .I(n3834), .Z(n3833) );
  BUFFD0 U3818 ( .I(n3835), .Z(n3834) );
  BUFFD0 U3819 ( .I(n3836), .Z(n3835) );
  BUFFD0 U3820 ( .I(n3837), .Z(n3836) );
  BUFFD0 U3821 ( .I(n3838), .Z(n3837) );
  BUFFD0 U3822 ( .I(n3839), .Z(n3838) );
  BUFFD0 U3823 ( .I(n3840), .Z(n3839) );
  BUFFD0 U3824 ( .I(n3841), .Z(n3840) );
  BUFFD0 U3825 ( .I(n3842), .Z(n3841) );
  BUFFD0 U3826 ( .I(n3843), .Z(n3842) );
  BUFFD0 U3827 ( .I(n3844), .Z(n3843) );
  BUFFD0 U3828 ( .I(n3845), .Z(n3844) );
  BUFFD0 U3829 ( .I(n3846), .Z(n3845) );
  BUFFD0 U3830 ( .I(n3847), .Z(n3846) );
  BUFFD0 U3831 ( .I(n3848), .Z(n3847) );
  BUFFD0 U3832 ( .I(n3849), .Z(n3848) );
  BUFFD0 U3833 ( .I(n3850), .Z(n3849) );
  BUFFD0 U3834 ( .I(n3851), .Z(n3850) );
  BUFFD0 U3835 ( .I(n3852), .Z(n3851) );
  BUFFD0 U3836 ( .I(n3853), .Z(n3852) );
  BUFFD0 U3837 ( .I(n3854), .Z(n3853) );
  BUFFD0 U3838 ( .I(n3855), .Z(n3854) );
  BUFFD0 U3839 ( .I(n3856), .Z(n3855) );
  BUFFD0 U3840 ( .I(n3857), .Z(n3856) );
  BUFFD0 U3841 ( .I(n3858), .Z(n3857) );
  BUFFD0 U3842 ( .I(n3859), .Z(n3858) );
  BUFFD0 U3843 ( .I(n3860), .Z(n3859) );
  BUFFD0 U3844 ( .I(n3861), .Z(n3860) );
  BUFFD0 U3845 ( .I(n3862), .Z(n3861) );
  BUFFD0 U3846 ( .I(n3863), .Z(n3862) );
  BUFFD0 U3847 ( .I(n3864), .Z(n3863) );
  BUFFD0 U3848 ( .I(n3865), .Z(n3864) );
  BUFFD0 U3849 ( .I(n3866), .Z(n3865) );
  BUFFD0 U3850 ( .I(n3867), .Z(n3866) );
  BUFFD0 U3851 ( .I(n4007), .Z(n3867) );
  BUFFD0 U3852 ( .I(N75), .Z(n3868) );
  BUFFD0 U3853 ( .I(N68), .Z(n3869) );
  BUFFD0 U3854 ( .I(N74), .Z(n3870) );
  BUFFD0 U3855 ( .I(N82), .Z(n3871) );
  BUFFD0 U3856 ( .I(n3871), .Z(n3872) );
  BUFFD0 U3857 ( .I(n3874), .Z(n3873) );
  BUFFD0 U3858 ( .I(n3875), .Z(n3874) );
  BUFFD0 U3859 ( .I(n3876), .Z(n3875) );
  BUFFD0 U3860 ( .I(n3877), .Z(n3876) );
  BUFFD0 U3861 ( .I(n3878), .Z(n3877) );
  BUFFD0 U3862 ( .I(n3879), .Z(n3878) );
  BUFFD0 U3863 ( .I(n3880), .Z(n3879) );
  BUFFD0 U3864 ( .I(n3881), .Z(n3880) );
  BUFFD0 U3865 ( .I(n3882), .Z(n3881) );
  BUFFD0 U3866 ( .I(n3883), .Z(n3882) );
  BUFFD0 U3867 ( .I(n3884), .Z(n3883) );
  BUFFD0 U3868 ( .I(n3885), .Z(n3884) );
  BUFFD0 U3869 ( .I(n3886), .Z(n3885) );
  BUFFD0 U3870 ( .I(n3887), .Z(n3886) );
  BUFFD0 U3871 ( .I(n3888), .Z(n3887) );
  BUFFD0 U3872 ( .I(n3889), .Z(n3888) );
  BUFFD0 U3873 ( .I(n3890), .Z(n3889) );
  BUFFD0 U3874 ( .I(n3891), .Z(n3890) );
  BUFFD0 U3875 ( .I(n3892), .Z(n3891) );
  BUFFD0 U3876 ( .I(n3893), .Z(n3892) );
  BUFFD0 U3877 ( .I(n3894), .Z(n3893) );
  BUFFD0 U3878 ( .I(n3895), .Z(n3894) );
  BUFFD0 U3879 ( .I(n3896), .Z(n3895) );
  BUFFD0 U3880 ( .I(n3897), .Z(n3896) );
  BUFFD0 U3881 ( .I(n3898), .Z(n3897) );
  BUFFD0 U3882 ( .I(n3899), .Z(n3898) );
  BUFFD0 U3883 ( .I(n3900), .Z(n3899) );
  BUFFD0 U3884 ( .I(n3901), .Z(n3900) );
  BUFFD0 U3885 ( .I(n3902), .Z(n3901) );
  BUFFD0 U3886 ( .I(n3903), .Z(n3902) );
  BUFFD0 U3887 ( .I(n3904), .Z(n3903) );
  BUFFD0 U3888 ( .I(n3905), .Z(n3904) );
  BUFFD0 U3889 ( .I(n3906), .Z(n3905) );
  BUFFD0 U3890 ( .I(n3907), .Z(n3906) );
  BUFFD0 U3891 ( .I(n3908), .Z(n3907) );
  BUFFD0 U3892 ( .I(n3909), .Z(n3908) );
  BUFFD0 U3893 ( .I(n3910), .Z(n3909) );
  BUFFD0 U3894 ( .I(n3911), .Z(n3910) );
  BUFFD0 U3895 ( .I(n3912), .Z(n3911) );
  BUFFD0 U3896 ( .I(n3913), .Z(n3912) );
  BUFFD0 U3897 ( .I(n3914), .Z(n3913) );
  BUFFD0 U3898 ( .I(n3915), .Z(n3914) );
  BUFFD0 U3899 ( .I(n3916), .Z(n3915) );
  BUFFD0 U3900 ( .I(n3917), .Z(n3916) );
  BUFFD0 U3901 ( .I(n3918), .Z(n3917) );
  BUFFD0 U3902 ( .I(n3919), .Z(n3918) );
  BUFFD0 U3903 ( .I(n3920), .Z(n3919) );
  BUFFD0 U3904 ( .I(n3921), .Z(n3920) );
  BUFFD0 U3905 ( .I(n3922), .Z(n3921) );
  BUFFD0 U3906 ( .I(n3923), .Z(n3922) );
  BUFFD0 U3907 ( .I(n3951), .Z(n3923) );
  BUFFD0 U3908 ( .I(n2650), .Z(n3924) );
  BUFFD0 U3909 ( .I(n3948), .Z(n3925) );
  BUFFD0 U3910 ( .I(n3520), .Z(n3926) );
  BUFFD0 U3911 ( .I(N80), .Z(n3927) );
  BUFFD0 U3912 ( .I(N79), .Z(n3928) );
  BUFFD0 U3913 ( .I(n2975), .Z(n3929) );
  BUFFD0 U3914 ( .I(n3812), .Z(n3930) );
  BUFFD0 U3915 ( .I(n2716), .Z(n3931) );
  BUFFD0 U3916 ( .I(n2584), .Z(n3932) );
  BUFFD0 U3917 ( .I(n3955), .Z(n3933) );
  BUFFD0 U3918 ( .I(N65), .Z(n3934) );
  BUFFD0 U3919 ( .I(n2782), .Z(n3935) );
  BUFFD0 U3920 ( .I(n3579), .Z(n3936) );
  BUFFD0 U3921 ( .I(n3286), .Z(n3937) );
  BUFFD0 U3922 ( .I(N73), .Z(n3938) );
  BUFFD0 U3923 ( .I(n2971), .Z(n3939) );
  BUFFD0 U3924 ( .I(N69), .Z(n3940) );
  BUFFD0 U3925 ( .I(n3638), .Z(n3941) );
  BUFFD0 U3926 ( .I(n3221), .Z(n3942) );
  BUFFD0 U3927 ( .I(n2453), .Z(n3943) );
  BUFFD0 U3928 ( .I(n3868), .Z(n3944) );
  BUFFD0 U3929 ( .I(n3869), .Z(n3945) );
  BUFFD0 U3930 ( .I(n3225), .Z(n3946) );
  BUFFD0 U3931 ( .I(n3870), .Z(n3947) );
  BUFFD0 U3932 ( .I(n2518), .Z(n3948) );
  BUFFD0 U3933 ( .I(n3926), .Z(n3949) );
  BUFFD0 U3934 ( .I(n3927), .Z(n3950) );
  BUFFD0 U3935 ( .I(n3872), .Z(n3951) );
  BUFFD0 U3936 ( .I(n3928), .Z(n3952) );
  BUFFD0 U3937 ( .I(n3929), .Z(n3953) );
  BUFFD0 U3938 ( .I(n3930), .Z(n3954) );
  BUFFD0 U3939 ( .I(n3973), .Z(n3955) );
  BUFFD0 U3940 ( .I(n3974), .Z(n3956) );
  BUFFD0 U3941 ( .I(n3936), .Z(n3957) );
  BUFFD0 U3942 ( .I(n3937), .Z(n3958) );
  BUFFD0 U3943 ( .I(n3938), .Z(n3959) );
  BUFFD0 U3944 ( .I(n3978), .Z(n3960) );
  BUFFD0 U3945 ( .I(n3979), .Z(n3961) );
  BUFFD0 U3946 ( .I(n3941), .Z(n3962) );
  BUFFD0 U3947 ( .I(n3981), .Z(n3963) );
  BUFFD0 U3948 ( .I(n3944), .Z(n3964) );
  BUFFD0 U3949 ( .I(n3983), .Z(n3965) );
  BUFFD0 U3950 ( .I(n3947), .Z(n3966) );
  BUFFD0 U3951 ( .I(n3946), .Z(n3967) );
  BUFFD0 U3952 ( .I(n3949), .Z(n3968) );
  BUFFD0 U3953 ( .I(n3950), .Z(n3969) );
  BUFFD0 U3954 ( .I(n3952), .Z(n3970) );
  BUFFD0 U3955 ( .I(n3989), .Z(n3971) );
  BUFFD0 U3956 ( .I(n3954), .Z(n3972) );
  BUFFD0 U3957 ( .I(N64), .Z(n3973) );
  BUFFD0 U3958 ( .I(n3991), .Z(n3974) );
  BUFFD0 U3959 ( .I(n3957), .Z(n3975) );
  BUFFD0 U3960 ( .I(n3958), .Z(n3976) );
  BUFFD0 U3961 ( .I(n3959), .Z(n3977) );
  BUFFD0 U3962 ( .I(n3995), .Z(n3978) );
  BUFFD0 U3963 ( .I(n3996), .Z(n3979) );
  BUFFD0 U3964 ( .I(n3962), .Z(n3980) );
  BUFFD0 U3965 ( .I(n3998), .Z(n3981) );
  BUFFD0 U3966 ( .I(n3964), .Z(n3982) );
  BUFFD0 U3967 ( .I(n3999), .Z(n3983) );
  BUFFD0 U3968 ( .I(n3966), .Z(n3984) );
  BUFFD0 U3969 ( .I(n3967), .Z(n3985) );
  BUFFD0 U3970 ( .I(n3968), .Z(n3986) );
  BUFFD0 U3971 ( .I(n3969), .Z(n3987) );
  BUFFD0 U3972 ( .I(n3970), .Z(n3988) );
  BUFFD0 U3973 ( .I(n4005), .Z(n3989) );
  BUFFD0 U3974 ( .I(n3972), .Z(n3990) );
  BUFFD0 U3975 ( .I(n3934), .Z(n3991) );
  BUFFD0 U3976 ( .I(n3975), .Z(n3992) );
  BUFFD0 U3977 ( .I(n3976), .Z(n3993) );
  BUFFD0 U3978 ( .I(n3977), .Z(n3994) );
  BUFFD0 U3979 ( .I(n3939), .Z(n3995) );
  BUFFD0 U3980 ( .I(n3940), .Z(n3996) );
  BUFFD0 U3981 ( .I(n3980), .Z(n3997) );
  BUFFD0 U3982 ( .I(n3942), .Z(n3998) );
  BUFFD0 U3983 ( .I(n3945), .Z(n3999) );
  BUFFD0 U3984 ( .I(n3982), .Z(n4000) );
  BUFFD0 U3985 ( .I(n4013), .Z(n4001) );
  BUFFD0 U3986 ( .I(n4014), .Z(n4002) );
  BUFFD0 U3987 ( .I(n3986), .Z(n4003) );
  BUFFD0 U3988 ( .I(n4016), .Z(n4004) );
  BUFFD0 U3989 ( .I(n3953), .Z(n4005) );
  BUFFD0 U3990 ( .I(n4017), .Z(n4006) );
  BUFFD0 U3991 ( .I(n4018), .Z(n4007) );
  BUFFD0 U3992 ( .I(n4019), .Z(n4008) );
  BUFFD0 U3993 ( .I(n3993), .Z(n4009) );
  BUFFD0 U3994 ( .I(n3994), .Z(n4010) );
  BUFFD0 U3995 ( .I(n3997), .Z(n4011) );
  BUFFD0 U3996 ( .I(n4024), .Z(n4012) );
  BUFFD0 U3997 ( .I(n4023), .Z(n4013) );
  BUFFD0 U3998 ( .I(n4025), .Z(n4014) );
  BUFFD0 U3999 ( .I(n4028), .Z(n4015) );
  BUFFD0 U4000 ( .I(n4029), .Z(n4018) );
  BUFFD0 U4001 ( .I(n4030), .Z(n4019) );
  BUFFD0 U4002 ( .I(n4009), .Z(n4020) );
  BUFFD0 U4003 ( .I(n4010), .Z(n4021) );
  BUFFD0 U4004 ( .I(n4011), .Z(n4022) );
  BUFFD0 U4005 ( .I(n3984), .Z(n4023) );
  BUFFD0 U4006 ( .I(n4034), .Z(n4024) );
  BUFFD0 U4007 ( .I(n3985), .Z(n4025) );
  BUFFD0 U4008 ( .I(n3987), .Z(n4026) );
  BUFFD0 U4009 ( .I(n3988), .Z(n4027) );
  BUFFD0 U4010 ( .I(n4035), .Z(n4028) );
  BUFFD0 U4011 ( .I(n3990), .Z(n4029) );
  BUFFD0 U4012 ( .I(n3992), .Z(n4030) );
  BUFFD0 U4013 ( .I(n4036), .Z(n4031) );
  BUFFD0 U4014 ( .I(n4021), .Z(n4032) );
  BUFFD0 U4015 ( .I(n4022), .Z(n4033) );
  BUFFD0 U4016 ( .I(n4000), .Z(n4034) );
  BUFFD0 U4017 ( .I(n4003), .Z(n4035) );
  BUFFD0 U4018 ( .I(n4039), .Z(n4036) );
  BUFFD0 U4019 ( .I(n4040), .Z(n4037) );
  BUFFD0 U4020 ( .I(n4041), .Z(n4038) );
  BUFFD0 U4021 ( .I(n4020), .Z(n4039) );
  BUFFD0 U4022 ( .I(n4042), .Z(n4040) );
  BUFFD0 U4023 ( .I(n4043), .Z(n4041) );
  BUFFD0 U4024 ( .I(n4032), .Z(n4042) );
  BUFFD0 U4025 ( .I(n4033), .Z(n4043) );
  BUFFD0 U4026 ( .I(n4330), .Z(n4044) );
  BUFFD0 U4027 ( .I(n4046), .Z(n4045) );
  BUFFD0 U4028 ( .I(n4047), .Z(n4046) );
  BUFFD0 U4029 ( .I(n4048), .Z(n4047) );
  BUFFD0 U4030 ( .I(n4049), .Z(n4048) );
  BUFFD0 U4031 ( .I(n4050), .Z(n4049) );
  BUFFD0 U4032 ( .I(n4051), .Z(n4050) );
  BUFFD0 U4033 ( .I(n4052), .Z(n4051) );
  BUFFD0 U4034 ( .I(n4053), .Z(n4052) );
  BUFFD0 U4035 ( .I(n4054), .Z(n4053) );
  BUFFD0 U4036 ( .I(n4055), .Z(n4054) );
  BUFFD0 U4037 ( .I(n4056), .Z(n4055) );
  BUFFD0 U4038 ( .I(n4057), .Z(n4056) );
  BUFFD0 U4039 ( .I(n4058), .Z(n4057) );
  BUFFD0 U4040 ( .I(n4059), .Z(n4058) );
  BUFFD0 U4041 ( .I(n4060), .Z(n4059) );
  BUFFD0 U4042 ( .I(n4061), .Z(n4060) );
  BUFFD0 U4043 ( .I(n4062), .Z(n4061) );
  BUFFD0 U4044 ( .I(n4063), .Z(n4062) );
  BUFFD0 U4045 ( .I(n4064), .Z(n4063) );
  BUFFD0 U4046 ( .I(n4065), .Z(n4064) );
  BUFFD0 U4047 ( .I(n4066), .Z(n4065) );
  BUFFD0 U4048 ( .I(n4067), .Z(n4066) );
  BUFFD0 U4049 ( .I(n4068), .Z(n4067) );
  BUFFD0 U4050 ( .I(n4069), .Z(n4068) );
  BUFFD0 U4051 ( .I(n4070), .Z(n4069) );
  BUFFD0 U4052 ( .I(n4071), .Z(n4070) );
  BUFFD0 U4053 ( .I(n4072), .Z(n4071) );
  BUFFD0 U4054 ( .I(n4073), .Z(n4072) );
  BUFFD0 U4055 ( .I(n4074), .Z(n4073) );
  BUFFD0 U4056 ( .I(n4075), .Z(n4074) );
  BUFFD0 U4057 ( .I(n4076), .Z(n4075) );
  BUFFD0 U4058 ( .I(n4077), .Z(n4076) );
  BUFFD0 U4059 ( .I(n4078), .Z(n4077) );
  BUFFD0 U4060 ( .I(n4079), .Z(n4078) );
  BUFFD0 U4061 ( .I(n4080), .Z(n4079) );
  BUFFD0 U4062 ( .I(n4081), .Z(n4080) );
  BUFFD0 U4063 ( .I(n4082), .Z(n4081) );
  BUFFD0 U4064 ( .I(n4083), .Z(n4082) );
  BUFFD0 U4065 ( .I(n4084), .Z(n4083) );
  BUFFD0 U4066 ( .I(n4085), .Z(n4084) );
  BUFFD0 U4067 ( .I(n4086), .Z(n4085) );
  BUFFD0 U4068 ( .I(n4087), .Z(n4086) );
  BUFFD0 U4069 ( .I(n4088), .Z(n4087) );
  BUFFD0 U4070 ( .I(n4089), .Z(n4088) );
  BUFFD0 U4071 ( .I(n4090), .Z(n4089) );
  BUFFD0 U4072 ( .I(n4091), .Z(n4090) );
  BUFFD0 U4073 ( .I(n4092), .Z(n4091) );
  BUFFD0 U4074 ( .I(n4093), .Z(n4092) );
  BUFFD0 U4075 ( .I(n4094), .Z(n4093) );
  BUFFD0 U4076 ( .I(n4095), .Z(n4094) );
  BUFFD0 U4077 ( .I(n4096), .Z(n4095) );
  BUFFD0 U4078 ( .I(n4097), .Z(n4096) );
  BUFFD0 U4079 ( .I(n4098), .Z(n4097) );
  BUFFD0 U4080 ( .I(Read), .Z(n4098) );
  CKAN2D0 U4081 ( .A1(Dreadyr), .A2(ChipEna), .Z(Dready) );
  BUFFD1 U4082 ( .I(n4354), .Z(n4340) );
  BUFFD1 U4083 ( .I(n4354), .Z(n4341) );
  BUFFD1 U4084 ( .I(n4353), .Z(n4342) );
  BUFFD1 U4085 ( .I(n4359), .Z(n4343) );
  BUFFD1 U4086 ( .I(n4352), .Z(n4344) );
  BUFFD1 U4087 ( .I(n4352), .Z(n4345) );
  BUFFD1 U4088 ( .I(n4351), .Z(n4346) );
  BUFFD1 U4089 ( .I(n4351), .Z(n4347) );
  BUFFD1 U4090 ( .I(n4350), .Z(n4348) );
  BUFFD1 U4091 ( .I(n4350), .Z(n4349) );
  BUFFD1 U4092 ( .I(n4357), .Z(n4334) );
  BUFFD1 U4093 ( .I(n4357), .Z(n4335) );
  BUFFD1 U4094 ( .I(n4356), .Z(n4336) );
  BUFFD1 U4095 ( .I(n4356), .Z(n4337) );
  BUFFD1 U4096 ( .I(n4355), .Z(n4338) );
  BUFFD1 U4097 ( .I(n4355), .Z(n4339) );
  BUFFD1 U4098 ( .I(n4359), .Z(n4354) );
  BUFFD1 U4099 ( .I(n4359), .Z(n4353) );
  BUFFD1 U4100 ( .I(n4360), .Z(n4352) );
  BUFFD1 U4101 ( .I(n4360), .Z(n4351) );
  BUFFD1 U4102 ( .I(n4360), .Z(n4350) );
  BUFFD1 U4103 ( .I(n4358), .Z(n4356) );
  BUFFD1 U4104 ( .I(n4358), .Z(n4355) );
  BUFFD1 U4105 ( .I(n4358), .Z(n4357) );
  BUFFD1 U4106 ( .I(n4361), .Z(n4359) );
  BUFFD1 U4107 ( .I(n4361), .Z(n4360) );
  BUFFD1 U4108 ( .I(n4363), .Z(n4361) );
  BUFFD1 U4109 ( .I(n4362), .Z(n4358) );
  BUFFD1 U4110 ( .I(n4363), .Z(n4362) );
  INVD1 U4111 ( .I(Reset), .ZN(n4363) );
  BUFFD1 U4112 ( .I(n4319), .Z(n4307) );
  BUFFD1 U4113 ( .I(n4308), .Z(n4306) );
  BUFFD1 U4114 ( .I(n4308), .Z(n4305) );
  BUFFD1 U4115 ( .I(n4309), .Z(n4304) );
  BUFFD1 U4116 ( .I(n4309), .Z(n4303) );
  BUFFD1 U4117 ( .I(n4310), .Z(n4302) );
  BUFFD1 U4118 ( .I(n4311), .Z(n4301) );
  BUFFD1 U4119 ( .I(n4311), .Z(n4300) );
  BUFFD1 U4120 ( .I(n4312), .Z(n4299) );
  BUFFD1 U4121 ( .I(n4312), .Z(n4298) );
  BUFFD1 U4122 ( .I(n4313), .Z(n4297) );
  BUFFD1 U4123 ( .I(n4313), .Z(n4296) );
  BUFFD1 U4124 ( .I(n4314), .Z(n4295) );
  BUFFD1 U4125 ( .I(n4314), .Z(n4294) );
  BUFFD1 U4126 ( .I(n4315), .Z(n4293) );
  BUFFD1 U4127 ( .I(n4315), .Z(n4292) );
  BUFFD1 U4128 ( .I(n4316), .Z(n4291) );
  BUFFD1 U4129 ( .I(n4316), .Z(n4290) );
  BUFFD1 U4130 ( .I(n4317), .Z(n4289) );
  BUFFD1 U4131 ( .I(n4317), .Z(n4288) );
  BUFFD1 U4132 ( .I(n4318), .Z(n4287) );
  BUFFD1 U4133 ( .I(n4318), .Z(n4286) );
  BUFFD1 U4134 ( .I(n4319), .Z(n4285) );
  BUFFD1 U4135 ( .I(n4319), .Z(n4284) );
  BUFFD1 U4136 ( .I(n4320), .Z(n4283) );
  BUFFD1 U4137 ( .I(n4320), .Z(n4282) );
  INVD1 U4138 ( .I(n16), .ZN(n4277) );
  INVD1 U4139 ( .I(n16), .ZN(n4276) );
  INVD1 U4140 ( .I(n18), .ZN(n4261) );
  INVD1 U4141 ( .I(n18), .ZN(n4260) );
  BUFFD1 U4142 ( .I(n4321), .Z(n4281) );
  BUFFD1 U4143 ( .I(n4322), .Z(n4321) );
  BUFFD1 U4144 ( .I(n4317), .Z(n4308) );
  BUFFD1 U4145 ( .I(n4316), .Z(n4309) );
  BUFFD1 U4146 ( .I(n4325), .Z(n4310) );
  BUFFD1 U4147 ( .I(n4325), .Z(n4311) );
  BUFFD1 U4148 ( .I(n4325), .Z(n4312) );
  BUFFD1 U4149 ( .I(n4324), .Z(n4313) );
  BUFFD1 U4150 ( .I(n4324), .Z(n4314) );
  BUFFD1 U4151 ( .I(n4324), .Z(n4315) );
  BUFFD1 U4152 ( .I(n4323), .Z(n4316) );
  BUFFD1 U4153 ( .I(n4323), .Z(n4317) );
  BUFFD1 U4154 ( .I(n4323), .Z(n4318) );
  BUFFD1 U4155 ( .I(n4322), .Z(n4319) );
  BUFFD1 U4156 ( .I(n4322), .Z(n4320) );
  INVD1 U4157 ( .I(n20), .ZN(n4275) );
  INVD1 U4158 ( .I(n20), .ZN(n4274) );
  INVD1 U4159 ( .I(n25), .ZN(n4273) );
  INVD1 U4160 ( .I(n25), .ZN(n4272) );
  INVD1 U4161 ( .I(n22), .ZN(n4271) );
  INVD1 U4162 ( .I(n22), .ZN(n4270) );
  INVD1 U4163 ( .I(n19), .ZN(n4269) );
  INVD1 U4164 ( .I(n19), .ZN(n4268) );
  INVD1 U4165 ( .I(n21), .ZN(n4267) );
  INVD1 U4166 ( .I(n21), .ZN(n4266) );
  INVD1 U4167 ( .I(n26), .ZN(n4265) );
  INVD1 U4168 ( .I(n26), .ZN(n4264) );
  INVD1 U4169 ( .I(n23), .ZN(n4263) );
  INVD1 U4170 ( .I(n23), .ZN(n4262) );
  INVD1 U4171 ( .I(n17), .ZN(n4259) );
  INVD1 U4172 ( .I(n17), .ZN(n4258) );
  INVD1 U4173 ( .I(n13), .ZN(n4257) );
  INVD1 U4174 ( .I(n13), .ZN(n4256) );
  INVD1 U4175 ( .I(n11), .ZN(n4255) );
  INVD1 U4176 ( .I(n11), .ZN(n4254) );
  INVD1 U4177 ( .I(n12), .ZN(n4253) );
  INVD1 U4178 ( .I(n12), .ZN(n4252) );
  INVD1 U4179 ( .I(n14), .ZN(n4251) );
  INVD1 U4180 ( .I(n14), .ZN(n4250) );
  INVD1 U4181 ( .I(n24), .ZN(n4249) );
  INVD1 U4182 ( .I(n24), .ZN(n4248) );
  INVD1 U4183 ( .I(n15), .ZN(n4247) );
  INVD1 U4184 ( .I(n15), .ZN(n4246) );
  BUFFD1 U4185 ( .I(n4279), .Z(n4325) );
  BUFFD1 U4186 ( .I(n4279), .Z(n4324) );
  BUFFD1 U4187 ( .I(n4278), .Z(n4323) );
  BUFFD1 U4188 ( .I(n4278), .Z(n4322) );
  BUFFD1 U4189 ( .I(N44), .Z(n4241) );
  BUFFD1 U4190 ( .I(N44), .Z(n4242) );
  BUFFD1 U4191 ( .I(N44), .Z(n4243) );
  BUFFD1 U4192 ( .I(n4240), .Z(n4244) );
  BUFFD1 U4193 ( .I(n4240), .Z(n4245) );
  BUFFD1 U4194 ( .I(n4234), .Z(n4235) );
  BUFFD1 U4195 ( .I(n4234), .Z(n4236) );
  BUFFD1 U4196 ( .I(n4234), .Z(n4237) );
  BUFFD1 U4197 ( .I(n4233), .Z(n4238) );
  BUFFD1 U4198 ( .I(n4233), .Z(n4239) );
  INVD1 U4199 ( .I(n4331), .ZN(n4329) );
  INVD1 U4200 ( .I(n4331), .ZN(n4328) );
  INVD1 U4201 ( .I(n4331), .ZN(n4330) );
  BUFFD1 U4202 ( .I(n4280), .Z(n4279) );
  BUFFD1 U4203 ( .I(n4280), .Z(n4278) );
  INVD1 U4204 ( .I(n4327), .ZN(n4326) );
  XOR3D1 U4205 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n65), .Z(N84) );
  XOR3D1 U4206 ( .A1(DataI[0]), .A2(n66), .A3(n67), .Z(n65) );
  XOR3D1 U4207 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n68), .Z(n67) );
  XOR3D1 U4208 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n74), .Z(n73) );
  XOR3D1 U4209 ( .A1(n75), .A2(DataI[17]), .A3(n76), .Z(n74) );
  XOR3D1 U4210 ( .A1(n69), .A2(DataI[3]), .A3(n70), .Z(n68) );
  XOR3D1 U4211 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n71), .Z(n70) );
  XOR3D1 U4212 ( .A1(n72), .A2(DataI[10]), .A3(n73), .Z(n71) );
  XOR3D1 U4213 ( .A1(n87), .A2(N57), .A3(n88), .Z(n86) );
  XOR3D1 U4214 ( .A1(n3960), .A2(n3956), .A3(n83), .Z(n81) );
  XOR3D1 U4215 ( .A1(n4015), .A2(n4012), .A3(n80), .Z(n79) );
  BUFFD1 U4216 ( .I(N45), .Z(n4234) );
  INVD1 U4217 ( .I(n4231), .ZN(n4232) );
  BUFFD1 U4218 ( .I(n4332), .Z(n4240) );
  BUFFD1 U4219 ( .I(N45), .Z(n4233) );
  ND2D1 U4220 ( .A1(n101), .A2(n96), .ZN(n98) );
  ND2D1 U4221 ( .A1(n99), .A2(n100), .ZN(n94) );
  ND2D1 U4222 ( .A1(n95), .A2(n96), .ZN(n91) );
  INVD1 U4223 ( .I(n4045), .ZN(n4331) );
  INVD1 U4224 ( .I(ClockR), .ZN(n4327) );
  BUFFD1 U4225 ( .I(ClockW), .Z(n4280) );
  MUX4D0 U4226 ( .I0(n4106), .I1(n4104), .I2(n4105), .I3(n4103), .S0(N47), 
        .S1(N46), .Z(N80) );
  MUX4D0 U4227 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(N44), .S1(n4233), .Z(n4105) );
  MUX4D0 U4228 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n4244), .S1(n4234), .Z(
        n4104) );
  MUX4D0 U4229 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n4332), .S1(n4233), .Z(
        n4106) );
  MUX4D0 U4230 ( .I0(n4110), .I1(n4108), .I2(n4109), .I3(n4107), .S0(N47), 
        .S1(N46), .Z(N79) );
  MUX4D0 U4231 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(N44), .S1(n4237), .Z(n4109) );
  MUX4D0 U4232 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(N44), .S1(n4233), .Z(
        n4108) );
  MUX4D0 U4233 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(N44), .S1(n4239), .Z(n4110) );
  MUX4D0 U4234 ( .I0(n4130), .I1(n4128), .I2(n4129), .I3(n4127), .S0(N47), 
        .S1(N46), .Z(N74) );
  MUX4D0 U4235 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n4243), .S1(n4234), .Z(
        n4129) );
  MUX4D0 U4236 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n4243), .S1(n4234), .Z(
        n4128) );
  MUX4D0 U4237 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(N44), .S1(n4233), .Z(n4130) );
  MUX4D0 U4238 ( .I0(n4150), .I1(n4148), .I2(n4149), .I3(n4147), .S0(n4232), 
        .S1(n4333), .Z(N69) );
  MUX4D0 U4239 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n4240), .S1(n4236), .Z(
        n4149) );
  MUX4D0 U4240 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n4240), .S1(n4236), 
        .Z(n4148) );
  MUX4D0 U4241 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(N44), .S1(n4236), .Z(
        n4150) );
  MUX4D0 U4242 ( .I0(n4154), .I1(n4152), .I2(n4153), .I3(n4151), .S0(N47), 
        .S1(n4333), .Z(N68) );
  MUX4D0 U4243 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n4241), .S1(n4236), .Z(
        n4153) );
  MUX4D0 U4244 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n4242), .S1(n4236), 
        .Z(n4152) );
  MUX4D0 U4245 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n4244), .S1(n4236), .Z(
        n4154) );
  MUX4D0 U4246 ( .I0(n4178), .I1(n4176), .I2(n4177), .I3(n4175), .S0(N47), 
        .S1(n4333), .Z(N62) );
  MUX4D0 U4247 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n4241), .S1(n4236), .Z(
        n4177) );
  MUX4D0 U4248 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n4241), .S1(n4235), 
        .Z(n4176) );
  MUX4D0 U4249 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n4241), .S1(n4235), .Z(
        n4178) );
  MUX4D0 U4250 ( .I0(n4182), .I1(n4180), .I2(n4181), .I3(n4179), .S0(n4232), 
        .S1(N46), .Z(N61) );
  MUX4D0 U4251 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n4241), .S1(n4239), .Z(
        n4181) );
  MUX4D0 U4252 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n4241), .S1(n4237), 
        .Z(n4180) );
  MUX4D0 U4253 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n4241), .S1(n4238), .Z(
        n4182) );
  MUX4D0 U4254 ( .I0(n4206), .I1(n4204), .I2(n4205), .I3(n4203), .S0(n4232), 
        .S1(n4333), .Z(N55) );
  MUX4D0 U4255 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n4243), .S1(N45), .Z(
        n4205) );
  MUX4D0 U4256 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n4243), .S1(n4234), 
        .Z(n4204) );
  MUX4D0 U4257 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n4243), .S1(N45), .Z(
        n4206) );
  MUX4D0 U4258 ( .I0(n4210), .I1(n4208), .I2(n4209), .I3(n4207), .S0(n4232), 
        .S1(n4333), .Z(N54) );
  MUX4D0 U4259 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n4244), .S1(n4238), .Z(
        n4209) );
  MUX4D0 U4260 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n4244), .S1(n4238), 
        .Z(n4208) );
  MUX4D0 U4261 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n4244), .S1(n4238), .Z(
        n4210) );
  MUX4D0 U4262 ( .I0(n4222), .I1(n4220), .I2(n4221), .I3(n4219), .S0(n4232), 
        .S1(n4333), .Z(N51) );
  MUX4D0 U4263 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n4245), .S1(n4239), .Z(
        n4221) );
  MUX4D0 U4264 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n4245), .S1(n4239), 
        .Z(n4220) );
  MUX4D0 U4265 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n4245), .S1(n4239), .Z(
        n4222) );
  MUX4D0 U4266 ( .I0(n4226), .I1(n4224), .I2(n4225), .I3(n4223), .S0(n4232), 
        .S1(n4333), .Z(N50) );
  MUX4D0 U4267 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n4245), .S1(n4239), .Z(
        n4225) );
  MUX4D0 U4268 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n4245), .S1(n4239), 
        .Z(n4224) );
  MUX4D0 U4269 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n4245), .S1(n4239), .Z(
        n4226) );
  MUX4D0 U4270 ( .I0(n4126), .I1(n4124), .I2(n4125), .I3(n4123), .S0(N47), 
        .S1(N46), .Z(N75) );
  MUX4D0 U4271 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n4244), .S1(N45), .Z(n4125) );
  MUX4D0 U4272 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n4245), .S1(N45), .Z(
        n4124) );
  MUX4D0 U4273 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(N44), .S1(n4234), .Z(n4126) );
  MUX4D0 U4274 ( .I0(n4166), .I1(n4164), .I2(n4165), .I3(n4163), .S0(n4232), 
        .S1(n4333), .Z(N65) );
  MUX4D0 U4275 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(N44), .S1(n4237), .Z(
        n4165) );
  MUX4D0 U4276 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(N44), .S1(n4237), .Z(
        n4164) );
  MUX4D0 U4277 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n4245), .S1(n4237), .Z(
        n4166) );
  MUX4D0 U4278 ( .I0(n4194), .I1(n4192), .I2(n4193), .I3(n4191), .S0(n4232), 
        .S1(n4333), .Z(N58) );
  MUX4D0 U4279 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n4242), .S1(n4236), .Z(
        n4193) );
  MUX4D0 U4280 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n4242), .S1(n4237), 
        .Z(n4192) );
  MUX4D0 U4281 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n4242), .S1(n4238), .Z(
        n4194) );
  MUX4D0 U4282 ( .I0(n4198), .I1(n4196), .I2(n4197), .I3(n4195), .S0(n4232), 
        .S1(n4333), .Z(N57) );
  MUX4D0 U4283 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n4243), .S1(n4235), .Z(
        n4197) );
  MUX4D0 U4284 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n4243), .S1(N45), .Z(
        n4196) );
  MUX4D0 U4285 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n4243), .S1(N45), .Z(
        n4198) );
  MUX4D0 U4286 ( .I0(n4102), .I1(n4100), .I2(n4101), .I3(n4099), .S0(n4232), 
        .S1(n4333), .Z(N81) );
  MUX4D0 U4287 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n4240), .S1(n4233), .Z(
        n4101) );
  MUX4D0 U4288 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n4332), .S1(N45), .Z(
        n4100) );
  MUX4D0 U4289 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n4332), .S1(n4236), .Z(
        n4102) );
  MUX4D0 U4290 ( .I0(n4118), .I1(n4116), .I2(n4117), .I3(n4115), .S0(N47), 
        .S1(N46), .Z(N77) );
  MUX4D0 U4291 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n4240), .S1(N45), .Z(n4117) );
  MUX4D0 U4292 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n4332), .S1(n4239), .Z(
        n4116) );
  MUX4D0 U4293 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n4245), .S1(n4236), .Z(
        n4118) );
  MUX4D0 U4294 ( .I0(n4142), .I1(n4140), .I2(n4141), .I3(n4139), .S0(N47), 
        .S1(N46), .Z(N71) );
  MUX4D0 U4295 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n4242), .S1(n4235), .Z(
        n4141) );
  MUX4D0 U4296 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n4241), .S1(n4235), 
        .Z(n4140) );
  MUX4D0 U4297 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n4242), .S1(n4235), .Z(
        n4142) );
  MUX4D0 U4298 ( .I0(n4146), .I1(n4144), .I2(n4145), .I3(n4143), .S0(N47), 
        .S1(N46), .Z(N70) );
  MUX4D0 U4299 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n4241), .S1(n4235), .Z(
        n4145) );
  MUX4D0 U4300 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n4242), .S1(n4235), 
        .Z(n4144) );
  MUX4D0 U4301 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n4241), .S1(n4235), .Z(
        n4146) );
  MUX4D0 U4302 ( .I0(n4158), .I1(n4156), .I2(n4157), .I3(n4155), .S0(N47), 
        .S1(N46), .Z(N67) );
  MUX4D0 U4303 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n4245), .S1(n4236), .Z(
        n4157) );
  MUX4D0 U4304 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n4245), .S1(n4236), 
        .Z(n4156) );
  MUX4D0 U4305 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n4242), .S1(n4236), .Z(
        n4158) );
  MUX4D0 U4306 ( .I0(n4174), .I1(n4172), .I2(n4173), .I3(n4171), .S0(N47), 
        .S1(n4333), .Z(N63) );
  MUX4D0 U4307 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n4241), .S1(n4234), .Z(
        n4173) );
  MUX4D0 U4308 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n4241), .S1(n4233), 
        .Z(n4172) );
  MUX4D0 U4309 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n4241), .S1(n4234), .Z(
        n4174) );
  MUX4D0 U4310 ( .I0(n4186), .I1(n4184), .I2(n4185), .I3(n4183), .S0(n4232), 
        .S1(n4333), .Z(N60) );
  MUX4D0 U4311 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n4242), .S1(n4233), .Z(
        n4185) );
  MUX4D0 U4312 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n4242), .S1(n4233), 
        .Z(n4184) );
  MUX4D0 U4313 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n4242), .S1(n4233), .Z(
        n4186) );
  MUX4D0 U4314 ( .I0(n4202), .I1(n4200), .I2(n4201), .I3(n4199), .S0(n4232), 
        .S1(n4333), .Z(N56) );
  MUX4D0 U4315 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n4243), .S1(n4233), .Z(
        n4201) );
  MUX4D0 U4316 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n4243), .S1(n4234), 
        .Z(n4200) );
  MUX4D0 U4317 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n4243), .S1(n4233), .Z(
        n4202) );
  MUX4D0 U4318 ( .I0(n4214), .I1(n4212), .I2(n4213), .I3(n4211), .S0(n4232), 
        .S1(n4333), .Z(N53) );
  MUX4D0 U4319 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n4244), .S1(n4238), .Z(
        n4213) );
  MUX4D0 U4320 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n4244), .S1(n4238), 
        .Z(n4212) );
  MUX4D0 U4321 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n4244), .S1(n4238), .Z(
        n4214) );
  MUX4D0 U4322 ( .I0(n4218), .I1(n4216), .I2(n4217), .I3(n4215), .S0(n4232), 
        .S1(n4333), .Z(N52) );
  MUX4D0 U4323 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n4244), .S1(n4238), .Z(
        n4217) );
  MUX4D0 U4324 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n4244), .S1(n4238), 
        .Z(n4216) );
  MUX4D0 U4325 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n4244), .S1(n4238), .Z(
        n4218) );
  MUX4D0 U4326 ( .I0(n4122), .I1(n4120), .I2(n4121), .I3(n4119), .S0(N47), 
        .S1(n4333), .Z(N76) );
  MUX4D0 U4327 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n4243), .S1(n4234), .Z(
        n4121) );
  MUX4D0 U4328 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n4332), .S1(n4234), .Z(
        n4120) );
  MUX4D0 U4329 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n4243), .S1(n4237), .Z(
        n4122) );
  MUX4D0 U4330 ( .I0(n4138), .I1(n4136), .I2(n4137), .I3(n4135), .S0(n4232), 
        .S1(n4333), .Z(N72) );
  MUX4D0 U4331 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(N44), .S1(n4235), .Z(n4137) );
  MUX4D0 U4332 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n4241), .S1(n4235), .Z(
        n4136) );
  MUX4D0 U4333 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n4244), .S1(n4235), .Z(
        n4138) );
  MUX4D0 U4334 ( .I0(n4162), .I1(n4160), .I2(n4161), .I3(n4159), .S0(N47), 
        .S1(N46), .Z(N66) );
  MUX4D0 U4335 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n4332), .S1(n4237), .Z(
        n4161) );
  MUX4D0 U4336 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n4240), .S1(n4237), 
        .Z(n4160) );
  MUX4D0 U4337 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(N44), .S1(n4237), .Z(
        n4162) );
  MUX4D0 U4338 ( .I0(n4170), .I1(n4168), .I2(n4169), .I3(n4167), .S0(N47), 
        .S1(N46), .Z(N64) );
  MUX4D0 U4339 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n4240), .S1(n4237), .Z(
        n4169) );
  MUX4D0 U4340 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n4241), .S1(n4237), 
        .Z(n4168) );
  MUX4D0 U4341 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n4240), .S1(n4237), .Z(
        n4170) );
  MUX4D0 U4342 ( .I0(n4190), .I1(n4188), .I2(n4189), .I3(n4187), .S0(n4232), 
        .S1(n4333), .Z(N59) );
  MUX4D0 U4343 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n4242), .S1(n4233), .Z(
        n4189) );
  MUX4D0 U4344 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n4242), .S1(n4233), 
        .Z(n4188) );
  MUX4D0 U4345 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n4242), .S1(n4234), .Z(
        n4190) );
  MUX4D0 U4346 ( .I0(n4230), .I1(n4228), .I2(n4229), .I3(n4227), .S0(n4232), 
        .S1(n4333), .Z(N49) );
  MUX4D0 U4347 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n4245), .S1(n4239), .Z(
        n4229) );
  MUX4D0 U4348 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n4245), .S1(n4239), 
        .Z(n4228) );
  MUX4D0 U4349 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n4245), .S1(n4239), .Z(
        n4230) );
  MUX4D0 U4350 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n4245), .S1(n4239), 
        .Z(n4227) );
  MUX4D0 U4351 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n4332), .S1(n4234), .Z(
        n4099) );
  MUX4D0 U4352 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(N44), .S1(N45), .Z(n4103) );
  MUX4D0 U4353 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(N44), .S1(n4235), .Z(
        n4107) );
  MUX4D0 U4354 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n4240), .S1(n4238), .Z(
        n4115) );
  MUX4D0 U4355 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n4332), .S1(n4239), .Z(
        n4119) );
  MUX4D0 U4356 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n4240), .S1(n4233), .Z(
        n4123) );
  MUX4D0 U4357 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n4244), .S1(N45), .Z(
        n4127) );
  MUX4D0 U4358 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n4240), .S1(n4235), .Z(
        n4135) );
  MUX4D0 U4359 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n4241), .S1(n4235), 
        .Z(n4139) );
  MUX4D0 U4360 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n4242), .S1(n4235), 
        .Z(n4143) );
  MUX4D0 U4361 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n4240), .S1(n4236), 
        .Z(n4147) );
  MUX4D0 U4362 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n4245), .S1(n4236), 
        .Z(n4151) );
  MUX4D0 U4363 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n4245), .S1(n4236), 
        .Z(n4155) );
  MUX4D0 U4364 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n4332), .S1(n4237), 
        .Z(n4159) );
  MUX4D0 U4365 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n4240), .S1(n4237), 
        .Z(n4163) );
  MUX4D0 U4366 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n4240), .S1(n4237), 
        .Z(n4167) );
  MUX4D0 U4367 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n4241), .S1(N45), .Z(
        n4171) );
  MUX4D0 U4368 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n4241), .S1(n4236), 
        .Z(n4175) );
  MUX4D0 U4369 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n4241), .S1(n4235), 
        .Z(n4179) );
  MUX4D0 U4370 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n4242), .S1(n4234), 
        .Z(n4183) );
  MUX4D0 U4371 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n4242), .S1(n4233), 
        .Z(n4187) );
  MUX4D0 U4372 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n4242), .S1(n4237), 
        .Z(n4191) );
  MUX4D0 U4373 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n4243), .S1(N45), .Z(
        n4195) );
  MUX4D0 U4374 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n4243), .S1(n4234), 
        .Z(n4199) );
  MUX4D0 U4375 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n4243), .S1(n4233), 
        .Z(n4203) );
  MUX4D0 U4376 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n4244), .S1(n4238), 
        .Z(n4207) );
  MUX4D0 U4377 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n4244), .S1(n4238), 
        .Z(n4211) );
  MUX4D0 U4378 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n4244), .S1(n4238), 
        .Z(n4215) );
  MUX4D0 U4379 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n4245), .S1(n4239), 
        .Z(n4219) );
  MUX4D0 U4380 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n4245), .S1(n4239), 
        .Z(n4223) );
  BUFFD1 U4381 ( .I(N46), .Z(n4333) );
  MUX4D0 U4382 ( .I0(n4134), .I1(n4132), .I2(n4133), .I3(n4131), .S0(N47), 
        .S1(N46), .Z(N73) );
  MUX4D0 U4383 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n4243), .S1(n4233), .Z(
        n4133) );
  MUX4D0 U4384 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n4243), .S1(n4234), .Z(
        n4132) );
  MUX4D0 U4385 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n4240), .S1(n4237), .Z(
        n4134) );
  MUX4D0 U4386 ( .I0(n4114), .I1(n4112), .I2(n4113), .I3(n4111), .S0(N47), 
        .S1(N46), .Z(N78) );
  MUX4D0 U4387 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n4242), .S1(n4233), .Z(
        n4113) );
  MUX4D0 U4388 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n4240), .S1(n4239), .Z(
        n4112) );
  MUX4D0 U4389 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n4240), .S1(n4234), .Z(
        n4114) );
  MUX4D0 U4390 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n4243), .S1(n4234), .Z(
        n4111) );
  MUX4D0 U4391 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n4240), .S1(n4239), .Z(
        n4131) );
  ND2D1 U4392 ( .A1(AddrW[1]), .A2(n100), .ZN(n93) );
  ND2D1 U4393 ( .A1(AddrW[2]), .A2(AddrW[1]), .ZN(n90) );
  ND2D1 U4394 ( .A1(n101), .A2(AddrW[0]), .ZN(n97) );
  ND2D1 U4395 ( .A1(AddrW[2]), .A2(n99), .ZN(n92) );
  ND2D1 U4396 ( .A1(AddrW[0]), .A2(n95), .ZN(n89) );
  INR2D1 U4397 ( .A1(Write), .B1(AddrW[3]), .ZN(n101) );
  INVD1 U4398 ( .I(AddrW[1]), .ZN(n99) );
  INVD1 U4399 ( .I(AddrW[0]), .ZN(n96) );
  INVD1 U4400 ( .I(AddrW[2]), .ZN(n100) );
  AN2D1 U4401 ( .A1(Write), .A2(AddrW[3]), .Z(n95) );
  INR2D1 U4402 ( .A1(ClkW), .B1(N9), .ZN(ClockW) );
  INR2D1 U4403 ( .A1(ClkR), .B1(N9), .ZN(ClockR) );
  INVD0 U4404 ( .I(ChipEna), .ZN(N9) );
endmodule


module ClockComparator_0 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n5,
         n7, n8, n9, n1, n2, n3, n4, n6, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n152;

  AO211D1 U8 ( .A1(n7), .A2(n8), .B(N8), .C(N5), .Z(n9) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n5), .QN(N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n5), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n152), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n152), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(n1), .CP(ClockIn), .CDN(n5), .Q(\ClockInN[0] ), 
        .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(n27), .CP(ClockIn), .CDN(n5), .QN(n7) );
  DFSND1 ZeroCounters_reg ( .D(n49), .CP(ClockIn), .SDN(n152), .QN(n5) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(n6), .Z(n4) );
  BUFFD0 U7 ( .I(n10), .Z(n6) );
  BUFFD0 U9 ( .I(n11), .Z(n10) );
  BUFFD0 U10 ( .I(n12), .Z(n11) );
  BUFFD0 U11 ( .I(n13), .Z(n12) );
  BUFFD0 U12 ( .I(n14), .Z(n13) );
  BUFFD0 U13 ( .I(n15), .Z(n14) );
  BUFFD0 U14 ( .I(n16), .Z(n15) );
  BUFFD0 U15 ( .I(n17), .Z(n16) );
  BUFFD0 U16 ( .I(n18), .Z(n17) );
  BUFFD0 U17 ( .I(n19), .Z(n18) );
  BUFFD0 U18 ( .I(n20), .Z(n19) );
  BUFFD0 U19 ( .I(n21), .Z(n20) );
  BUFFD0 U20 ( .I(n22), .Z(n21) );
  BUFFD0 U21 ( .I(n23), .Z(n22) );
  BUFFD0 U22 ( .I(n24), .Z(n23) );
  BUFFD0 U23 ( .I(n25), .Z(n24) );
  BUFFD0 U24 ( .I(n148), .Z(n25) );
  BUFFD0 U25 ( .I(N5), .Z(n26) );
  BUFFD0 U26 ( .I(n28), .Z(n27) );
  BUFFD0 U27 ( .I(n29), .Z(n28) );
  BUFFD0 U28 ( .I(n30), .Z(n29) );
  BUFFD0 U29 ( .I(n31), .Z(n30) );
  BUFFD0 U30 ( .I(n32), .Z(n31) );
  BUFFD0 U31 ( .I(n33), .Z(n32) );
  BUFFD0 U32 ( .I(n34), .Z(n33) );
  BUFFD0 U33 ( .I(n35), .Z(n34) );
  BUFFD0 U34 ( .I(n36), .Z(n35) );
  BUFFD0 U35 ( .I(n37), .Z(n36) );
  BUFFD0 U36 ( .I(n38), .Z(n37) );
  BUFFD0 U37 ( .I(n39), .Z(n38) );
  BUFFD0 U38 ( .I(n40), .Z(n39) );
  BUFFD0 U39 ( .I(n41), .Z(n40) );
  BUFFD0 U40 ( .I(n42), .Z(n41) );
  BUFFD0 U41 ( .I(n43), .Z(n42) );
  BUFFD0 U42 ( .I(n44), .Z(n43) );
  BUFFD0 U43 ( .I(n45), .Z(n44) );
  BUFFD0 U44 ( .I(n46), .Z(n45) );
  BUFFD0 U45 ( .I(n47), .Z(n46) );
  BUFFD0 U46 ( .I(n145), .Z(n47) );
  BUFFD0 U47 ( .I(N6), .Z(n48) );
  BUFFD0 U48 ( .I(n52), .Z(n49) );
  BUFFD0 U49 ( .I(n26), .Z(n50) );
  BUFFD0 U50 ( .I(n48), .Z(n51) );
  BUFFD0 U51 ( .I(n55), .Z(n52) );
  BUFFD0 U52 ( .I(n50), .Z(n53) );
  BUFFD0 U53 ( .I(n51), .Z(n54) );
  BUFFD0 U54 ( .I(n58), .Z(n55) );
  BUFFD0 U55 ( .I(n53), .Z(n56) );
  BUFFD0 U56 ( .I(n54), .Z(n57) );
  BUFFD0 U57 ( .I(n61), .Z(n58) );
  BUFFD0 U58 ( .I(n56), .Z(n59) );
  BUFFD0 U59 ( .I(n57), .Z(n60) );
  BUFFD0 U60 ( .I(n64), .Z(n61) );
  BUFFD0 U61 ( .I(n59), .Z(n62) );
  BUFFD0 U62 ( .I(n60), .Z(n63) );
  BUFFD0 U63 ( .I(n67), .Z(n64) );
  BUFFD0 U64 ( .I(n62), .Z(n65) );
  BUFFD0 U65 ( .I(n63), .Z(n66) );
  BUFFD0 U66 ( .I(n70), .Z(n67) );
  BUFFD0 U67 ( .I(n65), .Z(n68) );
  BUFFD0 U68 ( .I(n66), .Z(n69) );
  BUFFD0 U69 ( .I(n73), .Z(n70) );
  BUFFD0 U70 ( .I(n68), .Z(n71) );
  BUFFD0 U71 ( .I(n69), .Z(n72) );
  BUFFD0 U72 ( .I(n76), .Z(n73) );
  BUFFD0 U73 ( .I(n71), .Z(n74) );
  BUFFD0 U74 ( .I(n72), .Z(n75) );
  BUFFD0 U75 ( .I(n77), .Z(n76) );
  BUFFD0 U76 ( .I(n82), .Z(n77) );
  BUFFD0 U77 ( .I(n74), .Z(n78) );
  BUFFD0 U78 ( .I(n75), .Z(n79) );
  BUFFD0 U79 ( .I(n78), .Z(n80) );
  BUFFD0 U80 ( .I(n79), .Z(n81) );
  BUFFD0 U81 ( .I(n85), .Z(n82) );
  BUFFD0 U82 ( .I(n80), .Z(n83) );
  BUFFD0 U83 ( .I(n81), .Z(n84) );
  BUFFD0 U84 ( .I(n86), .Z(n85) );
  BUFFD0 U85 ( .I(n91), .Z(n86) );
  BUFFD0 U86 ( .I(n83), .Z(n87) );
  BUFFD0 U87 ( .I(n84), .Z(n88) );
  BUFFD0 U88 ( .I(n87), .Z(n89) );
  BUFFD0 U89 ( .I(n88), .Z(n90) );
  BUFFD0 U90 ( .I(n94), .Z(n91) );
  BUFFD0 U91 ( .I(n89), .Z(n92) );
  BUFFD0 U92 ( .I(n90), .Z(n93) );
  BUFFD0 U93 ( .I(n95), .Z(n94) );
  BUFFD0 U94 ( .I(n96), .Z(n95) );
  BUFFD0 U95 ( .I(n97), .Z(n96) );
  BUFFD0 U96 ( .I(N9), .Z(n97) );
  BUFFD0 U97 ( .I(n92), .Z(n98) );
  BUFFD0 U98 ( .I(n93), .Z(n99) );
  BUFFD0 U99 ( .I(n98), .Z(n100) );
  BUFFD0 U100 ( .I(n99), .Z(n101) );
  BUFFD0 U101 ( .I(n100), .Z(n102) );
  BUFFD0 U102 ( .I(n101), .Z(n103) );
  BUFFD0 U103 ( .I(n102), .Z(n104) );
  BUFFD0 U104 ( .I(n103), .Z(n105) );
  BUFFD0 U105 ( .I(n104), .Z(n106) );
  BUFFD0 U106 ( .I(n105), .Z(n107) );
  BUFFD0 U107 ( .I(n106), .Z(n108) );
  BUFFD0 U108 ( .I(n107), .Z(n109) );
  BUFFD0 U109 ( .I(n108), .Z(n110) );
  BUFFD0 U110 ( .I(n109), .Z(n111) );
  BUFFD0 U111 ( .I(n110), .Z(n112) );
  BUFFD0 U112 ( .I(n111), .Z(n113) );
  BUFFD0 U113 ( .I(n112), .Z(n114) );
  BUFFD0 U114 ( .I(n113), .Z(n115) );
  BUFFD0 U115 ( .I(n114), .Z(n116) );
  BUFFD0 U116 ( .I(n115), .Z(n117) );
  BUFFD0 U117 ( .I(n116), .Z(n118) );
  BUFFD0 U118 ( .I(n117), .Z(n119) );
  BUFFD0 U119 ( .I(n118), .Z(n120) );
  BUFFD0 U120 ( .I(n119), .Z(n121) );
  BUFFD0 U121 ( .I(n120), .Z(n122) );
  BUFFD0 U122 ( .I(n121), .Z(n123) );
  BUFFD0 U123 ( .I(n122), .Z(n124) );
  BUFFD0 U124 ( .I(n123), .Z(n125) );
  BUFFD0 U125 ( .I(n124), .Z(n126) );
  BUFFD0 U126 ( .I(n125), .Z(n127) );
  BUFFD0 U127 ( .I(n126), .Z(n128) );
  BUFFD0 U128 ( .I(n127), .Z(n129) );
  BUFFD0 U129 ( .I(n128), .Z(n130) );
  BUFFD0 U130 ( .I(n129), .Z(n131) );
  BUFFD0 U131 ( .I(n130), .Z(n132) );
  BUFFD0 U132 ( .I(n131), .Z(n133) );
  BUFFD0 U133 ( .I(n132), .Z(n134) );
  BUFFD0 U134 ( .I(n133), .Z(n135) );
  BUFFD0 U135 ( .I(n134), .Z(n136) );
  BUFFD0 U136 ( .I(n135), .Z(n137) );
  BUFFD0 U137 ( .I(n136), .Z(n138) );
  BUFFD0 U138 ( .I(n137), .Z(n139) );
  BUFFD0 U139 ( .I(n138), .Z(n140) );
  BUFFD0 U140 ( .I(n139), .Z(n141) );
  BUFFD0 U141 ( .I(n140), .Z(n142) );
  BUFFD0 U142 ( .I(n141), .Z(n143) );
  BUFFD0 U143 ( .I(n142), .Z(n144) );
  CKBD0 U144 ( .CLK(n143), .C(n145) );
  BUFFD0 U145 ( .I(n144), .Z(n146) );
  BUFFD0 U146 ( .I(\ClockInN[0] ), .Z(n147) );
  XNR2D0 U147 ( .A1(n147), .A2(n7), .ZN(N6) );
  CKBD0 U148 ( .CLK(n146), .C(n148) );
  INVD1 U149 ( .I(Reset), .ZN(n152) );
  NR2D1 U150 ( .A1(n145), .A2(n148), .ZN(N9) );
  OAI21D1 U151 ( .A1(n8), .A2(n7), .B(n9), .ZN(N20) );
  NR2D1 U152 ( .A1(N19), .A2(N7), .ZN(n8) );
  XNR2D1 U153 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module VFO_0 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n17, n18, n19, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n20, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_0_DW01_dec_0 \Sampler/sub_193  ( .A({n64, n182, DivideFactor[3], n123, 
        n240, n300}), .SUM({N40, N39, N38, N37, N36, N35}) );
  VFO_0_DW01_inc_0 \Sampler/add_190  ( .A({n64, n182, DivideFactor[3], n123, 
        n240, n300}), .SUM({N32, N31, N30, N29, N28, N27}) );
  VFO_0_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n17), .CP(FastClock), .CDN(n416), .Q(ClockOut)
         );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(n2), .E(n361), .CP(Sample), .CDN(n416), 
        .Q(DivideFactor[5]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(n65), .E(n361), .CP(Sample), .CDN(n416), 
        .Q(DivideFactor[2]) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n124), .CP(Sample), .SDN(n416), .Q(
        DivideFactor[4]), .QN(n428) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n183), .CP(Sample), .SDN(n416), .Q(
        DivideFactor[1]), .QN(n440) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n242), .CP(Sample), .SDN(n416), .Q(
        DivideFactor[0]), .QN(n438) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(n301), .E(n361), .CP(Sample), .CDN(n416), 
        .Q(DivideFactor[3]), .QN(n433) );
  INVD4 U3 ( .I(n1), .ZN(N54) );
  MUX2D0 U4 ( .I0(n415), .I1(n427), .S(AdjustFreq[0]), .Z(n1) );
  BUFFD0 U5 ( .I(n5), .Z(n2) );
  BUFFD0 U6 ( .I(N55), .Z(n3) );
  BUFFD0 U7 ( .I(n3), .Z(n4) );
  BUFFD0 U8 ( .I(n6), .Z(n5) );
  BUFFD0 U9 ( .I(n7), .Z(n6) );
  BUFFD0 U10 ( .I(n8), .Z(n7) );
  BUFFD0 U11 ( .I(n9), .Z(n8) );
  BUFFD0 U12 ( .I(n10), .Z(n9) );
  BUFFD0 U13 ( .I(n11), .Z(n10) );
  BUFFD0 U14 ( .I(n12), .Z(n11) );
  BUFFD0 U15 ( .I(n13), .Z(n12) );
  BUFFD0 U16 ( .I(n14), .Z(n13) );
  BUFFD0 U17 ( .I(n15), .Z(n14) );
  BUFFD0 U18 ( .I(n16), .Z(n15) );
  BUFFD0 U19 ( .I(n20), .Z(n16) );
  BUFFD0 U20 ( .I(n22), .Z(n20) );
  BUFFD0 U21 ( .I(n23), .Z(n22) );
  BUFFD0 U22 ( .I(n24), .Z(n23) );
  BUFFD0 U23 ( .I(n25), .Z(n24) );
  BUFFD0 U24 ( .I(n26), .Z(n25) );
  BUFFD0 U25 ( .I(n27), .Z(n26) );
  BUFFD0 U26 ( .I(n28), .Z(n27) );
  BUFFD0 U27 ( .I(n29), .Z(n28) );
  BUFFD0 U28 ( .I(n30), .Z(n29) );
  BUFFD0 U29 ( .I(n31), .Z(n30) );
  BUFFD0 U30 ( .I(n32), .Z(n31) );
  BUFFD0 U31 ( .I(n33), .Z(n32) );
  BUFFD0 U32 ( .I(n34), .Z(n33) );
  BUFFD0 U33 ( .I(n35), .Z(n34) );
  BUFFD0 U34 ( .I(n36), .Z(n35) );
  BUFFD0 U35 ( .I(n37), .Z(n36) );
  BUFFD0 U36 ( .I(n38), .Z(n37) );
  BUFFD0 U37 ( .I(n39), .Z(n38) );
  BUFFD0 U38 ( .I(n40), .Z(n39) );
  BUFFD0 U39 ( .I(n41), .Z(n40) );
  BUFFD0 U40 ( .I(n42), .Z(n41) );
  BUFFD0 U41 ( .I(n43), .Z(n42) );
  BUFFD0 U42 ( .I(n44), .Z(n43) );
  BUFFD0 U43 ( .I(n45), .Z(n44) );
  BUFFD0 U44 ( .I(n46), .Z(n45) );
  BUFFD0 U45 ( .I(n47), .Z(n46) );
  BUFFD0 U46 ( .I(n48), .Z(n47) );
  BUFFD0 U47 ( .I(n49), .Z(n48) );
  BUFFD0 U48 ( .I(n50), .Z(n49) );
  BUFFD0 U49 ( .I(n51), .Z(n50) );
  BUFFD0 U50 ( .I(n52), .Z(n51) );
  BUFFD0 U51 ( .I(n53), .Z(n52) );
  BUFFD0 U52 ( .I(n54), .Z(n53) );
  BUFFD0 U53 ( .I(n55), .Z(n54) );
  BUFFD0 U54 ( .I(n56), .Z(n55) );
  BUFFD0 U55 ( .I(n57), .Z(n56) );
  BUFFD0 U56 ( .I(n58), .Z(n57) );
  BUFFD0 U57 ( .I(n59), .Z(n58) );
  BUFFD0 U58 ( .I(n60), .Z(n59) );
  BUFFD0 U59 ( .I(n61), .Z(n60) );
  BUFFD0 U60 ( .I(n62), .Z(n61) );
  BUFFD0 U61 ( .I(n4), .Z(n62) );
  BUFFD0 U62 ( .I(DivideFactor[5]), .Z(n63) );
  CKBD0 U63 ( .CLK(n63), .C(n64) );
  BUFFD0 U64 ( .I(n69), .Z(n65) );
  BUFFD0 U65 ( .I(N49), .Z(n66) );
  BUFFD0 U66 ( .I(n66), .Z(n67) );
  BUFFD0 U67 ( .I(n67), .Z(n68) );
  BUFFD0 U68 ( .I(n70), .Z(n69) );
  BUFFD0 U69 ( .I(n71), .Z(n70) );
  BUFFD0 U70 ( .I(n72), .Z(n71) );
  BUFFD0 U71 ( .I(n73), .Z(n72) );
  BUFFD0 U72 ( .I(n74), .Z(n73) );
  BUFFD0 U73 ( .I(n75), .Z(n74) );
  BUFFD0 U74 ( .I(n76), .Z(n75) );
  BUFFD0 U75 ( .I(n77), .Z(n76) );
  BUFFD0 U76 ( .I(n78), .Z(n77) );
  BUFFD0 U77 ( .I(n79), .Z(n78) );
  BUFFD0 U78 ( .I(n80), .Z(n79) );
  BUFFD0 U79 ( .I(n81), .Z(n80) );
  BUFFD0 U80 ( .I(n82), .Z(n81) );
  BUFFD0 U81 ( .I(n83), .Z(n82) );
  BUFFD0 U82 ( .I(n84), .Z(n83) );
  BUFFD0 U83 ( .I(n85), .Z(n84) );
  BUFFD0 U84 ( .I(n86), .Z(n85) );
  BUFFD0 U85 ( .I(n87), .Z(n86) );
  BUFFD0 U86 ( .I(n88), .Z(n87) );
  BUFFD0 U87 ( .I(n89), .Z(n88) );
  BUFFD0 U88 ( .I(n90), .Z(n89) );
  BUFFD0 U89 ( .I(n91), .Z(n90) );
  BUFFD0 U90 ( .I(n92), .Z(n91) );
  BUFFD0 U91 ( .I(n93), .Z(n92) );
  BUFFD0 U92 ( .I(n94), .Z(n93) );
  BUFFD0 U93 ( .I(n95), .Z(n94) );
  BUFFD0 U94 ( .I(n96), .Z(n95) );
  BUFFD0 U95 ( .I(n97), .Z(n96) );
  BUFFD0 U96 ( .I(n98), .Z(n97) );
  BUFFD0 U97 ( .I(n99), .Z(n98) );
  BUFFD0 U98 ( .I(n100), .Z(n99) );
  BUFFD0 U99 ( .I(n101), .Z(n100) );
  BUFFD0 U100 ( .I(n102), .Z(n101) );
  BUFFD0 U101 ( .I(n103), .Z(n102) );
  BUFFD0 U102 ( .I(n104), .Z(n103) );
  BUFFD0 U103 ( .I(n105), .Z(n104) );
  BUFFD0 U104 ( .I(n106), .Z(n105) );
  BUFFD0 U105 ( .I(n107), .Z(n106) );
  BUFFD0 U106 ( .I(n108), .Z(n107) );
  BUFFD0 U107 ( .I(n109), .Z(n108) );
  BUFFD0 U108 ( .I(n110), .Z(n109) );
  BUFFD0 U109 ( .I(n111), .Z(n110) );
  BUFFD0 U110 ( .I(n112), .Z(n111) );
  BUFFD0 U111 ( .I(n113), .Z(n112) );
  BUFFD0 U112 ( .I(n114), .Z(n113) );
  BUFFD0 U113 ( .I(n115), .Z(n114) );
  BUFFD0 U114 ( .I(n116), .Z(n115) );
  BUFFD0 U115 ( .I(n117), .Z(n116) );
  BUFFD0 U116 ( .I(n118), .Z(n117) );
  BUFFD0 U117 ( .I(n119), .Z(n118) );
  BUFFD0 U118 ( .I(n120), .Z(n119) );
  BUFFD0 U119 ( .I(n121), .Z(n120) );
  BUFFD0 U120 ( .I(n68), .Z(n121) );
  BUFFD0 U121 ( .I(DivideFactor[2]), .Z(n122) );
  CKBD0 U122 ( .CLK(n122), .C(n123) );
  BUFFD0 U123 ( .I(n127), .Z(n124) );
  BUFFD0 U124 ( .I(n19), .Z(n125) );
  BUFFD0 U125 ( .I(n125), .Z(n126) );
  BUFFD0 U126 ( .I(n128), .Z(n127) );
  BUFFD0 U127 ( .I(n129), .Z(n128) );
  BUFFD0 U128 ( .I(n130), .Z(n129) );
  BUFFD0 U129 ( .I(n131), .Z(n130) );
  BUFFD0 U130 ( .I(n132), .Z(n131) );
  BUFFD0 U131 ( .I(n133), .Z(n132) );
  BUFFD0 U132 ( .I(n134), .Z(n133) );
  BUFFD0 U133 ( .I(n135), .Z(n134) );
  BUFFD0 U134 ( .I(n136), .Z(n135) );
  BUFFD0 U135 ( .I(n137), .Z(n136) );
  BUFFD0 U136 ( .I(n138), .Z(n137) );
  BUFFD0 U137 ( .I(n139), .Z(n138) );
  BUFFD0 U138 ( .I(n140), .Z(n139) );
  BUFFD0 U139 ( .I(n141), .Z(n140) );
  BUFFD0 U140 ( .I(n142), .Z(n141) );
  BUFFD0 U141 ( .I(n143), .Z(n142) );
  BUFFD0 U142 ( .I(n144), .Z(n143) );
  BUFFD0 U143 ( .I(n145), .Z(n144) );
  BUFFD0 U144 ( .I(n146), .Z(n145) );
  BUFFD0 U145 ( .I(n147), .Z(n146) );
  BUFFD0 U146 ( .I(n148), .Z(n147) );
  BUFFD0 U147 ( .I(n149), .Z(n148) );
  BUFFD0 U148 ( .I(n150), .Z(n149) );
  BUFFD0 U149 ( .I(n151), .Z(n150) );
  BUFFD0 U150 ( .I(n152), .Z(n151) );
  BUFFD0 U151 ( .I(n153), .Z(n152) );
  BUFFD0 U152 ( .I(n154), .Z(n153) );
  BUFFD0 U153 ( .I(n155), .Z(n154) );
  BUFFD0 U154 ( .I(n156), .Z(n155) );
  BUFFD0 U155 ( .I(n157), .Z(n156) );
  BUFFD0 U156 ( .I(n158), .Z(n157) );
  BUFFD0 U157 ( .I(n159), .Z(n158) );
  BUFFD0 U158 ( .I(n160), .Z(n159) );
  BUFFD0 U159 ( .I(n161), .Z(n160) );
  CKBXD0 U160 ( .I(DivideFactor[4]), .Z(n182) );
  BUFFD0 U161 ( .I(n162), .Z(n161) );
  BUFFD0 U162 ( .I(n163), .Z(n162) );
  BUFFD0 U163 ( .I(n164), .Z(n163) );
  BUFFD0 U164 ( .I(n165), .Z(n164) );
  BUFFD0 U165 ( .I(n166), .Z(n165) );
  BUFFD0 U166 ( .I(n167), .Z(n166) );
  BUFFD0 U167 ( .I(n168), .Z(n167) );
  BUFFD0 U168 ( .I(n169), .Z(n168) );
  BUFFD0 U169 ( .I(n170), .Z(n169) );
  BUFFD0 U170 ( .I(n171), .Z(n170) );
  BUFFD0 U171 ( .I(n172), .Z(n171) );
  BUFFD0 U172 ( .I(n173), .Z(n172) );
  BUFFD0 U173 ( .I(n174), .Z(n173) );
  BUFFD0 U174 ( .I(n175), .Z(n174) );
  BUFFD0 U175 ( .I(n176), .Z(n175) );
  BUFFD0 U176 ( .I(n177), .Z(n176) );
  BUFFD0 U177 ( .I(n178), .Z(n177) );
  BUFFD0 U178 ( .I(n179), .Z(n178) );
  BUFFD0 U179 ( .I(n180), .Z(n179) );
  BUFFD0 U180 ( .I(n181), .Z(n180) );
  BUFFD0 U181 ( .I(n126), .Z(n181) );
  BUFFD0 U182 ( .I(n186), .Z(n183) );
  BUFFD0 U183 ( .I(n18), .Z(n184) );
  BUFFD0 U184 ( .I(n184), .Z(n185) );
  BUFFD0 U185 ( .I(n187), .Z(n186) );
  BUFFD0 U186 ( .I(n188), .Z(n187) );
  BUFFD0 U187 ( .I(n189), .Z(n188) );
  BUFFD0 U188 ( .I(n190), .Z(n189) );
  BUFFD0 U189 ( .I(n191), .Z(n190) );
  BUFFD0 U190 ( .I(n192), .Z(n191) );
  BUFFD0 U191 ( .I(n193), .Z(n192) );
  BUFFD0 U192 ( .I(n194), .Z(n193) );
  BUFFD0 U193 ( .I(n195), .Z(n194) );
  BUFFD0 U194 ( .I(n196), .Z(n195) );
  BUFFD0 U195 ( .I(n197), .Z(n196) );
  BUFFD0 U196 ( .I(n198), .Z(n197) );
  BUFFD0 U197 ( .I(n199), .Z(n198) );
  BUFFD0 U198 ( .I(n200), .Z(n199) );
  BUFFD0 U199 ( .I(n201), .Z(n200) );
  BUFFD0 U200 ( .I(n202), .Z(n201) );
  BUFFD0 U201 ( .I(n203), .Z(n202) );
  BUFFD0 U202 ( .I(n204), .Z(n203) );
  BUFFD0 U203 ( .I(n205), .Z(n204) );
  BUFFD0 U204 ( .I(n206), .Z(n205) );
  BUFFD0 U205 ( .I(n207), .Z(n206) );
  BUFFD0 U206 ( .I(n208), .Z(n207) );
  BUFFD0 U207 ( .I(n209), .Z(n208) );
  BUFFD0 U208 ( .I(n210), .Z(n209) );
  BUFFD0 U209 ( .I(n211), .Z(n210) );
  BUFFD0 U210 ( .I(n212), .Z(n211) );
  BUFFD0 U211 ( .I(n213), .Z(n212) );
  BUFFD0 U212 ( .I(n214), .Z(n213) );
  BUFFD0 U213 ( .I(n215), .Z(n214) );
  BUFFD0 U214 ( .I(n216), .Z(n215) );
  BUFFD0 U215 ( .I(n217), .Z(n216) );
  BUFFD0 U216 ( .I(n218), .Z(n217) );
  BUFFD0 U217 ( .I(n219), .Z(n218) );
  BUFFD0 U218 ( .I(n220), .Z(n219) );
  BUFFD0 U219 ( .I(n221), .Z(n220) );
  BUFFD0 U220 ( .I(n222), .Z(n221) );
  BUFFD0 U221 ( .I(n223), .Z(n222) );
  BUFFD0 U222 ( .I(n224), .Z(n223) );
  BUFFD0 U223 ( .I(n225), .Z(n224) );
  BUFFD0 U224 ( .I(n226), .Z(n225) );
  BUFFD0 U225 ( .I(n227), .Z(n226) );
  BUFFD0 U226 ( .I(n228), .Z(n227) );
  BUFFD0 U227 ( .I(n229), .Z(n228) );
  BUFFD0 U228 ( .I(n230), .Z(n229) );
  BUFFD0 U229 ( .I(n231), .Z(n230) );
  BUFFD0 U230 ( .I(n232), .Z(n231) );
  BUFFD0 U231 ( .I(n233), .Z(n232) );
  BUFFD0 U232 ( .I(n234), .Z(n233) );
  BUFFD0 U233 ( .I(n235), .Z(n234) );
  BUFFD0 U234 ( .I(n236), .Z(n235) );
  BUFFD0 U235 ( .I(n237), .Z(n236) );
  BUFFD0 U236 ( .I(n238), .Z(n237) );
  BUFFD0 U237 ( .I(n239), .Z(n238) );
  BUFFD0 U238 ( .I(n185), .Z(n239) );
  BUFFD0 U239 ( .I(n241), .Z(n240) );
  BUFFD0 U240 ( .I(DivideFactor[1]), .Z(n241) );
  BUFFD0 U241 ( .I(n245), .Z(n242) );
  BUFFD0 U242 ( .I(n21), .Z(n243) );
  BUFFD0 U243 ( .I(n243), .Z(n244) );
  BUFFD0 U244 ( .I(n246), .Z(n245) );
  BUFFD0 U245 ( .I(n247), .Z(n246) );
  BUFFD0 U246 ( .I(n248), .Z(n247) );
  BUFFD0 U247 ( .I(n249), .Z(n248) );
  BUFFD0 U248 ( .I(n250), .Z(n249) );
  BUFFD0 U249 ( .I(n251), .Z(n250) );
  BUFFD0 U250 ( .I(n252), .Z(n251) );
  BUFFD0 U251 ( .I(n253), .Z(n252) );
  BUFFD0 U252 ( .I(n254), .Z(n253) );
  BUFFD0 U253 ( .I(n255), .Z(n254) );
  BUFFD0 U254 ( .I(n256), .Z(n255) );
  BUFFD0 U255 ( .I(n257), .Z(n256) );
  BUFFD0 U256 ( .I(n258), .Z(n257) );
  BUFFD0 U257 ( .I(n259), .Z(n258) );
  BUFFD0 U258 ( .I(n260), .Z(n259) );
  BUFFD0 U259 ( .I(n261), .Z(n260) );
  BUFFD0 U260 ( .I(n262), .Z(n261) );
  BUFFD0 U261 ( .I(n263), .Z(n262) );
  BUFFD0 U262 ( .I(n264), .Z(n263) );
  BUFFD0 U263 ( .I(n265), .Z(n264) );
  BUFFD0 U264 ( .I(n266), .Z(n265) );
  BUFFD0 U265 ( .I(n267), .Z(n266) );
  BUFFD0 U266 ( .I(n268), .Z(n267) );
  BUFFD0 U267 ( .I(n269), .Z(n268) );
  BUFFD0 U268 ( .I(n270), .Z(n269) );
  BUFFD0 U269 ( .I(n271), .Z(n270) );
  BUFFD0 U270 ( .I(n272), .Z(n271) );
  BUFFD0 U271 ( .I(n273), .Z(n272) );
  BUFFD0 U272 ( .I(n274), .Z(n273) );
  BUFFD0 U273 ( .I(n275), .Z(n274) );
  BUFFD0 U274 ( .I(n276), .Z(n275) );
  BUFFD0 U275 ( .I(n277), .Z(n276) );
  BUFFD0 U276 ( .I(n278), .Z(n277) );
  BUFFD0 U277 ( .I(n279), .Z(n278) );
  BUFFD0 U278 ( .I(n280), .Z(n279) );
  BUFFD0 U279 ( .I(n281), .Z(n280) );
  BUFFD0 U280 ( .I(n282), .Z(n281) );
  BUFFD0 U281 ( .I(n283), .Z(n282) );
  BUFFD0 U282 ( .I(n284), .Z(n283) );
  BUFFD0 U283 ( .I(n285), .Z(n284) );
  BUFFD0 U284 ( .I(n286), .Z(n285) );
  BUFFD0 U285 ( .I(n287), .Z(n286) );
  BUFFD0 U286 ( .I(n288), .Z(n287) );
  BUFFD0 U287 ( .I(n289), .Z(n288) );
  BUFFD0 U288 ( .I(n290), .Z(n289) );
  BUFFD0 U289 ( .I(n291), .Z(n290) );
  BUFFD0 U290 ( .I(n292), .Z(n291) );
  BUFFD0 U291 ( .I(n293), .Z(n292) );
  BUFFD0 U292 ( .I(n294), .Z(n293) );
  BUFFD0 U293 ( .I(n295), .Z(n294) );
  BUFFD0 U294 ( .I(n296), .Z(n295) );
  BUFFD0 U295 ( .I(n297), .Z(n296) );
  BUFFD0 U296 ( .I(n298), .Z(n297) );
  BUFFD0 U297 ( .I(n244), .Z(n298) );
  BUFFD0 U298 ( .I(DivideFactor[0]), .Z(n299) );
  CKBXD0 U299 ( .I(n299), .Z(n300) );
  BUFFD0 U300 ( .I(n305), .Z(n301) );
  BUFFD0 U301 ( .I(N51), .Z(n302) );
  BUFFD0 U302 ( .I(n302), .Z(n303) );
  BUFFD0 U303 ( .I(n303), .Z(n304) );
  BUFFD0 U304 ( .I(n306), .Z(n305) );
  BUFFD0 U305 ( .I(n307), .Z(n306) );
  BUFFD0 U306 ( .I(n308), .Z(n307) );
  BUFFD0 U307 ( .I(n309), .Z(n308) );
  BUFFD0 U308 ( .I(n310), .Z(n309) );
  BUFFD0 U309 ( .I(n311), .Z(n310) );
  BUFFD0 U310 ( .I(n312), .Z(n311) );
  BUFFD0 U311 ( .I(n313), .Z(n312) );
  BUFFD0 U312 ( .I(n314), .Z(n313) );
  BUFFD0 U313 ( .I(n315), .Z(n314) );
  BUFFD0 U314 ( .I(n316), .Z(n315) );
  BUFFD0 U315 ( .I(n317), .Z(n316) );
  BUFFD0 U316 ( .I(n318), .Z(n317) );
  BUFFD0 U317 ( .I(n319), .Z(n318) );
  BUFFD0 U318 ( .I(n320), .Z(n319) );
  BUFFD0 U319 ( .I(n321), .Z(n320) );
  BUFFD0 U320 ( .I(n322), .Z(n321) );
  BUFFD0 U321 ( .I(n323), .Z(n322) );
  BUFFD0 U322 ( .I(n324), .Z(n323) );
  BUFFD0 U323 ( .I(n325), .Z(n324) );
  BUFFD0 U324 ( .I(n326), .Z(n325) );
  BUFFD0 U325 ( .I(n327), .Z(n326) );
  BUFFD0 U326 ( .I(n328), .Z(n327) );
  BUFFD0 U327 ( .I(n329), .Z(n328) );
  BUFFD0 U328 ( .I(n330), .Z(n329) );
  BUFFD0 U329 ( .I(n331), .Z(n330) );
  BUFFD0 U330 ( .I(n332), .Z(n331) );
  BUFFD0 U331 ( .I(n333), .Z(n332) );
  BUFFD0 U332 ( .I(n334), .Z(n333) );
  BUFFD0 U333 ( .I(n335), .Z(n334) );
  BUFFD0 U334 ( .I(n336), .Z(n335) );
  BUFFD0 U335 ( .I(n337), .Z(n336) );
  BUFFD0 U336 ( .I(n338), .Z(n337) );
  BUFFD0 U337 ( .I(n339), .Z(n338) );
  BUFFD0 U338 ( .I(n340), .Z(n339) );
  BUFFD0 U339 ( .I(n341), .Z(n340) );
  BUFFD0 U340 ( .I(n342), .Z(n341) );
  BUFFD0 U341 ( .I(n343), .Z(n342) );
  BUFFD0 U342 ( .I(n344), .Z(n343) );
  BUFFD0 U343 ( .I(n345), .Z(n344) );
  BUFFD0 U344 ( .I(n346), .Z(n345) );
  BUFFD0 U345 ( .I(n347), .Z(n346) );
  BUFFD0 U346 ( .I(n348), .Z(n347) );
  BUFFD0 U347 ( .I(n349), .Z(n348) );
  BUFFD0 U348 ( .I(n350), .Z(n349) );
  BUFFD0 U349 ( .I(n351), .Z(n350) );
  BUFFD0 U350 ( .I(n352), .Z(n351) );
  BUFFD0 U351 ( .I(n353), .Z(n352) );
  BUFFD0 U352 ( .I(n354), .Z(n353) );
  BUFFD0 U353 ( .I(n355), .Z(n354) );
  BUFFD0 U354 ( .I(n356), .Z(n355) );
  BUFFD0 U355 ( .I(n357), .Z(n356) );
  BUFFD0 U356 ( .I(n358), .Z(n357) );
  BUFFD0 U357 ( .I(n359), .Z(n358) );
  BUFFD0 U358 ( .I(n304), .Z(n359) );
  BUFFD0 U359 ( .I(n362), .Z(n360) );
  BUFFD0 U360 ( .I(n360), .Z(n361) );
  BUFFD0 U361 ( .I(n363), .Z(n362) );
  BUFFD0 U362 ( .I(n364), .Z(n363) );
  BUFFD0 U363 ( .I(n365), .Z(n364) );
  BUFFD0 U364 ( .I(n366), .Z(n365) );
  BUFFD0 U365 ( .I(n367), .Z(n366) );
  BUFFD0 U366 ( .I(n368), .Z(n367) );
  BUFFD0 U367 ( .I(n369), .Z(n368) );
  BUFFD0 U368 ( .I(n370), .Z(n369) );
  BUFFD0 U369 ( .I(n371), .Z(n370) );
  BUFFD0 U370 ( .I(n372), .Z(n371) );
  BUFFD0 U371 ( .I(n373), .Z(n372) );
  BUFFD0 U372 ( .I(n374), .Z(n373) );
  BUFFD0 U373 ( .I(n375), .Z(n374) );
  BUFFD0 U374 ( .I(n376), .Z(n375) );
  BUFFD0 U375 ( .I(n377), .Z(n376) );
  BUFFD0 U376 ( .I(n378), .Z(n377) );
  BUFFD0 U377 ( .I(n379), .Z(n378) );
  BUFFD0 U378 ( .I(n380), .Z(n379) );
  BUFFD0 U379 ( .I(n381), .Z(n380) );
  BUFFD0 U380 ( .I(n382), .Z(n381) );
  BUFFD0 U381 ( .I(n383), .Z(n382) );
  BUFFD0 U382 ( .I(n384), .Z(n383) );
  BUFFD0 U383 ( .I(n385), .Z(n384) );
  BUFFD0 U384 ( .I(n386), .Z(n385) );
  BUFFD0 U385 ( .I(n387), .Z(n386) );
  BUFFD0 U386 ( .I(n388), .Z(n387) );
  BUFFD0 U387 ( .I(n389), .Z(n388) );
  BUFFD0 U388 ( .I(n390), .Z(n389) );
  BUFFD0 U389 ( .I(n391), .Z(n390) );
  BUFFD0 U390 ( .I(n392), .Z(n391) );
  BUFFD0 U391 ( .I(n393), .Z(n392) );
  BUFFD0 U392 ( .I(n394), .Z(n393) );
  BUFFD0 U393 ( .I(n395), .Z(n394) );
  BUFFD0 U394 ( .I(n396), .Z(n395) );
  BUFFD0 U395 ( .I(n397), .Z(n396) );
  BUFFD0 U396 ( .I(n398), .Z(n397) );
  BUFFD0 U397 ( .I(n399), .Z(n398) );
  BUFFD0 U398 ( .I(n400), .Z(n399) );
  BUFFD0 U399 ( .I(n401), .Z(n400) );
  BUFFD0 U400 ( .I(n402), .Z(n401) );
  BUFFD0 U401 ( .I(n403), .Z(n402) );
  BUFFD0 U402 ( .I(n404), .Z(n403) );
  BUFFD0 U403 ( .I(n405), .Z(n404) );
  BUFFD0 U404 ( .I(n406), .Z(n405) );
  BUFFD0 U405 ( .I(n407), .Z(n406) );
  BUFFD0 U406 ( .I(n408), .Z(n407) );
  BUFFD0 U407 ( .I(n409), .Z(n408) );
  BUFFD0 U408 ( .I(n410), .Z(n409) );
  BUFFD0 U409 ( .I(n411), .Z(n410) );
  BUFFD0 U410 ( .I(n412), .Z(n411) );
  BUFFD0 U411 ( .I(n413), .Z(n412) );
  BUFFD0 U412 ( .I(n414), .Z(n413) );
  BUFFD0 U413 ( .I(N54), .Z(n414) );
  BUFFD0 U414 ( .I(n426), .Z(n415) );
  INVD1 U415 ( .I(Reset), .ZN(n416) );
  AO222D0 U416 ( .A1(N27), .A2(n417), .B1(N35), .B2(n418), .C1(n300), .C2(n419), .Z(n21) );
  AO222D0 U417 ( .A1(N31), .A2(n417), .B1(N39), .B2(n418), .C1(n182), .C2(n419), .Z(n19) );
  AO222D0 U418 ( .A1(N28), .A2(n417), .B1(N36), .B2(n418), .C1(n240), .C2(n419), .Z(n18) );
  CKND0 U419 ( .CLK(n360), .CN(n419) );
  AN2D0 U420 ( .A1(n420), .A2(n421), .Z(n418) );
  AN3D0 U421 ( .A1(n422), .A2(n423), .A3(n424), .Z(n417) );
  CKXOR2D0 U422 ( .A1(ClockOut), .A2(n425), .Z(n17) );
  AO22D0 U423 ( .A1(N32), .A2(n424), .B1(N40), .B2(n420), .Z(N55) );
  CKND2D0 U424 ( .A1(AdjustFreq[1]), .A2(n421), .ZN(n427) );
  ND3D0 U425 ( .A1(n428), .A2(n423), .A3(n429), .ZN(n421) );
  ND4D0 U426 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(n240), .A4(n300), .ZN(n429) );
  IND3D0 U427 ( .A1(AdjustFreq[1]), .B1(n423), .B2(n422), .ZN(n426) );
  CKND2D0 U428 ( .A1(n182), .A2(DivideFactor[3]), .ZN(n422) );
  AO22D0 U429 ( .A1(N30), .A2(n424), .B1(N38), .B2(n420), .Z(N51) );
  AO22D0 U430 ( .A1(N29), .A2(n424), .B1(N37), .B2(n420), .Z(N49) );
  AN2D0 U431 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n420) );
  NR2D0 U432 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n424) );
  INR2D0 U433 ( .A1(N14), .B1(n425), .ZN(N21) );
  INR2D0 U434 ( .A1(N13), .B1(n425), .ZN(N20) );
  INR2D0 U435 ( .A1(N12), .B1(n425), .ZN(N19) );
  INR2D0 U436 ( .A1(N11), .B1(n425), .ZN(N18) );
  INR2D0 U437 ( .A1(N10), .B1(n425), .ZN(N17) );
  INR2D0 U438 ( .A1(N9), .B1(n425), .ZN(N16) );
  OA21D0 U439 ( .A1(FastDivvy[5]), .A2(n423), .B(n430), .Z(n425) );
  IOA22D0 U440 ( .B1(n431), .B2(n432), .A1(n423), .A2(FastDivvy[5]), .ZN(n430)
         );
  AOI221D0 U441 ( .A1(FastDivvy[4]), .A2(n428), .B1(FastDivvy[3]), .B2(n433), 
        .C(n434), .ZN(n432) );
  AOI221D0 U442 ( .A1(DivideFactor[3]), .A2(n435), .B1(DivideFactor[2]), .B2(
        n436), .C(n437), .ZN(n434) );
  IAO21D0 U443 ( .A1(n436), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n437)
         );
  OAI32D0 U444 ( .A1(n438), .A2(FastDivvy[0]), .A3(n439), .B1(FastDivvy[1]), 
        .B2(n440), .ZN(n436) );
  AN2D0 U445 ( .A1(FastDivvy[1]), .A2(n440), .Z(n439) );
  CKND0 U446 ( .CLK(FastDivvy[3]), .CN(n435) );
  NR2D0 U447 ( .A1(FastDivvy[4]), .A2(n428), .ZN(n431) );
  CKND0 U448 ( .CLK(DivideFactor[5]), .CN(n423) );
  CKND0 U449 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U450 ( .A1(WireD[5]), .A2(n416), .ZN(WireD[0]) );
endmodule


module MultiCounter_0 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [3:0] Ctr;

  MultiCounter_0_DW01_inc_0 add_16 ( .A({CarryOut, n10, n5, n1, n6}), .SUM({N5, 
        N4, N3, N2, N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n11), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n11), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n11), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n11), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n11), .Q(CarryOut) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(Ctr[1]), .Z(n4) );
  BUFFD0 U7 ( .I(Ctr[2]), .Z(n5) );
  BUFFD0 U8 ( .I(n7), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(Ctr[0]), .Z(n9) );
  BUFFD0 U12 ( .I(Ctr[3]), .Z(n10) );
  INVD1 U13 ( .I(Reset), .ZN(n11) );
endmodule


module FIFOTop_AWid3_DWid32_1 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4;
  wire   [2:0] SM_ReadAddr;
  wire   [2:0] SM_WriteAddr;

  FIFOStateM_AWid3_1 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(n1), .ClkW(ClkW), .Reset(n3) );
  DPMem1kx32_AWid3_DWid32_1 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(n1), .ClkW(ClkW), .ChipEna(
        \*Logic1* ), .Read(n2), .Write(SM_MemWriteCmd), .Reset(n3) );
  BUFFD0 U2 ( .I(ClkR), .Z(n1) );
  INVD1 U3 ( .I(n4), .ZN(n3) );
  INVD1 U4 ( .I(Reseter), .ZN(n4) );
  BUFFD1 U5 ( .I(SM_MemReadCmd), .Z(n2) );
  TIEH U6 ( .Z(\*Logic1* ) );
endmodule


module SerEncoder_DWid32_1 ( SerOut, SerValid, FIFO_ReadReq, ParIn, F_Empty, 
        ParClk, SerClk, ParValid, Reset );
  input [31:0] ParIn;
  input F_Empty, ParClk, SerClk, ParValid, Reset;
  output SerOut, SerValid, FIFO_ReadReq;
  wire   N2, N3, N4, N5, N6, HalfParClkr, \Sh_N[5] , N8, N9, N10, N11, N12,
         N13, N23, N24, N25, N26, N27, N28, N29, N31, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88;
  wire   [31:0] InBuf;

  SerEncoder_DWid32_1_DW01_dec_0 \ShifterBlock/sub_132  ( .A({n32, n49, n43, 
        n34, n46, n45}), .SUM({N13, N12, N11, N10, N9, N8}) );
  DFCNQD1 SerValidr_reg ( .D(n63), .CP(n23), .CDN(n70), .Q(SerValid) );
  DFCNQD1 HalfParClkr_reg ( .D(n6), .CP(ParClk), .CDN(n68), .Q(HalfParClkr) );
  DFCNQD1 \InBuf_reg[30]  ( .D(N83), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[30]) );
  DFCNQD1 \InBuf_reg[29]  ( .D(N82), .CP(n23), .CDN(n68), .Q(InBuf[29]) );
  DFCNQD1 \InBuf_reg[26]  ( .D(N79), .CP(n23), .CDN(n69), .Q(InBuf[26]) );
  DFCNQD1 \InBuf_reg[25]  ( .D(N78), .CP(n23), .CDN(n69), .Q(InBuf[25]) );
  DFCNQD1 \InBuf_reg[22]  ( .D(N75), .CP(n65), .CDN(n69), .Q(InBuf[22]) );
  DFCNQD1 \InBuf_reg[21]  ( .D(N74), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[21]) );
  DFCNQD1 \InBuf_reg[18]  ( .D(N71), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[18]) );
  DFCNQD1 \InBuf_reg[17]  ( .D(N70), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[17]) );
  DFCNQD1 \InBuf_reg[14]  ( .D(N67), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[14]) );
  DFCNQD1 \InBuf_reg[13]  ( .D(N66), .CP(n65), .CDN(n70), .Q(InBuf[13]) );
  DFCNQD1 \InBuf_reg[10]  ( .D(N63), .CP(n23), .CDN(n70), .Q(InBuf[10]) );
  DFCNQD1 \InBuf_reg[9]  ( .D(N62), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[9])
         );
  DFCNQD1 \InBuf_reg[6]  ( .D(N59), .CP(n23), .CDN(n69), .Q(InBuf[6]) );
  DFCNQD1 \InBuf_reg[5]  ( .D(N58), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[5])
         );
  DFCNQD1 \InBuf_reg[2]  ( .D(N55), .CP(n23), .CDN(n69), .Q(InBuf[2]) );
  DFCNQD1 \InBuf_reg[1]  ( .D(N54), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[1])
         );
  DFCNQD1 \InBuf_reg[31]  ( .D(N84), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[31]) );
  DFCNQD1 \InBuf_reg[28]  ( .D(N81), .CP(n23), .CDN(n69), .Q(InBuf[28]) );
  DFCNQD1 \InBuf_reg[27]  ( .D(N80), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[27]) );
  DFCNQD1 \InBuf_reg[24]  ( .D(N77), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[24]) );
  DFCNQD1 \InBuf_reg[23]  ( .D(N76), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[23]) );
  DFCNQD1 \InBuf_reg[20]  ( .D(N73), .CP(n23), .CDN(n69), .Q(InBuf[20]) );
  DFCNQD1 \InBuf_reg[19]  ( .D(N72), .CP(n23), .CDN(n69), .Q(InBuf[19]) );
  DFCNQD1 \InBuf_reg[16]  ( .D(N69), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[16]) );
  DFCNQD1 \InBuf_reg[15]  ( .D(N68), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[15]) );
  DFCNQD1 \InBuf_reg[12]  ( .D(N65), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[12]) );
  DFCNQD1 \InBuf_reg[11]  ( .D(N64), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[11]) );
  DFCNQD1 \InBuf_reg[8]  ( .D(N61), .CP(HalfParClkr), .CDN(n68), .Q(InBuf[8])
         );
  DFCNQD1 \InBuf_reg[7]  ( .D(N60), .CP(n23), .CDN(n69), .Q(InBuf[7]) );
  DFCNQD1 \InBuf_reg[4]  ( .D(N57), .CP(HalfParClkr), .CDN(n70), .Q(InBuf[4])
         );
  DFCNQD1 \InBuf_reg[3]  ( .D(N56), .CP(n23), .CDN(n68), .Q(InBuf[3]) );
  DFCNQD1 \InBuf_reg[0]  ( .D(N53), .CP(HalfParClkr), .CDN(n69), .Q(InBuf[0])
         );
  DFCNQD1 \Sh_N_reg[5]  ( .D(N13), .CP(SerClk), .CDN(n68), .Q(\Sh_N[5] ) );
  DFCNQD1 \Sh_N_reg[4]  ( .D(N12), .CP(SerClk), .CDN(n68), .Q(N6) );
  DFCNQD1 \Sh_N_reg[2]  ( .D(N10), .CP(SerClk), .CDN(n68), .Q(N4) );
  DFCNQD1 \Sh_N_reg[3]  ( .D(N11), .CP(SerClk), .CDN(n68), .Q(N5) );
  DFCNQD1 \Sh_N_reg[1]  ( .D(N9), .CP(SerClk), .CDN(n68), .Q(N3) );
  DFCNQD1 \Sh_N_reg[0]  ( .D(N8), .CP(SerClk), .CDN(n68), .Q(N2) );
  DFCNQD1 SerOutr_reg ( .D(n42), .CP(SerClk), .CDN(n70), .Q(SerOut) );
  INR2D1 U3 ( .A1(ParValid), .B1(F_Empty), .ZN(N85) );
  CKND0 U4 ( .CLK(n29), .CN(n67) );
  MUX2ND0 U5 ( .I0(n57), .I1(n58), .S(n48), .ZN(n1) );
  MUX2ND0 U6 ( .I0(n53), .I1(n54), .S(n48), .ZN(n2) );
  MUX2ND0 U7 ( .I0(n55), .I1(n56), .S(n48), .ZN(n3) );
  MUX2ND0 U8 ( .I0(n51), .I1(n52), .S(n48), .ZN(n4) );
  CKBD0 U9 ( .CLK(HalfParClkr), .C(n23) );
  BUFFD0 U10 ( .I(n65), .Z(n5) );
  BUFFD0 U11 ( .I(n8), .Z(n6) );
  BUFFD0 U12 ( .I(n5), .Z(n7) );
  BUFFD0 U13 ( .I(n10), .Z(n8) );
  BUFFD0 U14 ( .I(n7), .Z(n9) );
  BUFFD0 U15 ( .I(n11), .Z(n10) );
  BUFFD0 U16 ( .I(n13), .Z(n11) );
  BUFFD0 U17 ( .I(n9), .Z(n12) );
  BUFFD0 U18 ( .I(n15), .Z(n13) );
  BUFFD0 U19 ( .I(n12), .Z(n14) );
  BUFFD0 U20 ( .I(n17), .Z(n15) );
  BUFFD0 U21 ( .I(n14), .Z(n16) );
  BUFFD0 U22 ( .I(n21), .Z(n17) );
  BUFFD0 U23 ( .I(n16), .Z(n18) );
  BUFFD0 U24 ( .I(n67), .Z(n19) );
  BUFFD0 U25 ( .I(n18), .Z(n20) );
  BUFFD0 U26 ( .I(n24), .Z(n21) );
  BUFFD0 U27 ( .I(n20), .Z(n22) );
  BUFFD0 U28 ( .I(n30), .Z(n24) );
  BUFFD0 U29 ( .I(n23), .Z(n25) );
  BUFFD0 U30 ( .I(n25), .Z(n26) );
  BUFFD0 U31 ( .I(n26), .Z(n27) );
  BUFFD0 U32 ( .I(n27), .Z(n28) );
  BUFFD0 U33 ( .I(n22), .Z(n29) );
  BUFFD0 U34 ( .I(n19), .Z(n30) );
  CKBD0 U35 ( .CLK(\Sh_N[5] ), .C(n31) );
  BUFFD0 U36 ( .I(n44), .Z(n32) );
  BUFFD0 U37 ( .I(N6), .Z(n33) );
  CKBD0 U38 ( .CLK(n50), .C(n43) );
  CKBXD0 U39 ( .I(N5), .Z(n50) );
  BUFFD0 U40 ( .I(n48), .Z(n34) );
  CKBXD0 U41 ( .I(N4), .Z(n48) );
  CKBD0 U42 ( .CLK(N3), .C(n35) );
  CKBD0 U43 ( .CLK(n35), .C(n36) );
  CKBD0 U44 ( .CLK(n36), .C(n37) );
  CKBD0 U45 ( .CLK(N2), .C(n38) );
  CKBD0 U46 ( .CLK(n38), .C(n39) );
  CKBD0 U47 ( .CLK(n39), .C(n40) );
  CKBD0 U48 ( .CLK(n40), .C(n41) );
  BUFFD0 U49 ( .I(N31), .Z(n42) );
  CKBD0 U50 ( .CLK(n37), .C(n46) );
  CKBD0 U51 ( .CLK(n47), .C(n44) );
  CKBXD0 U52 ( .I(n31), .Z(n47) );
  CKBD0 U53 ( .CLK(n41), .C(n45) );
  OR2D0 U54 ( .A1(n45), .A2(n46), .Z(n72) );
  CKND2D0 U55 ( .A1(n46), .A2(n45), .ZN(n73) );
  CKBXD0 U56 ( .I(n33), .Z(n49) );
  INVD1 U57 ( .I(Reset), .ZN(n70) );
  INVD1 U58 ( .I(Reset), .ZN(n69) );
  INVD1 U59 ( .I(Reset), .ZN(n68) );
  INVD1 U60 ( .I(n64), .ZN(n63) );
  INVD1 U61 ( .I(n72), .ZN(n71) );
  AN2D1 U62 ( .A1(n48), .A2(n71), .Z(N26) );
  MUX4ND0 U63 ( .I0(InBuf[8]), .I1(InBuf[9]), .I2(InBuf[10]), .I3(InBuf[11]), 
        .S0(N2), .S1(N3), .ZN(n51) );
  MUX4ND0 U64 ( .I0(InBuf[12]), .I1(InBuf[13]), .I2(InBuf[14]), .I3(InBuf[15]), 
        .S0(N2), .S1(N3), .ZN(n52) );
  MUX4ND0 U65 ( .I0(InBuf[16]), .I1(InBuf[17]), .I2(InBuf[18]), .I3(InBuf[19]), 
        .S0(N2), .S1(N3), .ZN(n53) );
  MUX4ND0 U66 ( .I0(InBuf[20]), .I1(InBuf[21]), .I2(InBuf[22]), .I3(InBuf[23]), 
        .S0(N2), .S1(N3), .ZN(n54) );
  MUX4ND0 U67 ( .I0(InBuf[24]), .I1(InBuf[25]), .I2(InBuf[26]), .I3(InBuf[27]), 
        .S0(N2), .S1(N3), .ZN(n55) );
  MUX4ND0 U68 ( .I0(InBuf[28]), .I1(InBuf[29]), .I2(InBuf[30]), .I3(InBuf[31]), 
        .S0(N2), .S1(N3), .ZN(n56) );
  MUX4ND0 U69 ( .I0(InBuf[0]), .I1(InBuf[1]), .I2(InBuf[2]), .I3(InBuf[3]), 
        .S0(N2), .S1(N3), .ZN(n57) );
  MUX4ND0 U70 ( .I0(InBuf[4]), .I1(InBuf[5]), .I2(InBuf[6]), .I3(InBuf[7]), 
        .S0(N2), .S1(N3), .ZN(n58) );
  NR2D1 U71 ( .A1(n73), .A2(n48), .ZN(N24) );
  INVD1 U72 ( .I(N85), .ZN(n64) );
  INVD1 U73 ( .I(n66), .ZN(n65) );
  INVD1 U74 ( .I(n28), .ZN(n66) );
  MUX2ND0 U75 ( .I0(n59), .I1(n60), .S(n49), .ZN(N29) );
  MUX2ND0 U76 ( .I0(n61), .I1(n62), .S(n49), .ZN(N27) );
  MUX2ND0 U77 ( .I0(n60), .I1(n59), .S(n49), .ZN(N25) );
  MUX2ND0 U78 ( .I0(n62), .I1(n61), .S(n49), .ZN(N23) );
  MUX2ND0 U79 ( .I0(n2), .I1(n3), .S(n50), .ZN(n60) );
  MUX2ND0 U80 ( .I0(n1), .I1(n4), .S(n50), .ZN(n59) );
  MUX2ND0 U81 ( .I0(n3), .I1(n1), .S(n50), .ZN(n62) );
  MUX2ND0 U82 ( .I0(n4), .I1(n2), .S(n50), .ZN(n61) );
  MUX2ND0 U83 ( .I0(n73), .I1(n72), .S(n48), .ZN(N28) );
  AN2D0 U84 ( .A1(ParIn[31]), .A2(N85), .Z(N84) );
  AN2D0 U85 ( .A1(ParIn[30]), .A2(n63), .Z(N83) );
  AN2D0 U86 ( .A1(ParIn[29]), .A2(N85), .Z(N82) );
  AN2D0 U87 ( .A1(ParIn[28]), .A2(n63), .Z(N81) );
  AN2D0 U88 ( .A1(ParIn[27]), .A2(N85), .Z(N80) );
  AN2D0 U89 ( .A1(ParIn[26]), .A2(N85), .Z(N79) );
  AN2D0 U90 ( .A1(ParIn[25]), .A2(N85), .Z(N78) );
  AN2D0 U91 ( .A1(ParIn[24]), .A2(N85), .Z(N77) );
  AN2D0 U92 ( .A1(ParIn[23]), .A2(n63), .Z(N76) );
  AN2D0 U93 ( .A1(ParIn[22]), .A2(n63), .Z(N75) );
  AN2D0 U94 ( .A1(ParIn[21]), .A2(n63), .Z(N74) );
  AN2D0 U95 ( .A1(ParIn[20]), .A2(n63), .Z(N73) );
  AN2D0 U96 ( .A1(ParIn[19]), .A2(n63), .Z(N72) );
  AN2D0 U97 ( .A1(ParIn[18]), .A2(n63), .Z(N71) );
  AN2D0 U98 ( .A1(ParIn[17]), .A2(n63), .Z(N70) );
  AN2D0 U99 ( .A1(ParIn[16]), .A2(N85), .Z(N69) );
  AN2D0 U100 ( .A1(ParIn[15]), .A2(N85), .Z(N68) );
  AN2D0 U101 ( .A1(ParIn[14]), .A2(N85), .Z(N67) );
  AN2D0 U102 ( .A1(ParIn[13]), .A2(N85), .Z(N66) );
  AN2D0 U103 ( .A1(ParIn[12]), .A2(N85), .Z(N65) );
  AN2D0 U104 ( .A1(ParIn[11]), .A2(N85), .Z(N64) );
  AN2D0 U105 ( .A1(ParIn[10]), .A2(n63), .Z(N63) );
  AN2D0 U106 ( .A1(ParIn[9]), .A2(N85), .Z(N62) );
  AN2D0 U107 ( .A1(ParIn[8]), .A2(N85), .Z(N61) );
  AN2D0 U108 ( .A1(ParIn[7]), .A2(n63), .Z(N60) );
  AN2D0 U109 ( .A1(ParIn[6]), .A2(n63), .Z(N59) );
  AN2D0 U110 ( .A1(ParIn[5]), .A2(n63), .Z(N58) );
  AN2D0 U111 ( .A1(ParIn[4]), .A2(n63), .Z(N57) );
  AN2D0 U112 ( .A1(ParIn[3]), .A2(n63), .Z(N56) );
  AN2D0 U113 ( .A1(ParIn[2]), .A2(n63), .Z(N55) );
  AN2D0 U114 ( .A1(ParIn[1]), .A2(n63), .Z(N54) );
  AN2D0 U115 ( .A1(ParIn[0]), .A2(n63), .Z(N53) );
  IND2D0 U116 ( .A1(n74), .B1(n75), .ZN(N31) );
  OAI21D0 U117 ( .A1(N23), .A2(n76), .B(n77), .ZN(n75) );
  MUX2ND0 U118 ( .I0(n78), .I1(n79), .S(n76), .ZN(n77) );
  MUX3ND0 U119 ( .I0(N25), .I1(n80), .I2(N24), .S0(n44), .S1(n81), .ZN(n79) );
  NR2D0 U120 ( .A1(n44), .A2(n50), .ZN(n81) );
  MUX2D0 U121 ( .I0(n82), .I1(N26), .S(n83), .Z(n80) );
  NR2D0 U122 ( .A1(n49), .A2(n50), .ZN(n83) );
  INR2D0 U123 ( .A1(N27), .B1(n49), .ZN(n82) );
  CKND0 U124 ( .CLK(n43), .CN(n78) );
  CKND2D0 U125 ( .A1(n84), .A2(n85), .ZN(n76) );
  MUX2ND0 U126 ( .I0(n86), .I1(n87), .S(n43), .ZN(n74) );
  CKND2D0 U127 ( .A1(N29), .A2(n88), .ZN(n87) );
  CKND2D0 U128 ( .A1(N28), .A2(n88), .ZN(n86) );
  NR2D0 U129 ( .A1(n85), .A2(n84), .ZN(n88) );
  CKND0 U130 ( .CLK(n49), .CN(n84) );
  CKND0 U131 ( .CLK(n44), .CN(n85) );
  INR3D0 U132 ( .A1(n63), .B1(Reset), .B2(n30), .ZN(FIFO_ReadReq) );
endmodule


module SerialTx_1 ( SerOut, SerClk, SerIn, ParClk, Reset );
  input SerIn, ParClk, Reset;
  output SerOut, SerClk;
  wire   n2;

  PLLTop_2 PLL_TxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerIn), .Z(SerOut) );
endmodule


module FIFOTop_AWid4_DWid32_1 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [3:0] SM_ReadAddr;
  wire   [3:0] SM_WriteAddr;

  FIFOStateM_AWid4_1 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid4_DWid32_1 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  CKBD0 U2 ( .CLK(SM_MemReadCmd), .C(n1) );
  INVD1 U3 ( .I(n3), .ZN(n2) );
  INVD1 U4 ( .I(Reseter), .ZN(n3) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32_1 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   SerClock, N30, N31, N32, N33, N34, N37, N38, N39, N40, N41, N42, N43,
         N47, n1, n4, n5, n30, n31, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9026, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294;
  wire   [3:0] ParValidTimer;
  wire   [31:0] Decoder;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  MOAI22D1 U29 ( .A1(n9128), .A2(n9256), .B1(n9129), .B2(Decoder[19]), .ZN(
        n9219) );
  MOAI22D1 U36 ( .A1(n9127), .A2(n9249), .B1(n9129), .B2(Decoder[12]), .ZN(
        n9212) );
  OR3D1 U92 ( .A1(n8152), .A2(n8561), .A3(n8211), .Z(n9276) );
  OR3D1 U94 ( .A1(n8550), .A2(n8359), .A3(n8299), .Z(n9275) );
  OR3D1 U96 ( .A1(n8808), .A2(n8162), .A3(n8009), .Z(n9274) );
  OA21D1 U99 ( .A1(n9272), .A2(n9271), .B(SerValid), .Z(N43) );
  OR2D1 U101 ( .A1(Count32[1]), .A2(Count32[0]), .Z(n9270) );
  DesDecoder_DWid32_1_DW01_inc_0 \ClkGen/add_206  ( .A({Count32[4:2], n6969, 
        n6977}), .SUM({N34, N33, N32, N31, N30}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(n4), .CPN(n9149), .CDN(n9159), .Q(FrameSR[63]) );
  DFNCND1 \FrameSR_reg[22]  ( .D(n30), .CPN(n9154), .CDN(n9159), .Q(
        FrameSR[22]) );
  DFNCND1 \FrameSR_reg[23]  ( .D(n233), .CPN(n9154), .CDN(n9159), .Q(
        FrameSR[23]) );
  DFNCND1 \FrameSR_reg[37]  ( .D(n333), .CPN(n9152), .CDN(n9160), .Q(
        FrameSR[37]) );
  DFNCND1 \FrameSR_reg[38]  ( .D(n432), .CPN(n9152), .CDN(n9160), .Q(
        FrameSR[38]) );
  DFNCND1 \FrameSR_reg[53]  ( .D(n532), .CPN(n9150), .CDN(n9163), .Q(
        FrameSR[53]) );
  DFNCND1 \FrameSR_reg[54]  ( .D(n631), .CPN(n9150), .CDN(n9161), .Q(
        FrameSR[54]) );
  DFNCND1 \FrameSR_reg[32]  ( .D(n731), .CPN(n9153), .CDN(n9160), .Q(
        FrameSR[32]) );
  DFNCND1 \FrameSR_reg[39]  ( .D(n733), .CPN(n9152), .CDN(n9160), .Q(
        FrameSR[39]) );
  DFNCND1 \FrameSR_reg[55]  ( .D(n833), .CPN(n9150), .CDN(n9161), .Q(
        FrameSR[55]) );
  DFNCND1 \FrameSR_reg[8]  ( .D(n933), .CPN(n9155), .CDN(n9157), .Q(FrameSR[8]) );
  DFNCND1 \FrameSR_reg[9]  ( .D(n937), .CPN(n9155), .CDN(n9157), .Q(FrameSR[9]) );
  DFNCND1 \FrameSR_reg[10]  ( .D(n939), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[10]) );
  DFNCND1 \FrameSR_reg[11]  ( .D(n941), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[11]) );
  DFNCND1 \FrameSR_reg[12]  ( .D(n943), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[12]) );
  DFNCND1 \FrameSR_reg[13]  ( .D(n945), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[13]) );
  DFNCND1 \FrameSR_reg[14]  ( .D(n947), .CPN(n9155), .CDN(n9158), .Q(
        FrameSR[14]) );
  DFNCND1 \FrameSR_reg[15]  ( .D(n949), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[15]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(n951), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[19]) );
  DFNCND1 \FrameSR_reg[24]  ( .D(n1050), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[24]) );
  DFNCND1 \FrameSR_reg[25]  ( .D(n1150), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[25]) );
  DFNCND1 \FrameSR_reg[26]  ( .D(n1152), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[26]) );
  DFNCND1 \FrameSR_reg[27]  ( .D(n1154), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[27]) );
  DFNCND1 \FrameSR_reg[28]  ( .D(n1156), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[28]) );
  DFNCND1 \FrameSR_reg[29]  ( .D(n1158), .CPN(n9153), .CDN(n9159), .Q(
        FrameSR[29]) );
  DFNCND1 \FrameSR_reg[30]  ( .D(n1160), .CPN(n9153), .CDN(n9160), .Q(
        FrameSR[30]) );
  DFNCND1 \FrameSR_reg[31]  ( .D(n1162), .CPN(n9153), .CDN(n9160), .Q(
        FrameSR[31]) );
  DFNCND1 \FrameSR_reg[40]  ( .D(n1164), .CPN(n9152), .CDN(n9158), .Q(
        FrameSR[40]) );
  DFNCND1 \FrameSR_reg[41]  ( .D(n1264), .CPN(n9152), .CDN(n9161), .Q(
        FrameSR[41]) );
  DFNCND1 \FrameSR_reg[42]  ( .D(n1266), .CPN(n9151), .CDN(n9163), .Q(
        FrameSR[42]) );
  DFNCND1 \FrameSR_reg[43]  ( .D(n1268), .CPN(n9151), .CDN(n9163), .Q(
        FrameSR[43]) );
  DFNCND1 \FrameSR_reg[44]  ( .D(n1270), .CPN(n9151), .CDN(n9163), .Q(
        FrameSR[44]) );
  DFNCND1 \FrameSR_reg[45]  ( .D(n1272), .CPN(n9151), .CDN(n9164), .Q(
        FrameSR[45]) );
  DFNCND1 \FrameSR_reg[46]  ( .D(n1274), .CPN(n9151), .CDN(n9159), .Q(
        FrameSR[46]) );
  DFNCND1 \FrameSR_reg[47]  ( .D(n1276), .CPN(n9151), .CDN(n9163), .Q(
        FrameSR[47]) );
  DFNCND1 \FrameSR_reg[56]  ( .D(n1278), .CPN(n9150), .CDN(n9163), .Q(
        FrameSR[56]) );
  DFNCND1 \FrameSR_reg[57]  ( .D(n1378), .CPN(n9150), .CDN(n9164), .Q(
        FrameSR[57]) );
  DFNCND1 \FrameSR_reg[58]  ( .D(n1380), .CPN(n9150), .CDN(n9157), .Q(
        FrameSR[58]) );
  DFNCND1 \FrameSR_reg[59]  ( .D(n1382), .CPN(n9150), .CDN(n9163), .Q(
        FrameSR[59]) );
  DFNCND1 \FrameSR_reg[60]  ( .D(n1384), .CPN(n9149), .CDN(n9162), .Q(
        FrameSR[60]) );
  DFNCND1 \FrameSR_reg[61]  ( .D(n1386), .CPN(n9149), .CDN(n9161), .Q(
        FrameSR[61]) );
  DFNCND1 \FrameSR_reg[62]  ( .D(n1388), .CPN(n9149), .CDN(n9164), .Q(
        FrameSR[62]) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[0]) );
  DFNCND1 \FrameSR_reg[4]  ( .D(n1390), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(n1393), .CPN(n9154), .CDN(n9159), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(n1492), .CPN(n9152), .CDN(n9160), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(n1591), .CPN(n9151), .CDN(n9162), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(n1690), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(n1693), .CPN(n9155), .CDN(n9157), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(n1697), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(n1796), .CPN(n9152), .CDN(n9160), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(n1896), .CPN(n9151), .CDN(n9161), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(n1898), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(n1901), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(n1904), .CPN(n9156), .CDN(n9157), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(n1907), .CPN(n9155), .CDN(n9157), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(n1911), .CPN(n9154), .CDN(n9159), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(n2010), .CPN(n9152), .CDN(n9160), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(n2109), .CPN(n9151), .CDN(n9162), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[51]  ( .D(n2208), .CPN(n9150), .CDN(n9161), .Q(
        FrameSR[51]) );
  DFNCND1 \FrameSR_reg[36]  ( .D(n2307), .CPN(n9152), .CDN(n9160), .Q(
        FrameSR[36]) );
  DFNCND1 \FrameSR_reg[52]  ( .D(n2406), .CPN(n9150), .CDN(n9157), .Q(
        FrameSR[52]) );
  DFNCND1 \FrameSR_reg[17]  ( .D(n2505), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[17]) );
  DFNCND1 \FrameSR_reg[16]  ( .D(n2604), .CPN(n9154), .CDN(n9158), .Q(
        FrameSR[16]) );
  EDFCNQD1 \Count32_reg[4]  ( .D(n2606), .E(SerValid), .CP(n9141), .CDN(n9160), 
        .Q(Count32[4]) );
  DFNCND1 \Decoder_reg[31]  ( .D(n2607), .CPN(n9149), .CDN(n9160), .Q(
        Decoder[31]) );
  DFNCND1 \Decoder_reg[30]  ( .D(n2741), .CPN(n9149), .CDN(n9159), .Q(
        Decoder[30]) );
  DFNCND1 \Decoder_reg[29]  ( .D(n2877), .CPN(n9149), .CDN(n9159), .Q(
        Decoder[29]) );
  DFNCND1 \Decoder_reg[28]  ( .D(n3013), .CPN(n9149), .CDN(n9158), .Q(
        Decoder[28]) );
  DFNCND1 \Decoder_reg[27]  ( .D(n3149), .CPN(n9149), .CDN(n9158), .Q(
        Decoder[27]) );
  DFNCND1 \Decoder_reg[26]  ( .D(n3285), .CPN(n9148), .CDN(n9157), .Q(
        Decoder[26]) );
  DFNCND1 \Decoder_reg[25]  ( .D(n3421), .CPN(n9148), .CDN(n9162), .Q(
        Decoder[25]) );
  DFNCND1 \Decoder_reg[24]  ( .D(n3557), .CPN(n9148), .CDN(n9163), .Q(
        Decoder[24]) );
  DFNCND1 \Decoder_reg[23]  ( .D(n3693), .CPN(n9148), .CDN(n9162), .Q(
        Decoder[23]) );
  DFNCND1 \Decoder_reg[22]  ( .D(n3829), .CPN(n9148), .CDN(n9161), .Q(
        Decoder[22]) );
  DFNCND1 \Decoder_reg[21]  ( .D(n3965), .CPN(n9148), .CDN(n9161), .Q(
        Decoder[21]) );
  DFNCND1 \Decoder_reg[20]  ( .D(n4101), .CPN(n9148), .CDN(n9160), .Q(
        Decoder[20]) );
  DFNCND1 \Decoder_reg[19]  ( .D(n4237), .CPN(n9148), .CDN(n9164), .Q(
        Decoder[19]) );
  DFNCND1 \Decoder_reg[18]  ( .D(n4374), .CPN(n9148), .CDN(n9157), .Q(
        Decoder[18]) );
  DFNCND1 \Decoder_reg[17]  ( .D(n4510), .CPN(n9147), .CDN(n9160), .Q(
        Decoder[17]) );
  DFNCND1 \Decoder_reg[16]  ( .D(n4646), .CPN(n9147), .CDN(n9159), .Q(
        Decoder[16]) );
  DFNCND1 \Decoder_reg[15]  ( .D(n4782), .CPN(n9147), .CDN(n9157), .Q(
        Decoder[15]) );
  DFNCND1 \Decoder_reg[14]  ( .D(n4918), .CPN(n9147), .CDN(n9158), .Q(
        Decoder[14]) );
  DFNCND1 \Decoder_reg[13]  ( .D(n5054), .CPN(n9147), .CDN(n9158), .Q(
        Decoder[13]) );
  DFNCND1 \Decoder_reg[12]  ( .D(n5191), .CPN(n9147), .CDN(n9163), .Q(
        Decoder[12]) );
  DFNCND1 \Decoder_reg[11]  ( .D(n5327), .CPN(n9147), .CDN(n9161), .Q(
        Decoder[11]) );
  DFNCND1 \Decoder_reg[10]  ( .D(n5463), .CPN(n9147), .CDN(n9162), .Q(
        Decoder[10]) );
  DFNCND1 \Decoder_reg[9]  ( .D(n5599), .CPN(n9147), .CDN(n9162), .Q(
        Decoder[9]) );
  DFNCND1 \Decoder_reg[8]  ( .D(n5735), .CPN(n9146), .CDN(n9162), .Q(
        Decoder[8]) );
  DFNCND1 \Decoder_reg[7]  ( .D(n5871), .CPN(n9146), .CDN(n9160), .Q(
        Decoder[7]) );
  DFNCND1 \Decoder_reg[6]  ( .D(n6007), .CPN(n9146), .CDN(n9164), .Q(
        Decoder[6]) );
  DFNCND1 \Decoder_reg[5]  ( .D(n6144), .CPN(n9146), .CDN(n9157), .Q(
        Decoder[5]) );
  DFNCND1 \Decoder_reg[4]  ( .D(n6281), .CPN(n9146), .CDN(n9160), .Q(
        Decoder[4]) );
  DFNCND1 \Decoder_reg[3]  ( .D(n6418), .CPN(n9146), .CDN(n9164), .Q(
        Decoder[3]) );
  DFNCND1 \Decoder_reg[2]  ( .D(n6555), .CPN(n9146), .CDN(n9163), .Q(
        Decoder[2]) );
  DFNCND1 \Decoder_reg[1]  ( .D(n6692), .CPN(n9146), .CDN(n9162), .Q(
        Decoder[1]) );
  DFNCND1 \Decoder_reg[0]  ( .D(n6829), .CPN(n9146), .CDN(n9161), .Q(
        Decoder[0]) );
  DFNCND1 \ParValidTimer_reg[1]  ( .D(n6966), .CPN(n9142), .CDN(n9162), .Q(
        ParValidTimer[1]) );
  EDFCNQD1 \Count32_reg[1]  ( .D(n6968), .E(SerValid), .CP(n9141), .CDN(n9163), 
        .Q(Count32[1]) );
  DFNCND1 \ParValidTimer_reg[0]  ( .D(n6970), .CPN(n9142), .CDN(n9162), .Q(
        ParValidTimer[0]) );
  EDFCNQD1 \Count32_reg[3]  ( .D(n6972), .E(SerValid), .CP(n9141), .CDN(n9161), 
        .Q(Count32[3]) );
  EDFCNQD1 \Count32_reg[2]  ( .D(n6974), .E(SerValid), .CP(n9141), .CDN(n9160), 
        .Q(Count32[2]) );
  EDFCNQD1 \Count32_reg[0]  ( .D(n6976), .E(SerValid), .CP(n9141), .CDN(n9161), 
        .Q(Count32[0]) );
  DFNCND1 \ParOutr_reg[2]  ( .D(n6978), .CPN(n9145), .CDN(n9163), .Q(ParOut[2]), .QN(n9239) );
  DFNCND1 \ParOutr_reg[1]  ( .D(n6982), .CPN(n9145), .CDN(n9163), .Q(ParOut[1]), .QN(n9238) );
  EDFCNQD1 ParClkr_reg ( .D(n6986), .E(n6988), .CP(n9141), .CDN(n9164), .Q(
        ParClk) );
  DFNCND1 \ParOutr_reg[0]  ( .D(n6990), .CPN(n9145), .CDN(n9158), .Q(ParOut[0]), .QN(n9237) );
  DFNCND1 \ParOutr_reg[5]  ( .D(n6994), .CPN(n9145), .CDN(n9159), .Q(ParOut[5]), .QN(n9242) );
  DFNCND1 \ParOutr_reg[12]  ( .D(n6998), .CPN(n9144), .CDN(n9164), .Q(
        ParOut[12]), .QN(n9249) );
  DFNCND1 \ParOutr_reg[19]  ( .D(n7002), .CPN(n9143), .CDN(n9157), .Q(
        ParOut[19]), .QN(n9256) );
  DFNCND1 \ParOutr_reg[6]  ( .D(n7006), .CPN(n9145), .CDN(n9163), .Q(ParOut[6]), .QN(n9243) );
  DFNCND1 \ParOutr_reg[9]  ( .D(n7010), .CPN(n9144), .CDN(n9162), .Q(ParOut[9]), .QN(n9246) );
  DFNCND1 \ParOutr_reg[13]  ( .D(n7014), .CPN(n9144), .CDN(n9158), .Q(
        ParOut[13]), .QN(n9250) );
  DFNCND1 \ParOutr_reg[16]  ( .D(n7018), .CPN(n9143), .CDN(n9163), .Q(
        ParOut[16]), .QN(n9253) );
  DFNCND1 \ParOutr_reg[20]  ( .D(n7022), .CPN(n9143), .CDN(n9162), .Q(
        ParOut[20]), .QN(n9257) );
  DFNCND1 \ParOutr_reg[23]  ( .D(n7026), .CPN(n9143), .CDN(n9162), .Q(
        ParOut[23]), .QN(n9260) );
  DFNCND1 \ParOutr_reg[24]  ( .D(n7030), .CPN(n9143), .CDN(n9164), .Q(
        ParOut[24]), .QN(n9261) );
  DFNCND1 \ParOutr_reg[27]  ( .D(n7034), .CPN(n9142), .CDN(n9162), .Q(
        ParOut[27]), .QN(n9264) );
  DFNCND1 \ParOutr_reg[28]  ( .D(n7038), .CPN(n9142), .CDN(n9164), .Q(
        ParOut[28]), .QN(n9265) );
  DFNCND1 \ParOutr_reg[31]  ( .D(n7042), .CPN(n9142), .CDN(n9161), .Q(
        ParOut[31]), .QN(n9268) );
  DFNCND1 \ParOutr_reg[3]  ( .D(n7046), .CPN(n9145), .CDN(n9161), .Q(ParOut[3]), .QN(n9240) );
  DFNCND1 \ParOutr_reg[4]  ( .D(n7050), .CPN(n9145), .CDN(n9164), .Q(ParOut[4]), .QN(n9241) );
  DFNCND1 \ParOutr_reg[10]  ( .D(n7054), .CPN(n9144), .CDN(n9164), .Q(
        ParOut[10]), .QN(n9247) );
  DFNCND1 \ParOutr_reg[11]  ( .D(n7058), .CPN(n9144), .CDN(n9164), .Q(
        ParOut[11]), .QN(n9248) );
  DFNCND1 \ParOutr_reg[17]  ( .D(n7062), .CPN(n9143), .CDN(n9161), .Q(
        ParOut[17]), .QN(n9254) );
  DFNCND1 \ParOutr_reg[18]  ( .D(n7066), .CPN(n9143), .CDN(n9161), .Q(
        ParOut[18]), .QN(n9255) );
  DFNCND1 \ParOutr_reg[7]  ( .D(n7070), .CPN(n9144), .CDN(n9163), .Q(ParOut[7]), .QN(n9244) );
  DFNCND1 \ParOutr_reg[8]  ( .D(n7074), .CPN(n9144), .CDN(n9159), .Q(ParOut[8]), .QN(n9245) );
  DFNCND1 \ParOutr_reg[14]  ( .D(n7078), .CPN(n9144), .CDN(n9159), .Q(
        ParOut[14]), .QN(n9251) );
  DFNCND1 \ParOutr_reg[15]  ( .D(n7082), .CPN(n9144), .CDN(n9162), .Q(
        ParOut[15]), .QN(n9252) );
  DFNCND1 \ParOutr_reg[21]  ( .D(n7086), .CPN(n9143), .CDN(n9160), .Q(
        ParOut[21]), .QN(n9258) );
  DFNCND1 \ParOutr_reg[22]  ( .D(n7090), .CPN(n9143), .CDN(n9162), .Q(
        ParOut[22]), .QN(n9259) );
  DFNCND1 \ParOutr_reg[25]  ( .D(n7094), .CPN(n9142), .CDN(n9157), .Q(
        ParOut[25]), .QN(n9262) );
  DFNCND1 \ParOutr_reg[26]  ( .D(n7098), .CPN(n9142), .CDN(n9164), .Q(
        ParOut[26]), .QN(n9263) );
  DFNCND1 \ParOutr_reg[29]  ( .D(n7102), .CPN(n9142), .CDN(n9161), .Q(
        ParOut[29]), .QN(n9266) );
  DFNCND1 \ParOutr_reg[30]  ( .D(n7106), .CPN(n9142), .CDN(n9163), .Q(
        ParOut[30]), .QN(n9267) );
  DFNCND1 ParValidr_reg ( .D(n7110), .CPN(n9141), .CDN(n9158), .Q(ParValid), 
        .QN(n9269) );
  DFNCND1 doParSync_reg ( .D(N47), .CPN(n9145), .CDN(n9164), .Q(n9271), .QN(
        n9294) );
  DFNCND1 UnLoad_reg ( .D(n9017), .CPN(n9145), .CDN(n9164), .Q(n1), .QN(n9166)
         );
  DFNCND1 \ParValidTimer_reg[3]  ( .D(n9018), .CPN(n9141), .CDN(n9164), .QN(
        n9165) );
  DFNCND1 \ParValidTimer_reg[2]  ( .D(n9021), .CPN(n9141), .CDN(n9164), .QN(
        n9167) );
  IOA22D0 U3 ( .B1(n9128), .B2(n9268), .A1(n1), .A2(Decoder[31]), .ZN(n9231)
         );
  AO22D0 U4 ( .A1(n6143), .A2(n9017), .B1(Decoder[6]), .B2(n9126), .Z(n9193)
         );
  CKAN2D0 U5 ( .A1(N30), .A2(n9294), .Z(N38) );
  INVD0 U6 ( .I(ParValidTimer[0]), .ZN(n9292) );
  BUFFD0 U7 ( .I(n2876), .Z(n4) );
  CKBD0 U8 ( .CLK(FrameSR[62]), .C(n5) );
  BUFFD0 U9 ( .I(n8197), .Z(n30) );
  CKBD0 U10 ( .CLK(FrameSR[21]), .C(n31) );
  CKBD0 U11 ( .CLK(n31), .C(n64) );
  CKBD0 U12 ( .CLK(n64), .C(n65) );
  CKBD0 U13 ( .CLK(n65), .C(n66) );
  CKBD0 U14 ( .CLK(n66), .C(n67) );
  CKBD0 U15 ( .CLK(n67), .C(n68) );
  CKBD0 U16 ( .CLK(n68), .C(n69) );
  CKBD0 U17 ( .CLK(n69), .C(n70) );
  CKBD0 U18 ( .CLK(n70), .C(n71) );
  CKBD0 U19 ( .CLK(n71), .C(n72) );
  BUFFD0 U20 ( .I(n72), .Z(n73) );
  CKBD0 U21 ( .CLK(n73), .C(n74) );
  CKBD0 U22 ( .CLK(n74), .C(n75) );
  CKBD0 U23 ( .CLK(n75), .C(n76) );
  CKBD0 U24 ( .CLK(n76), .C(n77) );
  CKBD0 U25 ( .CLK(n77), .C(n78) );
  CKBD0 U26 ( .CLK(n78), .C(n79) );
  CKBD0 U27 ( .CLK(n79), .C(n80) );
  CKBD0 U28 ( .CLK(n80), .C(n81) );
  CKBD0 U30 ( .CLK(n81), .C(n82) );
  CKBD0 U31 ( .CLK(n82), .C(n83) );
  BUFFD0 U32 ( .I(n83), .Z(n84) );
  CKBD0 U33 ( .CLK(n84), .C(n85) );
  CKBD0 U34 ( .CLK(n85), .C(n86) );
  CKBD0 U35 ( .CLK(n86), .C(n87) );
  CKBD0 U37 ( .CLK(n87), .C(n88) );
  CKBD0 U38 ( .CLK(n88), .C(n89) );
  CKBD0 U39 ( .CLK(n89), .C(n90) );
  CKBD0 U40 ( .CLK(n90), .C(n91) );
  CKBD0 U41 ( .CLK(n91), .C(n92) );
  CKBD0 U42 ( .CLK(n92), .C(n93) );
  CKBD0 U43 ( .CLK(n93), .C(n94) );
  BUFFD0 U44 ( .I(n94), .Z(n95) );
  CKBD0 U45 ( .CLK(n95), .C(n165) );
  CKBD0 U46 ( .CLK(n165), .C(n166) );
  CKBD0 U47 ( .CLK(n166), .C(n167) );
  CKBD0 U48 ( .CLK(n167), .C(n168) );
  CKBD0 U49 ( .CLK(n168), .C(n169) );
  CKBD0 U50 ( .CLK(n169), .C(n170) );
  CKBD0 U51 ( .CLK(n170), .C(n171) );
  CKBD0 U52 ( .CLK(n171), .C(n172) );
  CKBD0 U53 ( .CLK(n172), .C(n173) );
  CKBD0 U54 ( .CLK(n173), .C(n174) );
  BUFFD0 U55 ( .I(n174), .Z(n175) );
  CKBD0 U56 ( .CLK(n175), .C(n176) );
  CKBD0 U57 ( .CLK(n176), .C(n177) );
  CKBD0 U58 ( .CLK(n177), .C(n178) );
  CKBD0 U59 ( .CLK(n178), .C(n179) );
  CKBD0 U60 ( .CLK(n179), .C(n180) );
  CKBD0 U61 ( .CLK(n180), .C(n181) );
  CKBD0 U62 ( .CLK(n181), .C(n182) );
  CKBD0 U63 ( .CLK(n182), .C(n183) );
  CKBD0 U64 ( .CLK(n183), .C(n184) );
  CKBD0 U65 ( .CLK(n184), .C(n185) );
  BUFFD0 U66 ( .I(n185), .Z(n186) );
  CKBD0 U67 ( .CLK(n186), .C(n187) );
  CKBD0 U68 ( .CLK(n187), .C(n188) );
  CKBD0 U69 ( .CLK(n188), .C(n189) );
  CKBD0 U70 ( .CLK(n189), .C(n190) );
  CKBD0 U71 ( .CLK(n190), .C(n191) );
  CKBD0 U72 ( .CLK(n191), .C(n192) );
  CKBD0 U73 ( .CLK(n192), .C(n193) );
  CKBD0 U74 ( .CLK(n193), .C(n194) );
  CKBD0 U75 ( .CLK(n194), .C(n195) );
  BUFFD0 U76 ( .I(n195), .Z(n196) );
  CKBD0 U77 ( .CLK(n196), .C(n197) );
  CKBD0 U78 ( .CLK(n197), .C(n198) );
  CKBD0 U79 ( .CLK(n198), .C(n199) );
  CKBD0 U80 ( .CLK(n199), .C(n200) );
  CKBD0 U81 ( .CLK(n200), .C(n201) );
  CKBD0 U82 ( .CLK(n201), .C(n202) );
  CKBD0 U83 ( .CLK(n202), .C(n203) );
  CKBD0 U84 ( .CLK(n203), .C(n204) );
  CKBD0 U85 ( .CLK(n204), .C(n205) );
  CKBD0 U86 ( .CLK(n205), .C(n206) );
  BUFFD0 U87 ( .I(n206), .Z(n207) );
  CKBD0 U88 ( .CLK(n207), .C(n208) );
  CKBD0 U89 ( .CLK(n208), .C(n209) );
  CKBD0 U90 ( .CLK(n209), .C(n210) );
  CKBD0 U91 ( .CLK(n210), .C(n211) );
  CKBD0 U93 ( .CLK(n211), .C(n212) );
  CKBD0 U95 ( .CLK(n212), .C(n213) );
  CKBD0 U97 ( .CLK(n213), .C(n214) );
  CKBD0 U98 ( .CLK(n214), .C(n215) );
  CKBD0 U100 ( .CLK(n215), .C(n216) );
  CKBD0 U102 ( .CLK(n216), .C(n217) );
  BUFFD0 U103 ( .I(n217), .Z(n218) );
  CKBD0 U104 ( .CLK(n218), .C(n219) );
  CKBD0 U105 ( .CLK(n219), .C(n220) );
  CKBD0 U106 ( .CLK(n220), .C(n221) );
  CKBD0 U107 ( .CLK(n221), .C(n222) );
  CKBD0 U108 ( .CLK(n222), .C(n223) );
  CKBD0 U109 ( .CLK(n223), .C(n224) );
  CKBD0 U110 ( .CLK(n224), .C(n225) );
  CKBD0 U111 ( .CLK(n225), .C(n226) );
  CKBD0 U112 ( .CLK(n226), .C(n227) );
  CKBD0 U113 ( .CLK(n227), .C(n228) );
  CKBD0 U114 ( .CLK(n228), .C(n229) );
  BUFFD0 U115 ( .I(n8009), .Z(n233) );
  CKBD0 U116 ( .CLK(FrameSR[22]), .C(n234) );
  CKBD0 U117 ( .CLK(n234), .C(n235) );
  CKBD0 U118 ( .CLK(n235), .C(n236) );
  CKBD0 U119 ( .CLK(n236), .C(n237) );
  CKBD0 U120 ( .CLK(n237), .C(n238) );
  BUFFD0 U121 ( .I(n238), .Z(n239) );
  CKBD0 U122 ( .CLK(n239), .C(n240) );
  CKBD0 U123 ( .CLK(n240), .C(n241) );
  CKBD0 U124 ( .CLK(n241), .C(n242) );
  CKBD0 U125 ( .CLK(n242), .C(n243) );
  CKBD0 U126 ( .CLK(n243), .C(n244) );
  CKBD0 U127 ( .CLK(n244), .C(n245) );
  CKBD0 U128 ( .CLK(n245), .C(n246) );
  CKBD0 U129 ( .CLK(n246), .C(n247) );
  CKBD0 U130 ( .CLK(n247), .C(n248) );
  CKBD0 U131 ( .CLK(n248), .C(n249) );
  BUFFD0 U132 ( .I(n249), .Z(n250) );
  CKBD0 U133 ( .CLK(n250), .C(n251) );
  CKBD0 U134 ( .CLK(n251), .C(n252) );
  CKBD0 U135 ( .CLK(n252), .C(n253) );
  CKBD0 U136 ( .CLK(n253), .C(n254) );
  CKBD0 U137 ( .CLK(n254), .C(n255) );
  CKBD0 U138 ( .CLK(n255), .C(n256) );
  CKBD0 U139 ( .CLK(n256), .C(n257) );
  CKBD0 U140 ( .CLK(n257), .C(n258) );
  CKBD0 U141 ( .CLK(n258), .C(n259) );
  CKBD0 U142 ( .CLK(n259), .C(n260) );
  BUFFD0 U143 ( .I(n260), .Z(n261) );
  CKBD0 U144 ( .CLK(n261), .C(n262) );
  CKBD0 U145 ( .CLK(n262), .C(n263) );
  CKBD0 U146 ( .CLK(n263), .C(n264) );
  CKBD0 U147 ( .CLK(n264), .C(n265) );
  CKBD0 U148 ( .CLK(n265), .C(n266) );
  CKBD0 U149 ( .CLK(n266), .C(n267) );
  CKBD0 U150 ( .CLK(n267), .C(n268) );
  CKBD0 U151 ( .CLK(n268), .C(n269) );
  CKBD0 U152 ( .CLK(n269), .C(n270) );
  CKBD0 U153 ( .CLK(n270), .C(n271) );
  BUFFD0 U154 ( .I(n271), .Z(n272) );
  CKBD0 U155 ( .CLK(n272), .C(n273) );
  CKBD0 U156 ( .CLK(n273), .C(n274) );
  CKBD0 U157 ( .CLK(n274), .C(n275) );
  CKBD0 U158 ( .CLK(n275), .C(n276) );
  CKBD0 U159 ( .CLK(n276), .C(n277) );
  CKBD0 U160 ( .CLK(n277), .C(n278) );
  CKBD0 U161 ( .CLK(n278), .C(n279) );
  CKBD0 U162 ( .CLK(n279), .C(n280) );
  CKBD0 U163 ( .CLK(n280), .C(n281) );
  CKBD0 U164 ( .CLK(n281), .C(n282) );
  BUFFD0 U165 ( .I(n282), .Z(n283) );
  CKBD0 U166 ( .CLK(n283), .C(n284) );
  CKBD0 U167 ( .CLK(n284), .C(n285) );
  CKBD0 U168 ( .CLK(n285), .C(n286) );
  CKBD0 U169 ( .CLK(n286), .C(n287) );
  CKBD0 U170 ( .CLK(n287), .C(n288) );
  CKBD0 U171 ( .CLK(n288), .C(n289) );
  CKBD0 U172 ( .CLK(n289), .C(n290) );
  CKBD0 U173 ( .CLK(n290), .C(n291) );
  CKBD0 U174 ( .CLK(n291), .C(n292) );
  BUFFD0 U175 ( .I(n292), .Z(n293) );
  CKBD0 U176 ( .CLK(n293), .C(n294) );
  CKBD0 U177 ( .CLK(n294), .C(n295) );
  CKBD0 U178 ( .CLK(n295), .C(n296) );
  CKBD0 U179 ( .CLK(n296), .C(n297) );
  CKBD0 U180 ( .CLK(n297), .C(n298) );
  CKBD0 U181 ( .CLK(n298), .C(n299) );
  CKBD0 U182 ( .CLK(n299), .C(n300) );
  CKBD0 U183 ( .CLK(n300), .C(n301) );
  CKBD0 U184 ( .CLK(n301), .C(n302) );
  CKBD0 U185 ( .CLK(n302), .C(n303) );
  BUFFD0 U186 ( .I(n303), .Z(n304) );
  CKBD0 U187 ( .CLK(n304), .C(n305) );
  CKBD0 U188 ( .CLK(n305), .C(n306) );
  CKBD0 U189 ( .CLK(n306), .C(n307) );
  CKBD0 U190 ( .CLK(n307), .C(n308) );
  CKBD0 U191 ( .CLK(n308), .C(n309) );
  CKBD0 U192 ( .CLK(n309), .C(n310) );
  CKBD0 U193 ( .CLK(n310), .C(n311) );
  CKBD0 U194 ( .CLK(n311), .C(n312) );
  CKBD0 U195 ( .CLK(n312), .C(n313) );
  CKBD0 U196 ( .CLK(n313), .C(n314) );
  BUFFD0 U197 ( .I(n314), .Z(n315) );
  CKBD0 U198 ( .CLK(n315), .C(n316) );
  CKBD0 U199 ( .CLK(n316), .C(n317) );
  CKBD0 U200 ( .CLK(n317), .C(n318) );
  CKBD0 U201 ( .CLK(n318), .C(n319) );
  CKBD0 U202 ( .CLK(n319), .C(n320) );
  CKBD0 U203 ( .CLK(n320), .C(n321) );
  CKBD0 U204 ( .CLK(n321), .C(n322) );
  CKBD0 U205 ( .CLK(n322), .C(n323) );
  CKBD0 U206 ( .CLK(n323), .C(n324) );
  CKBD0 U207 ( .CLK(n324), .C(n325) );
  BUFFD0 U208 ( .I(n325), .Z(n326) );
  CKBD0 U209 ( .CLK(n326), .C(n327) );
  CKBD0 U210 ( .CLK(n327), .C(n328) );
  CKBD0 U211 ( .CLK(n328), .C(n329) );
  CKBD0 U212 ( .CLK(n329), .C(n330) );
  CKBD0 U213 ( .CLK(n330), .C(n331) );
  CKBD0 U214 ( .CLK(n331), .C(n332) );
  BUFFD0 U215 ( .I(n8892), .Z(n333) );
  CKBD0 U216 ( .CLK(FrameSR[36]), .C(n334) );
  BUFFD0 U217 ( .I(n334), .Z(n335) );
  CKBD0 U218 ( .CLK(n335), .C(n336) );
  CKBD0 U219 ( .CLK(n336), .C(n337) );
  CKBD0 U220 ( .CLK(n337), .C(n338) );
  CKBD0 U221 ( .CLK(n338), .C(n339) );
  CKBD0 U222 ( .CLK(n339), .C(n340) );
  CKBD0 U223 ( .CLK(n340), .C(n341) );
  CKBD0 U224 ( .CLK(n341), .C(n342) );
  CKBD0 U225 ( .CLK(n342), .C(n343) );
  CKBD0 U226 ( .CLK(n343), .C(n344) );
  CKBD0 U227 ( .CLK(n344), .C(n345) );
  BUFFD0 U228 ( .I(n345), .Z(n346) );
  CKBD0 U229 ( .CLK(n346), .C(n347) );
  CKBD0 U230 ( .CLK(n347), .C(n348) );
  CKBD0 U231 ( .CLK(n348), .C(n349) );
  CKBD0 U232 ( .CLK(n349), .C(n350) );
  CKBD0 U233 ( .CLK(n350), .C(n351) );
  CKBD0 U234 ( .CLK(n351), .C(n352) );
  CKBD0 U235 ( .CLK(n352), .C(n353) );
  CKBD0 U236 ( .CLK(n353), .C(n354) );
  CKBD0 U237 ( .CLK(n354), .C(n355) );
  CKBD0 U238 ( .CLK(n355), .C(n356) );
  BUFFD0 U239 ( .I(n356), .Z(n357) );
  CKBD0 U240 ( .CLK(n357), .C(n358) );
  CKBD0 U241 ( .CLK(n358), .C(n359) );
  CKBD0 U242 ( .CLK(n359), .C(n360) );
  CKBD0 U243 ( .CLK(n360), .C(n361) );
  CKBD0 U244 ( .CLK(n361), .C(n362) );
  CKBD0 U245 ( .CLK(n362), .C(n363) );
  CKBD0 U246 ( .CLK(n363), .C(n364) );
  CKBD0 U247 ( .CLK(n364), .C(n365) );
  CKBD0 U248 ( .CLK(n365), .C(n366) );
  CKBD0 U249 ( .CLK(n366), .C(n367) );
  BUFFD0 U250 ( .I(n367), .Z(n368) );
  CKBD0 U251 ( .CLK(n368), .C(n369) );
  CKBD0 U252 ( .CLK(n369), .C(n370) );
  CKBD0 U253 ( .CLK(n370), .C(n371) );
  CKBD0 U254 ( .CLK(n371), .C(n372) );
  CKBD0 U255 ( .CLK(n372), .C(n373) );
  CKBD0 U256 ( .CLK(n373), .C(n374) );
  CKBD0 U257 ( .CLK(n374), .C(n375) );
  CKBD0 U258 ( .CLK(n375), .C(n376) );
  CKBD0 U259 ( .CLK(n376), .C(n377) );
  CKBD0 U260 ( .CLK(n377), .C(n378) );
  BUFFD0 U261 ( .I(n378), .Z(n379) );
  CKBD0 U262 ( .CLK(n379), .C(n380) );
  CKBD0 U263 ( .CLK(n380), .C(n381) );
  CKBD0 U264 ( .CLK(n381), .C(n382) );
  CKBD0 U265 ( .CLK(n382), .C(n383) );
  CKBD0 U266 ( .CLK(n383), .C(n384) );
  CKBD0 U267 ( .CLK(n384), .C(n385) );
  CKBD0 U268 ( .CLK(n385), .C(n386) );
  CKBD0 U269 ( .CLK(n386), .C(n387) );
  CKBD0 U270 ( .CLK(n387), .C(n388) );
  BUFFD0 U271 ( .I(n388), .Z(n389) );
  CKBD0 U272 ( .CLK(n389), .C(n390) );
  CKBD0 U273 ( .CLK(n390), .C(n391) );
  CKBD0 U274 ( .CLK(n391), .C(n392) );
  CKBD0 U275 ( .CLK(n392), .C(n393) );
  CKBD0 U276 ( .CLK(n393), .C(n394) );
  CKBD0 U277 ( .CLK(n394), .C(n395) );
  CKBD0 U278 ( .CLK(n395), .C(n396) );
  CKBD0 U279 ( .CLK(n396), .C(n397) );
  CKBD0 U280 ( .CLK(n397), .C(n398) );
  CKBD0 U281 ( .CLK(n398), .C(n399) );
  BUFFD0 U282 ( .I(n399), .Z(n400) );
  CKBD0 U283 ( .CLK(n400), .C(n401) );
  CKBD0 U284 ( .CLK(n401), .C(n402) );
  CKBD0 U285 ( .CLK(n402), .C(n403) );
  CKBD0 U286 ( .CLK(n403), .C(n404) );
  CKBD0 U287 ( .CLK(n404), .C(n405) );
  CKBD0 U288 ( .CLK(n405), .C(n406) );
  CKBD0 U289 ( .CLK(n406), .C(n407) );
  CKBD0 U290 ( .CLK(n407), .C(n408) );
  CKBD0 U291 ( .CLK(n408), .C(n409) );
  CKBD0 U292 ( .CLK(n409), .C(n410) );
  BUFFD0 U293 ( .I(n410), .Z(n411) );
  CKBD0 U294 ( .CLK(n411), .C(n412) );
  CKBD0 U295 ( .CLK(n412), .C(n413) );
  CKBD0 U296 ( .CLK(n413), .C(n414) );
  CKBD0 U297 ( .CLK(n414), .C(n415) );
  CKBD0 U298 ( .CLK(n415), .C(n416) );
  CKBD0 U299 ( .CLK(n416), .C(n417) );
  CKBD0 U300 ( .CLK(n417), .C(n418) );
  CKBD0 U301 ( .CLK(n418), .C(n419) );
  CKBD0 U302 ( .CLK(n419), .C(n420) );
  CKBD0 U303 ( .CLK(n420), .C(n421) );
  BUFFD0 U304 ( .I(n421), .Z(n422) );
  CKBD0 U305 ( .CLK(n422), .C(n423) );
  CKBD0 U306 ( .CLK(n423), .C(n424) );
  CKBD0 U307 ( .CLK(n424), .C(n425) );
  CKBD0 U308 ( .CLK(n425), .C(n426) );
  CKBD0 U309 ( .CLK(n426), .C(n427) );
  CKBD0 U310 ( .CLK(n427), .C(n428) );
  CKBD0 U311 ( .CLK(n428), .C(n429) );
  CKBD0 U312 ( .CLK(n429), .C(n430) );
  BUFFD0 U313 ( .I(n430), .Z(n431) );
  BUFFD0 U314 ( .I(n8299), .Z(n432) );
  CKBD0 U315 ( .CLK(FrameSR[37]), .C(n433) );
  CKBD0 U316 ( .CLK(n433), .C(n434) );
  CKBD0 U317 ( .CLK(n434), .C(n435) );
  CKBD0 U318 ( .CLK(n435), .C(n436) );
  CKBD0 U319 ( .CLK(n436), .C(n437) );
  CKBD0 U320 ( .CLK(n437), .C(n438) );
  CKBD0 U321 ( .CLK(n438), .C(n439) );
  CKBD0 U322 ( .CLK(n439), .C(n440) );
  CKBD0 U323 ( .CLK(n440), .C(n441) );
  BUFFD0 U324 ( .I(n441), .Z(n442) );
  CKBD0 U325 ( .CLK(n442), .C(n443) );
  CKBD0 U326 ( .CLK(n443), .C(n444) );
  CKBD0 U327 ( .CLK(n444), .C(n445) );
  CKBD0 U328 ( .CLK(n445), .C(n446) );
  CKBD0 U329 ( .CLK(n446), .C(n447) );
  CKBD0 U330 ( .CLK(n447), .C(n448) );
  CKBD0 U331 ( .CLK(n448), .C(n449) );
  CKBD0 U332 ( .CLK(n449), .C(n450) );
  CKBD0 U333 ( .CLK(n450), .C(n451) );
  CKBD0 U334 ( .CLK(n451), .C(n452) );
  BUFFD0 U335 ( .I(n452), .Z(n453) );
  CKBD0 U336 ( .CLK(n453), .C(n454) );
  CKBD0 U337 ( .CLK(n454), .C(n455) );
  CKBD0 U338 ( .CLK(n455), .C(n456) );
  CKBD0 U339 ( .CLK(n456), .C(n457) );
  CKBD0 U340 ( .CLK(n457), .C(n458) );
  CKBD0 U341 ( .CLK(n458), .C(n459) );
  CKBD0 U342 ( .CLK(n459), .C(n460) );
  CKBD0 U343 ( .CLK(n460), .C(n461) );
  CKBD0 U344 ( .CLK(n461), .C(n462) );
  CKBD0 U345 ( .CLK(n462), .C(n463) );
  BUFFD0 U346 ( .I(n463), .Z(n464) );
  CKBD0 U347 ( .CLK(n464), .C(n465) );
  CKBD0 U348 ( .CLK(n465), .C(n466) );
  CKBD0 U349 ( .CLK(n466), .C(n467) );
  CKBD0 U350 ( .CLK(n467), .C(n468) );
  CKBD0 U351 ( .CLK(n468), .C(n469) );
  CKBD0 U352 ( .CLK(n469), .C(n470) );
  CKBD0 U353 ( .CLK(n470), .C(n471) );
  CKBD0 U354 ( .CLK(n471), .C(n472) );
  CKBD0 U355 ( .CLK(n472), .C(n473) );
  CKBD0 U356 ( .CLK(n473), .C(n474) );
  BUFFD0 U357 ( .I(n474), .Z(n475) );
  CKBD0 U358 ( .CLK(n475), .C(n476) );
  CKBD0 U359 ( .CLK(n476), .C(n477) );
  CKBD0 U360 ( .CLK(n477), .C(n478) );
  CKBD0 U361 ( .CLK(n478), .C(n479) );
  CKBD0 U362 ( .CLK(n479), .C(n480) );
  CKBD0 U363 ( .CLK(n480), .C(n481) );
  CKBD0 U364 ( .CLK(n481), .C(n482) );
  CKBD0 U365 ( .CLK(n482), .C(n483) );
  CKBD0 U366 ( .CLK(n483), .C(n484) );
  CKBD0 U367 ( .CLK(n484), .C(n485) );
  BUFFD0 U368 ( .I(n485), .Z(n486) );
  CKBD0 U369 ( .CLK(n486), .C(n487) );
  CKBD0 U370 ( .CLK(n487), .C(n488) );
  CKBD0 U371 ( .CLK(n488), .C(n489) );
  CKBD0 U372 ( .CLK(n489), .C(n490) );
  CKBD0 U373 ( .CLK(n490), .C(n491) );
  CKBD0 U374 ( .CLK(n491), .C(n492) );
  CKBD0 U375 ( .CLK(n492), .C(n493) );
  CKBD0 U376 ( .CLK(n493), .C(n494) );
  CKBD0 U377 ( .CLK(n494), .C(n495) );
  CKBD0 U378 ( .CLK(n495), .C(n496) );
  BUFFD0 U379 ( .I(n496), .Z(n497) );
  CKBD0 U380 ( .CLK(n497), .C(n498) );
  CKBD0 U381 ( .CLK(n498), .C(n499) );
  CKBD0 U382 ( .CLK(n499), .C(n500) );
  CKBD0 U383 ( .CLK(n500), .C(n501) );
  CKBD0 U384 ( .CLK(n501), .C(n502) );
  CKBD0 U385 ( .CLK(n502), .C(n503) );
  CKBD0 U386 ( .CLK(n503), .C(n504) );
  CKBD0 U387 ( .CLK(n504), .C(n505) );
  CKBD0 U388 ( .CLK(n505), .C(n506) );
  BUFFD0 U389 ( .I(n506), .Z(n507) );
  CKBD0 U390 ( .CLK(n507), .C(n508) );
  CKBD0 U391 ( .CLK(n508), .C(n509) );
  CKBD0 U392 ( .CLK(n509), .C(n510) );
  CKBD0 U393 ( .CLK(n510), .C(n511) );
  CKBD0 U394 ( .CLK(n511), .C(n512) );
  CKBD0 U395 ( .CLK(n512), .C(n513) );
  CKBD0 U396 ( .CLK(n513), .C(n514) );
  CKBD0 U397 ( .CLK(n514), .C(n515) );
  CKBD0 U398 ( .CLK(n515), .C(n516) );
  CKBD0 U399 ( .CLK(n516), .C(n517) );
  BUFFD0 U400 ( .I(n517), .Z(n518) );
  CKBD0 U401 ( .CLK(n518), .C(n519) );
  CKBD0 U402 ( .CLK(n519), .C(n520) );
  CKBD0 U403 ( .CLK(n520), .C(n521) );
  CKBD0 U404 ( .CLK(n521), .C(n522) );
  CKBD0 U405 ( .CLK(n522), .C(n523) );
  CKBD0 U406 ( .CLK(n523), .C(n524) );
  CKBD0 U407 ( .CLK(n524), .C(n525) );
  CKBD0 U408 ( .CLK(n525), .C(n526) );
  CKBD0 U409 ( .CLK(n526), .C(n527) );
  CKBD0 U410 ( .CLK(n527), .C(n528) );
  BUFFD0 U411 ( .I(n528), .Z(n529) );
  CKBD0 U412 ( .CLK(n529), .C(n530) );
  CKBD0 U413 ( .CLK(n530), .C(n531) );
  BUFFD0 U414 ( .I(n8224), .Z(n532) );
  CKBD0 U415 ( .CLK(FrameSR[52]), .C(n533) );
  CKBD0 U416 ( .CLK(n533), .C(n534) );
  CKBD0 U417 ( .CLK(n534), .C(n535) );
  CKBD0 U418 ( .CLK(n535), .C(n536) );
  CKBD0 U419 ( .CLK(n536), .C(n537) );
  CKBD0 U420 ( .CLK(n537), .C(n538) );
  CKBD0 U421 ( .CLK(n538), .C(n539) );
  CKBD0 U422 ( .CLK(n539), .C(n540) );
  BUFFD0 U423 ( .I(n540), .Z(n541) );
  CKBD0 U424 ( .CLK(n541), .C(n542) );
  CKBD0 U425 ( .CLK(n542), .C(n543) );
  CKBD0 U426 ( .CLK(n543), .C(n544) );
  CKBD0 U427 ( .CLK(n544), .C(n545) );
  CKBD0 U428 ( .CLK(n545), .C(n546) );
  CKBD0 U429 ( .CLK(n546), .C(n547) );
  CKBD0 U430 ( .CLK(n547), .C(n548) );
  CKBD0 U431 ( .CLK(n548), .C(n549) );
  CKBD0 U432 ( .CLK(n549), .C(n550) );
  CKBD0 U433 ( .CLK(n550), .C(n551) );
  BUFFD0 U434 ( .I(n551), .Z(n552) );
  CKBD0 U435 ( .CLK(n552), .C(n553) );
  CKBD0 U436 ( .CLK(n553), .C(n554) );
  CKBD0 U437 ( .CLK(n554), .C(n555) );
  CKBD0 U438 ( .CLK(n555), .C(n556) );
  CKBD0 U439 ( .CLK(n556), .C(n557) );
  CKBD0 U440 ( .CLK(n557), .C(n558) );
  CKBD0 U441 ( .CLK(n558), .C(n559) );
  CKBD0 U442 ( .CLK(n559), .C(n560) );
  CKBD0 U443 ( .CLK(n560), .C(n561) );
  BUFFD0 U444 ( .I(n561), .Z(n562) );
  CKBD0 U445 ( .CLK(n562), .C(n563) );
  CKBD0 U446 ( .CLK(n563), .C(n564) );
  CKBD0 U447 ( .CLK(n564), .C(n565) );
  CKBD0 U448 ( .CLK(n565), .C(n566) );
  CKBD0 U449 ( .CLK(n566), .C(n567) );
  CKBD0 U450 ( .CLK(n567), .C(n568) );
  CKBD0 U451 ( .CLK(n568), .C(n569) );
  CKBD0 U452 ( .CLK(n569), .C(n570) );
  CKBD0 U453 ( .CLK(n570), .C(n571) );
  CKBD0 U454 ( .CLK(n571), .C(n572) );
  BUFFD0 U455 ( .I(n572), .Z(n573) );
  CKBD0 U456 ( .CLK(n573), .C(n574) );
  CKBD0 U457 ( .CLK(n574), .C(n575) );
  CKBD0 U458 ( .CLK(n575), .C(n576) );
  CKBD0 U459 ( .CLK(n576), .C(n577) );
  CKBD0 U460 ( .CLK(n577), .C(n578) );
  CKBD0 U461 ( .CLK(n578), .C(n579) );
  CKBD0 U462 ( .CLK(n579), .C(n580) );
  CKBD0 U463 ( .CLK(n580), .C(n581) );
  CKBD0 U464 ( .CLK(n581), .C(n582) );
  CKBD0 U465 ( .CLK(n582), .C(n583) );
  BUFFD0 U466 ( .I(n583), .Z(n584) );
  CKBD0 U467 ( .CLK(n584), .C(n585) );
  CKBD0 U468 ( .CLK(n585), .C(n586) );
  CKBD0 U469 ( .CLK(n586), .C(n587) );
  CKBD0 U470 ( .CLK(n587), .C(n588) );
  CKBD0 U471 ( .CLK(n588), .C(n589) );
  CKBD0 U472 ( .CLK(n589), .C(n590) );
  CKBD0 U473 ( .CLK(n590), .C(n591) );
  CKBD0 U474 ( .CLK(n591), .C(n592) );
  CKBD0 U475 ( .CLK(n592), .C(n593) );
  CKBD0 U476 ( .CLK(n593), .C(n594) );
  BUFFD0 U477 ( .I(n594), .Z(n595) );
  CKBD0 U478 ( .CLK(n595), .C(n596) );
  CKBD0 U479 ( .CLK(n596), .C(n597) );
  CKBD0 U480 ( .CLK(n597), .C(n598) );
  CKBD0 U481 ( .CLK(n598), .C(n599) );
  CKBD0 U482 ( .CLK(n599), .C(n600) );
  CKBD0 U483 ( .CLK(n600), .C(n601) );
  CKBD0 U484 ( .CLK(n601), .C(n602) );
  CKBD0 U485 ( .CLK(n602), .C(n603) );
  CKBD0 U486 ( .CLK(n603), .C(n604) );
  CKBD0 U487 ( .CLK(n604), .C(n605) );
  BUFFD0 U488 ( .I(n605), .Z(n606) );
  CKBD0 U489 ( .CLK(n606), .C(n607) );
  CKBD0 U490 ( .CLK(n607), .C(n608) );
  CKBD0 U491 ( .CLK(n608), .C(n609) );
  CKBD0 U492 ( .CLK(n609), .C(n610) );
  CKBD0 U493 ( .CLK(n610), .C(n611) );
  CKBD0 U494 ( .CLK(n611), .C(n612) );
  CKBD0 U495 ( .CLK(n612), .C(n613) );
  CKBD0 U496 ( .CLK(n613), .C(n614) );
  CKBD0 U497 ( .CLK(n614), .C(n615) );
  CKBD0 U498 ( .CLK(n615), .C(n616) );
  BUFFD0 U499 ( .I(n616), .Z(n617) );
  CKBD0 U500 ( .CLK(n617), .C(n618) );
  CKBD0 U501 ( .CLK(n618), .C(n619) );
  CKBD0 U502 ( .CLK(n619), .C(n620) );
  CKBD0 U503 ( .CLK(n620), .C(n621) );
  CKBD0 U504 ( .CLK(n621), .C(n622) );
  CKBD0 U505 ( .CLK(n622), .C(n623) );
  CKBD0 U506 ( .CLK(n623), .C(n624) );
  CKBD0 U507 ( .CLK(n624), .C(n625) );
  CKBD0 U508 ( .CLK(n625), .C(n626) );
  CKBD0 U509 ( .CLK(n626), .C(n627) );
  BUFFD0 U510 ( .I(n627), .Z(n628) );
  CKBD0 U511 ( .CLK(n628), .C(n629) );
  CKBD0 U512 ( .CLK(n629), .C(n630) );
  BUFFD0 U513 ( .I(n8211), .Z(n631) );
  CKBD0 U514 ( .CLK(FrameSR[53]), .C(n632) );
  BUFFD0 U515 ( .I(n632), .Z(n633) );
  CKBD0 U516 ( .CLK(n633), .C(n634) );
  CKBD0 U517 ( .CLK(n634), .C(n635) );
  CKBD0 U518 ( .CLK(n635), .C(n636) );
  CKBD0 U519 ( .CLK(n636), .C(n637) );
  CKBD0 U520 ( .CLK(n637), .C(n638) );
  CKBD0 U521 ( .CLK(n638), .C(n639) );
  CKBD0 U522 ( .CLK(n639), .C(n640) );
  CKBD0 U523 ( .CLK(n640), .C(n641) );
  CKBD0 U524 ( .CLK(n641), .C(n642) );
  BUFFD0 U525 ( .I(n642), .Z(n643) );
  CKBD0 U526 ( .CLK(n643), .C(n644) );
  CKBD0 U527 ( .CLK(n644), .C(n645) );
  CKBD0 U528 ( .CLK(n645), .C(n646) );
  CKBD0 U529 ( .CLK(n646), .C(n647) );
  CKBD0 U530 ( .CLK(n647), .C(n648) );
  CKBD0 U531 ( .CLK(n648), .C(n649) );
  CKBD0 U532 ( .CLK(n649), .C(n650) );
  CKBD0 U533 ( .CLK(n650), .C(n651) );
  CKBD0 U534 ( .CLK(n651), .C(n652) );
  CKBD0 U535 ( .CLK(n652), .C(n653) );
  BUFFD0 U536 ( .I(n653), .Z(n654) );
  CKBD0 U537 ( .CLK(n654), .C(n655) );
  CKBD0 U538 ( .CLK(n655), .C(n656) );
  CKBD0 U539 ( .CLK(n656), .C(n657) );
  CKBD0 U540 ( .CLK(n657), .C(n658) );
  CKBD0 U541 ( .CLK(n658), .C(n659) );
  CKBD0 U542 ( .CLK(n659), .C(n660) );
  CKBD0 U543 ( .CLK(n660), .C(n661) );
  CKBD0 U544 ( .CLK(n661), .C(n662) );
  CKBD0 U545 ( .CLK(n662), .C(n663) );
  CKBD0 U546 ( .CLK(n663), .C(n664) );
  BUFFD0 U547 ( .I(n664), .Z(n665) );
  CKBD0 U548 ( .CLK(n665), .C(n666) );
  CKBD0 U549 ( .CLK(n666), .C(n667) );
  CKBD0 U550 ( .CLK(n667), .C(n668) );
  CKBD0 U551 ( .CLK(n668), .C(n669) );
  CKBD0 U552 ( .CLK(n669), .C(n670) );
  CKBD0 U553 ( .CLK(n670), .C(n671) );
  CKBD0 U554 ( .CLK(n671), .C(n672) );
  CKBD0 U555 ( .CLK(n672), .C(n673) );
  CKBD0 U556 ( .CLK(n673), .C(n674) );
  CKBD0 U557 ( .CLK(n674), .C(n675) );
  BUFFD0 U558 ( .I(n675), .Z(n676) );
  CKBD0 U559 ( .CLK(n676), .C(n677) );
  CKBD0 U560 ( .CLK(n677), .C(n678) );
  CKBD0 U561 ( .CLK(n678), .C(n679) );
  CKBD0 U562 ( .CLK(n679), .C(n680) );
  CKBD0 U563 ( .CLK(n680), .C(n681) );
  CKBD0 U564 ( .CLK(n681), .C(n682) );
  CKBD0 U565 ( .CLK(n682), .C(n683) );
  CKBD0 U566 ( .CLK(n683), .C(n684) );
  CKBD0 U567 ( .CLK(n684), .C(n685) );
  CKBD0 U568 ( .CLK(n685), .C(n686) );
  BUFFD0 U569 ( .I(n686), .Z(n687) );
  CKBD0 U570 ( .CLK(n687), .C(n688) );
  CKBD0 U571 ( .CLK(n688), .C(n689) );
  CKBD0 U572 ( .CLK(n689), .C(n690) );
  CKBD0 U573 ( .CLK(n690), .C(n691) );
  CKBD0 U574 ( .CLK(n691), .C(n692) );
  CKBD0 U575 ( .CLK(n692), .C(n693) );
  CKBD0 U576 ( .CLK(n693), .C(n694) );
  CKBD0 U577 ( .CLK(n694), .C(n695) );
  CKBD0 U578 ( .CLK(n695), .C(n696) );
  CKBD0 U579 ( .CLK(n696), .C(n697) );
  BUFFD0 U580 ( .I(n697), .Z(n698) );
  CKBD0 U581 ( .CLK(n698), .C(n699) );
  CKBD0 U582 ( .CLK(n699), .C(n700) );
  CKBD0 U583 ( .CLK(n700), .C(n701) );
  CKBD0 U584 ( .CLK(n701), .C(n702) );
  CKBD0 U585 ( .CLK(n702), .C(n703) );
  CKBD0 U586 ( .CLK(n703), .C(n704) );
  CKBD0 U587 ( .CLK(n704), .C(n705) );
  CKBD0 U588 ( .CLK(n705), .C(n706) );
  CKBD0 U589 ( .CLK(n706), .C(n707) );
  CKBD0 U590 ( .CLK(n707), .C(n708) );
  BUFFD0 U591 ( .I(n708), .Z(n709) );
  CKBD0 U592 ( .CLK(n709), .C(n710) );
  CKBD0 U593 ( .CLK(n710), .C(n711) );
  CKBD0 U594 ( .CLK(n711), .C(n712) );
  CKBD0 U595 ( .CLK(n712), .C(n713) );
  CKBD0 U596 ( .CLK(n713), .C(n714) );
  CKBD0 U597 ( .CLK(n714), .C(n715) );
  CKBD0 U598 ( .CLK(n715), .C(n716) );
  CKBD0 U599 ( .CLK(n716), .C(n717) );
  CKBD0 U600 ( .CLK(n717), .C(n718) );
  BUFFD0 U601 ( .I(n718), .Z(n719) );
  CKBD0 U602 ( .CLK(n719), .C(n720) );
  CKBD0 U603 ( .CLK(n720), .C(n721) );
  CKBD0 U604 ( .CLK(n721), .C(n722) );
  CKBD0 U605 ( .CLK(n722), .C(n723) );
  CKBD0 U606 ( .CLK(n723), .C(n724) );
  CKBD0 U607 ( .CLK(n724), .C(n725) );
  CKBD0 U608 ( .CLK(n725), .C(n726) );
  CKBD0 U609 ( .CLK(n726), .C(n727) );
  CKBD0 U610 ( .CLK(n727), .C(n728) );
  CKBD0 U611 ( .CLK(n728), .C(n729) );
  CKBD0 U612 ( .CLK(n729), .C(n730) );
  BUFFD0 U613 ( .I(n4917), .Z(n731) );
  CKBD0 U614 ( .CLK(FrameSR[31]), .C(n732) );
  BUFFD0 U615 ( .I(n8359), .Z(n733) );
  CKBD0 U616 ( .CLK(FrameSR[38]), .C(n734) );
  CKBD0 U617 ( .CLK(n734), .C(n735) );
  CKBD0 U618 ( .CLK(n735), .C(n736) );
  CKBD0 U619 ( .CLK(n736), .C(n737) );
  CKBD0 U620 ( .CLK(n737), .C(n738) );
  CKBD0 U621 ( .CLK(n738), .C(n739) );
  CKBD0 U622 ( .CLK(n739), .C(n740) );
  BUFFD0 U623 ( .I(n740), .Z(n741) );
  CKBD0 U624 ( .CLK(n741), .C(n742) );
  CKBD0 U625 ( .CLK(n742), .C(n743) );
  CKBD0 U626 ( .CLK(n743), .C(n744) );
  CKBD0 U627 ( .CLK(n744), .C(n745) );
  CKBD0 U628 ( .CLK(n745), .C(n746) );
  CKBD0 U629 ( .CLK(n746), .C(n747) );
  CKBD0 U630 ( .CLK(n747), .C(n748) );
  CKBD0 U631 ( .CLK(n748), .C(n749) );
  CKBD0 U632 ( .CLK(n749), .C(n750) );
  CKBD0 U633 ( .CLK(n750), .C(n751) );
  BUFFD0 U634 ( .I(n751), .Z(n752) );
  CKBD0 U635 ( .CLK(n752), .C(n753) );
  CKBD0 U636 ( .CLK(n753), .C(n754) );
  CKBD0 U637 ( .CLK(n754), .C(n755) );
  CKBD0 U638 ( .CLK(n755), .C(n756) );
  CKBD0 U639 ( .CLK(n756), .C(n757) );
  CKBD0 U640 ( .CLK(n757), .C(n758) );
  CKBD0 U641 ( .CLK(n758), .C(n759) );
  CKBD0 U642 ( .CLK(n759), .C(n760) );
  CKBD0 U643 ( .CLK(n760), .C(n761) );
  CKBD0 U644 ( .CLK(n761), .C(n762) );
  BUFFD0 U645 ( .I(n762), .Z(n763) );
  CKBD0 U646 ( .CLK(n763), .C(n764) );
  CKBD0 U647 ( .CLK(n764), .C(n765) );
  CKBD0 U648 ( .CLK(n765), .C(n766) );
  CKBD0 U649 ( .CLK(n766), .C(n767) );
  CKBD0 U650 ( .CLK(n767), .C(n768) );
  CKBD0 U651 ( .CLK(n768), .C(n769) );
  CKBD0 U652 ( .CLK(n769), .C(n770) );
  CKBD0 U653 ( .CLK(n770), .C(n771) );
  CKBD0 U654 ( .CLK(n771), .C(n772) );
  CKBD0 U655 ( .CLK(n772), .C(n773) );
  BUFFD0 U656 ( .I(n773), .Z(n774) );
  CKBD0 U657 ( .CLK(n774), .C(n775) );
  CKBD0 U658 ( .CLK(n775), .C(n776) );
  CKBD0 U659 ( .CLK(n776), .C(n777) );
  CKBD0 U660 ( .CLK(n777), .C(n778) );
  CKBD0 U661 ( .CLK(n778), .C(n779) );
  CKBD0 U662 ( .CLK(n779), .C(n780) );
  CKBD0 U663 ( .CLK(n780), .C(n781) );
  CKBD0 U664 ( .CLK(n781), .C(n782) );
  CKBD0 U665 ( .CLK(n782), .C(n783) );
  CKBD0 U666 ( .CLK(n783), .C(n784) );
  BUFFD0 U667 ( .I(n784), .Z(n785) );
  CKBD0 U668 ( .CLK(n785), .C(n786) );
  CKBD0 U669 ( .CLK(n786), .C(n787) );
  CKBD0 U670 ( .CLK(n787), .C(n788) );
  CKBD0 U671 ( .CLK(n788), .C(n789) );
  CKBD0 U672 ( .CLK(n789), .C(n790) );
  CKBD0 U673 ( .CLK(n790), .C(n791) );
  CKBD0 U674 ( .CLK(n791), .C(n792) );
  CKBD0 U675 ( .CLK(n792), .C(n793) );
  CKBD0 U676 ( .CLK(n793), .C(n794) );
  CKBD0 U677 ( .CLK(n794), .C(n795) );
  BUFFD0 U678 ( .I(n795), .Z(n796) );
  CKBD0 U679 ( .CLK(n796), .C(n797) );
  CKBD0 U680 ( .CLK(n797), .C(n798) );
  CKBD0 U681 ( .CLK(n798), .C(n799) );
  CKBD0 U682 ( .CLK(n799), .C(n800) );
  CKBD0 U683 ( .CLK(n800), .C(n801) );
  CKBD0 U684 ( .CLK(n801), .C(n802) );
  CKBD0 U685 ( .CLK(n802), .C(n803) );
  CKBD0 U686 ( .CLK(n803), .C(n804) );
  CKBD0 U687 ( .CLK(n804), .C(n805) );
  BUFFD0 U688 ( .I(n805), .Z(n806) );
  CKBD0 U689 ( .CLK(n806), .C(n807) );
  CKBD0 U690 ( .CLK(n807), .C(n808) );
  CKBD0 U691 ( .CLK(n808), .C(n809) );
  CKBD0 U692 ( .CLK(n809), .C(n810) );
  CKBD0 U693 ( .CLK(n810), .C(n811) );
  CKBD0 U694 ( .CLK(n811), .C(n812) );
  CKBD0 U695 ( .CLK(n812), .C(n813) );
  CKBD0 U696 ( .CLK(n813), .C(n814) );
  CKBD0 U697 ( .CLK(n814), .C(n815) );
  CKBD0 U698 ( .CLK(n815), .C(n816) );
  BUFFD0 U699 ( .I(n816), .Z(n817) );
  CKBD0 U700 ( .CLK(n817), .C(n818) );
  CKBD0 U701 ( .CLK(n818), .C(n819) );
  CKBD0 U702 ( .CLK(n819), .C(n820) );
  CKBD0 U703 ( .CLK(n820), .C(n821) );
  CKBD0 U704 ( .CLK(n821), .C(n822) );
  CKBD0 U705 ( .CLK(n822), .C(n823) );
  CKBD0 U706 ( .CLK(n823), .C(n824) );
  CKBD0 U707 ( .CLK(n824), .C(n825) );
  CKBD0 U708 ( .CLK(n825), .C(n826) );
  CKBD0 U709 ( .CLK(n826), .C(n827) );
  BUFFD0 U710 ( .I(n827), .Z(n828) );
  CKBD0 U711 ( .CLK(n828), .C(n829) );
  CKBD0 U712 ( .CLK(n829), .C(n830) );
  CKBD0 U713 ( .CLK(n830), .C(n831) );
  CKBD0 U714 ( .CLK(n831), .C(n832) );
  BUFFD0 U715 ( .I(n8561), .Z(n833) );
  CKBD0 U716 ( .CLK(FrameSR[54]), .C(n834) );
  CKBD0 U717 ( .CLK(n834), .C(n835) );
  CKBD0 U718 ( .CLK(n835), .C(n836) );
  CKBD0 U719 ( .CLK(n836), .C(n837) );
  CKBD0 U720 ( .CLK(n837), .C(n838) );
  CKBD0 U721 ( .CLK(n838), .C(n839) );
  CKBD0 U722 ( .CLK(n839), .C(n840) );
  BUFFD0 U723 ( .I(n840), .Z(n841) );
  CKBD0 U724 ( .CLK(n841), .C(n842) );
  CKBD0 U725 ( .CLK(n842), .C(n843) );
  CKBD0 U726 ( .CLK(n843), .C(n844) );
  CKBD0 U727 ( .CLK(n844), .C(n845) );
  CKBD0 U728 ( .CLK(n845), .C(n846) );
  CKBD0 U729 ( .CLK(n846), .C(n847) );
  CKBD0 U730 ( .CLK(n847), .C(n848) );
  CKBD0 U731 ( .CLK(n848), .C(n849) );
  CKBD0 U732 ( .CLK(n849), .C(n850) );
  CKBD0 U733 ( .CLK(n850), .C(n851) );
  BUFFD0 U734 ( .I(n851), .Z(n852) );
  CKBD0 U735 ( .CLK(n852), .C(n853) );
  CKBD0 U736 ( .CLK(n853), .C(n854) );
  CKBD0 U737 ( .CLK(n854), .C(n855) );
  CKBD0 U738 ( .CLK(n855), .C(n856) );
  CKBD0 U739 ( .CLK(n856), .C(n857) );
  CKBD0 U740 ( .CLK(n857), .C(n858) );
  CKBD0 U741 ( .CLK(n858), .C(n859) );
  CKBD0 U742 ( .CLK(n859), .C(n860) );
  CKBD0 U743 ( .CLK(n860), .C(n861) );
  CKBD0 U744 ( .CLK(n861), .C(n862) );
  BUFFD0 U745 ( .I(n862), .Z(n863) );
  CKBD0 U746 ( .CLK(n863), .C(n864) );
  CKBD0 U747 ( .CLK(n864), .C(n865) );
  CKBD0 U748 ( .CLK(n865), .C(n866) );
  CKBD0 U749 ( .CLK(n866), .C(n867) );
  CKBD0 U750 ( .CLK(n867), .C(n868) );
  CKBD0 U751 ( .CLK(n868), .C(n869) );
  CKBD0 U752 ( .CLK(n869), .C(n870) );
  CKBD0 U753 ( .CLK(n870), .C(n871) );
  CKBD0 U754 ( .CLK(n871), .C(n872) );
  CKBD0 U755 ( .CLK(n872), .C(n873) );
  BUFFD0 U756 ( .I(n873), .Z(n874) );
  CKBD0 U757 ( .CLK(n874), .C(n875) );
  CKBD0 U758 ( .CLK(n875), .C(n876) );
  CKBD0 U759 ( .CLK(n876), .C(n877) );
  CKBD0 U760 ( .CLK(n877), .C(n878) );
  CKBD0 U761 ( .CLK(n878), .C(n879) );
  CKBD0 U762 ( .CLK(n879), .C(n880) );
  CKBD0 U763 ( .CLK(n880), .C(n881) );
  CKBD0 U764 ( .CLK(n881), .C(n882) );
  CKBD0 U765 ( .CLK(n882), .C(n883) );
  CKBD0 U766 ( .CLK(n883), .C(n884) );
  BUFFD0 U767 ( .I(n884), .Z(n885) );
  CKBD0 U768 ( .CLK(n885), .C(n886) );
  CKBD0 U769 ( .CLK(n886), .C(n887) );
  CKBD0 U770 ( .CLK(n887), .C(n888) );
  CKBD0 U771 ( .CLK(n888), .C(n889) );
  CKBD0 U772 ( .CLK(n889), .C(n890) );
  CKBD0 U773 ( .CLK(n890), .C(n891) );
  CKBD0 U774 ( .CLK(n891), .C(n892) );
  CKBD0 U775 ( .CLK(n892), .C(n893) );
  CKBD0 U776 ( .CLK(n893), .C(n894) );
  CKBD0 U777 ( .CLK(n894), .C(n895) );
  BUFFD0 U778 ( .I(n895), .Z(n896) );
  CKBD0 U779 ( .CLK(n896), .C(n897) );
  CKBD0 U780 ( .CLK(n897), .C(n898) );
  CKBD0 U781 ( .CLK(n898), .C(n899) );
  CKBD0 U782 ( .CLK(n899), .C(n900) );
  CKBD0 U783 ( .CLK(n900), .C(n901) );
  CKBD0 U784 ( .CLK(n901), .C(n902) );
  CKBD0 U785 ( .CLK(n902), .C(n903) );
  CKBD0 U786 ( .CLK(n903), .C(n904) );
  CKBD0 U787 ( .CLK(n904), .C(n905) );
  BUFFD0 U788 ( .I(n905), .Z(n906) );
  CKBD0 U789 ( .CLK(n906), .C(n907) );
  CKBD0 U790 ( .CLK(n907), .C(n908) );
  CKBD0 U791 ( .CLK(n908), .C(n909) );
  CKBD0 U792 ( .CLK(n909), .C(n910) );
  CKBD0 U793 ( .CLK(n910), .C(n911) );
  CKBD0 U794 ( .CLK(n911), .C(n912) );
  CKBD0 U795 ( .CLK(n912), .C(n913) );
  CKBD0 U796 ( .CLK(n913), .C(n914) );
  CKBD0 U797 ( .CLK(n914), .C(n915) );
  CKBD0 U798 ( .CLK(n915), .C(n916) );
  BUFFD0 U799 ( .I(n916), .Z(n917) );
  CKBD0 U800 ( .CLK(n917), .C(n918) );
  CKBD0 U801 ( .CLK(n918), .C(n919) );
  CKBD0 U802 ( .CLK(n919), .C(n920) );
  CKBD0 U803 ( .CLK(n920), .C(n921) );
  CKBD0 U804 ( .CLK(n921), .C(n922) );
  CKBD0 U805 ( .CLK(n922), .C(n923) );
  CKBD0 U806 ( .CLK(n923), .C(n924) );
  CKBD0 U807 ( .CLK(n924), .C(n925) );
  CKBD0 U808 ( .CLK(n925), .C(n926) );
  CKBD0 U809 ( .CLK(n926), .C(n927) );
  BUFFD0 U810 ( .I(n927), .Z(n928) );
  CKBD0 U811 ( .CLK(n928), .C(n929) );
  CKBD0 U812 ( .CLK(n929), .C(n930) );
  CKBD0 U813 ( .CLK(n930), .C(n931) );
  CKBD0 U814 ( .CLK(n931), .C(n932) );
  BUFFD0 U815 ( .I(n8877), .Z(n933) );
  CKBD0 U816 ( .CLK(FrameSR[7]), .C(n934) );
  CKBD0 U817 ( .CLK(n934), .C(n935) );
  CKBD0 U818 ( .CLK(n935), .C(n936) );
  BUFFD0 U819 ( .I(n6965), .Z(n937) );
  CKBD0 U820 ( .CLK(FrameSR[8]), .C(n938) );
  BUFFD0 U821 ( .I(n6828), .Z(n939) );
  CKBD0 U822 ( .CLK(FrameSR[9]), .C(n940) );
  BUFFD0 U823 ( .I(n6691), .Z(n941) );
  CKBD0 U824 ( .CLK(FrameSR[10]), .C(n942) );
  BUFFD0 U825 ( .I(n6554), .Z(n943) );
  CKBD0 U826 ( .CLK(FrameSR[11]), .C(n944) );
  BUFFD0 U827 ( .I(n6417), .Z(n945) );
  CKBD0 U828 ( .CLK(FrameSR[12]), .C(n946) );
  BUFFD0 U829 ( .I(n6280), .Z(n947) );
  CKBD0 U830 ( .CLK(FrameSR[13]), .C(n948) );
  BUFFD0 U831 ( .I(n6143), .Z(n949) );
  CKBD0 U832 ( .CLK(FrameSR[14]), .C(n950) );
  BUFFD0 U833 ( .I(n8415), .Z(n951) );
  CKBD0 U834 ( .CLK(FrameSR[18]), .C(n952) );
  CKBD0 U835 ( .CLK(n952), .C(n953) );
  CKBD0 U836 ( .CLK(n953), .C(n954) );
  CKBD0 U837 ( .CLK(n954), .C(n955) );
  CKBD0 U838 ( .CLK(n955), .C(n956) );
  CKBD0 U839 ( .CLK(n956), .C(n957) );
  CKBD0 U840 ( .CLK(n957), .C(n958) );
  CKBD0 U841 ( .CLK(n958), .C(n959) );
  CKBD0 U842 ( .CLK(n959), .C(n960) );
  CKBD0 U843 ( .CLK(n960), .C(n961) );
  BUFFD0 U844 ( .I(n961), .Z(n962) );
  CKBD0 U845 ( .CLK(n962), .C(n963) );
  CKBD0 U846 ( .CLK(n963), .C(n964) );
  CKBD0 U847 ( .CLK(n964), .C(n965) );
  CKBD0 U848 ( .CLK(n965), .C(n966) );
  CKBD0 U849 ( .CLK(n966), .C(n967) );
  CKBD0 U850 ( .CLK(n967), .C(n968) );
  CKBD0 U851 ( .CLK(n968), .C(n969) );
  CKBD0 U852 ( .CLK(n969), .C(n970) );
  CKBD0 U853 ( .CLK(n970), .C(n971) );
  CKBD0 U854 ( .CLK(n971), .C(n972) );
  BUFFD0 U855 ( .I(n972), .Z(n973) );
  CKBD0 U856 ( .CLK(n973), .C(n974) );
  CKBD0 U857 ( .CLK(n974), .C(n975) );
  CKBD0 U858 ( .CLK(n975), .C(n976) );
  CKBD0 U859 ( .CLK(n976), .C(n977) );
  CKBD0 U860 ( .CLK(n977), .C(n978) );
  CKBD0 U861 ( .CLK(n978), .C(n979) );
  CKBD0 U862 ( .CLK(n979), .C(n980) );
  CKBD0 U863 ( .CLK(n980), .C(n981) );
  CKBD0 U864 ( .CLK(n981), .C(n982) );
  CKBD0 U865 ( .CLK(n982), .C(n983) );
  BUFFD0 U866 ( .I(n983), .Z(n984) );
  CKBD0 U867 ( .CLK(n984), .C(n985) );
  CKBD0 U868 ( .CLK(n985), .C(n986) );
  CKBD0 U869 ( .CLK(n986), .C(n987) );
  CKBD0 U870 ( .CLK(n987), .C(n988) );
  CKBD0 U871 ( .CLK(n988), .C(n989) );
  CKBD0 U872 ( .CLK(n989), .C(n990) );
  CKBD0 U873 ( .CLK(n990), .C(n991) );
  CKBD0 U874 ( .CLK(n991), .C(n992) );
  CKBD0 U875 ( .CLK(n992), .C(n993) );
  CKBD0 U876 ( .CLK(n993), .C(n994) );
  BUFFD0 U877 ( .I(n994), .Z(n995) );
  CKBD0 U878 ( .CLK(n995), .C(n996) );
  CKBD0 U879 ( .CLK(n996), .C(n997) );
  CKBD0 U880 ( .CLK(n997), .C(n998) );
  CKBD0 U881 ( .CLK(n998), .C(n999) );
  CKBD0 U882 ( .CLK(n999), .C(n1000) );
  CKBD0 U883 ( .CLK(n1000), .C(n1001) );
  CKBD0 U884 ( .CLK(n1001), .C(n1002) );
  CKBD0 U885 ( .CLK(n1002), .C(n1003) );
  CKBD0 U886 ( .CLK(n1003), .C(n1004) );
  CKBD0 U887 ( .CLK(n1004), .C(n1005) );
  BUFFD0 U888 ( .I(n1005), .Z(n1006) );
  CKBD0 U889 ( .CLK(n1006), .C(n1007) );
  CKBD0 U890 ( .CLK(n1007), .C(n1008) );
  CKBD0 U891 ( .CLK(n1008), .C(n1009) );
  CKBD0 U892 ( .CLK(n1009), .C(n1010) );
  CKBD0 U893 ( .CLK(n1010), .C(n1011) );
  CKBD0 U894 ( .CLK(n1011), .C(n1012) );
  CKBD0 U895 ( .CLK(n1012), .C(n1013) );
  CKBD0 U896 ( .CLK(n1013), .C(n1014) );
  CKBD0 U897 ( .CLK(n1014), .C(n1015) );
  BUFFD0 U898 ( .I(n1015), .Z(n1016) );
  CKBD0 U899 ( .CLK(n1016), .C(n1017) );
  CKBD0 U900 ( .CLK(n1017), .C(n1018) );
  CKBD0 U901 ( .CLK(n1018), .C(n1019) );
  CKBD0 U902 ( .CLK(n1019), .C(n1020) );
  CKBD0 U903 ( .CLK(n1020), .C(n1021) );
  CKBD0 U904 ( .CLK(n1021), .C(n1022) );
  CKBD0 U905 ( .CLK(n1022), .C(n1023) );
  CKBD0 U906 ( .CLK(n1023), .C(n1024) );
  CKBD0 U907 ( .CLK(n1024), .C(n1025) );
  CKBD0 U908 ( .CLK(n1025), .C(n1026) );
  BUFFD0 U909 ( .I(n1026), .Z(n1027) );
  CKBD0 U910 ( .CLK(n1027), .C(n1028) );
  CKBD0 U911 ( .CLK(n1028), .C(n1029) );
  CKBD0 U912 ( .CLK(n1029), .C(n1030) );
  CKBD0 U913 ( .CLK(n1030), .C(n1031) );
  CKBD0 U914 ( .CLK(n1031), .C(n1032) );
  CKBD0 U915 ( .CLK(n1032), .C(n1033) );
  CKBD0 U916 ( .CLK(n1033), .C(n1034) );
  CKBD0 U917 ( .CLK(n1034), .C(n1035) );
  CKBD0 U918 ( .CLK(n1035), .C(n1036) );
  CKBD0 U919 ( .CLK(n1036), .C(n1037) );
  BUFFD0 U920 ( .I(n1037), .Z(n1038) );
  CKBD0 U921 ( .CLK(n1038), .C(n1039) );
  CKBD0 U922 ( .CLK(n1039), .C(n1040) );
  CKBD0 U923 ( .CLK(n1040), .C(n1041) );
  CKBD0 U924 ( .CLK(n1041), .C(n1042) );
  CKBD0 U925 ( .CLK(n1042), .C(n1043) );
  CKBD0 U926 ( .CLK(n1043), .C(n1044) );
  CKBD0 U927 ( .CLK(n1044), .C(n1045) );
  CKBD0 U928 ( .CLK(n1045), .C(n1046) );
  CKBD0 U929 ( .CLK(n1046), .C(n1047) );
  CKBD0 U930 ( .CLK(n1047), .C(n1048) );
  CKBD0 U931 ( .CLK(n1048), .C(n1049) );
  BUFFD0 U932 ( .I(n8162), .Z(n1050) );
  CKBD0 U933 ( .CLK(FrameSR[23]), .C(n1051) );
  CKBD0 U934 ( .CLK(n1051), .C(n1052) );
  CKBD0 U935 ( .CLK(n1052), .C(n1053) );
  CKBD0 U936 ( .CLK(n1053), .C(n1054) );
  CKBD0 U937 ( .CLK(n1054), .C(n1055) );
  BUFFD0 U938 ( .I(n1055), .Z(n1056) );
  CKBD0 U939 ( .CLK(n1056), .C(n1057) );
  CKBD0 U940 ( .CLK(n1057), .C(n1058) );
  CKBD0 U941 ( .CLK(n1058), .C(n1059) );
  CKBD0 U942 ( .CLK(n1059), .C(n1060) );
  CKBD0 U943 ( .CLK(n1060), .C(n1061) );
  CKBD0 U944 ( .CLK(n1061), .C(n1062) );
  CKBD0 U945 ( .CLK(n1062), .C(n1063) );
  CKBD0 U946 ( .CLK(n1063), .C(n1064) );
  CKBD0 U947 ( .CLK(n1064), .C(n1065) );
  CKBD0 U948 ( .CLK(n1065), .C(n1066) );
  BUFFD0 U949 ( .I(n1066), .Z(n1067) );
  CKBD0 U950 ( .CLK(n1067), .C(n1068) );
  CKBD0 U951 ( .CLK(n1068), .C(n1069) );
  CKBD0 U952 ( .CLK(n1069), .C(n1070) );
  CKBD0 U953 ( .CLK(n1070), .C(n1071) );
  CKBD0 U954 ( .CLK(n1071), .C(n1072) );
  CKBD0 U955 ( .CLK(n1072), .C(n1073) );
  CKBD0 U956 ( .CLK(n1073), .C(n1074) );
  CKBD0 U957 ( .CLK(n1074), .C(n1075) );
  CKBD0 U958 ( .CLK(n1075), .C(n1076) );
  CKBD0 U959 ( .CLK(n1076), .C(n1077) );
  BUFFD0 U960 ( .I(n1077), .Z(n1078) );
  CKBD0 U961 ( .CLK(n1078), .C(n1079) );
  CKBD0 U962 ( .CLK(n1079), .C(n1080) );
  CKBD0 U963 ( .CLK(n1080), .C(n1081) );
  CKBD0 U964 ( .CLK(n1081), .C(n1082) );
  CKBD0 U965 ( .CLK(n1082), .C(n1083) );
  CKBD0 U966 ( .CLK(n1083), .C(n1084) );
  CKBD0 U967 ( .CLK(n1084), .C(n1085) );
  CKBD0 U968 ( .CLK(n1085), .C(n1086) );
  CKBD0 U969 ( .CLK(n1086), .C(n1087) );
  CKBD0 U970 ( .CLK(n1087), .C(n1088) );
  BUFFD0 U971 ( .I(n1088), .Z(n1089) );
  CKBD0 U972 ( .CLK(n1089), .C(n1090) );
  CKBD0 U973 ( .CLK(n1090), .C(n1091) );
  CKBD0 U974 ( .CLK(n1091), .C(n1092) );
  CKBD0 U975 ( .CLK(n1092), .C(n1093) );
  CKBD0 U976 ( .CLK(n1093), .C(n1094) );
  CKBD0 U977 ( .CLK(n1094), .C(n1095) );
  CKBD0 U978 ( .CLK(n1095), .C(n1096) );
  CKBD0 U979 ( .CLK(n1096), .C(n1097) );
  CKBD0 U980 ( .CLK(n1097), .C(n1098) );
  CKBD0 U981 ( .CLK(n1098), .C(n1099) );
  BUFFD0 U982 ( .I(n1099), .Z(n1100) );
  CKBD0 U983 ( .CLK(n1100), .C(n1101) );
  CKBD0 U984 ( .CLK(n1101), .C(n1102) );
  CKBD0 U985 ( .CLK(n1102), .C(n1103) );
  CKBD0 U986 ( .CLK(n1103), .C(n1104) );
  CKBD0 U987 ( .CLK(n1104), .C(n1105) );
  CKBD0 U988 ( .CLK(n1105), .C(n1106) );
  CKBD0 U989 ( .CLK(n1106), .C(n1107) );
  CKBD0 U990 ( .CLK(n1107), .C(n1108) );
  CKBD0 U991 ( .CLK(n1108), .C(n1109) );
  BUFFD0 U992 ( .I(n1109), .Z(n1110) );
  CKBD0 U993 ( .CLK(n1110), .C(n1111) );
  CKBD0 U994 ( .CLK(n1111), .C(n1112) );
  CKBD0 U995 ( .CLK(n1112), .C(n1113) );
  CKBD0 U996 ( .CLK(n1113), .C(n1114) );
  CKBD0 U997 ( .CLK(n1114), .C(n1115) );
  CKBD0 U998 ( .CLK(n1115), .C(n1116) );
  CKBD0 U999 ( .CLK(n1116), .C(n1117) );
  CKBD0 U1000 ( .CLK(n1117), .C(n1118) );
  CKBD0 U1001 ( .CLK(n1118), .C(n1119) );
  CKBD0 U1002 ( .CLK(n1119), .C(n1120) );
  BUFFD0 U1003 ( .I(n1120), .Z(n1121) );
  CKBD0 U1004 ( .CLK(n1121), .C(n1122) );
  CKBD0 U1005 ( .CLK(n1122), .C(n1123) );
  CKBD0 U1006 ( .CLK(n1123), .C(n1124) );
  CKBD0 U1007 ( .CLK(n1124), .C(n1125) );
  CKBD0 U1008 ( .CLK(n1125), .C(n1126) );
  CKBD0 U1009 ( .CLK(n1126), .C(n1127) );
  CKBD0 U1010 ( .CLK(n1127), .C(n1128) );
  CKBD0 U1011 ( .CLK(n1128), .C(n1129) );
  CKBD0 U1012 ( .CLK(n1129), .C(n1130) );
  CKBD0 U1013 ( .CLK(n1130), .C(n1131) );
  BUFFD0 U1014 ( .I(n1131), .Z(n1132) );
  CKBD0 U1015 ( .CLK(n1132), .C(n1133) );
  CKBD0 U1016 ( .CLK(n1133), .C(n1134) );
  CKBD0 U1017 ( .CLK(n1134), .C(n1135) );
  CKBD0 U1018 ( .CLK(n1135), .C(n1136) );
  CKBD0 U1019 ( .CLK(n1136), .C(n1137) );
  CKBD0 U1020 ( .CLK(n1137), .C(n1138) );
  CKBD0 U1021 ( .CLK(n1138), .C(n1139) );
  CKBD0 U1022 ( .CLK(n1139), .C(n1140) );
  CKBD0 U1023 ( .CLK(n1140), .C(n1141) );
  CKBD0 U1024 ( .CLK(n1141), .C(n1142) );
  BUFFD0 U1025 ( .I(n1142), .Z(n1143) );
  CKBD0 U1026 ( .CLK(n1143), .C(n1144) );
  CKBD0 U1027 ( .CLK(n1144), .C(n1145) );
  CKBD0 U1028 ( .CLK(n1145), .C(n1146) );
  CKBD0 U1029 ( .CLK(n1146), .C(n1147) );
  CKBD0 U1030 ( .CLK(n1147), .C(n1148) );
  CKBD0 U1031 ( .CLK(n1148), .C(n1149) );
  BUFFD0 U1032 ( .I(n5870), .Z(n1150) );
  CKBD0 U1033 ( .CLK(FrameSR[24]), .C(n1151) );
  BUFFD0 U1034 ( .I(n5734), .Z(n1152) );
  CKBD0 U1035 ( .CLK(FrameSR[25]), .C(n1153) );
  BUFFD0 U1036 ( .I(n5598), .Z(n1154) );
  CKBD0 U1037 ( .CLK(FrameSR[26]), .C(n1155) );
  BUFFD0 U1038 ( .I(n5462), .Z(n1156) );
  CKBD0 U1039 ( .CLK(FrameSR[27]), .C(n1157) );
  BUFFD0 U1040 ( .I(n5326), .Z(n1158) );
  CKBD0 U1041 ( .CLK(FrameSR[28]), .C(n1159) );
  BUFFD0 U1042 ( .I(n5189), .Z(n1160) );
  CKBD0 U1043 ( .CLK(FrameSR[29]), .C(n1161) );
  BUFFD0 U1044 ( .I(n5053), .Z(n1162) );
  CKBD0 U1045 ( .CLK(FrameSR[30]), .C(n1163) );
  BUFFD0 U1046 ( .I(n8550), .Z(n1164) );
  CKBD0 U1047 ( .CLK(FrameSR[39]), .C(n1165) );
  CKBD0 U1048 ( .CLK(n1165), .C(n1166) );
  CKBD0 U1049 ( .CLK(n1166), .C(n1167) );
  BUFFD0 U1050 ( .I(n1167), .Z(n1168) );
  CKBD0 U1051 ( .CLK(n1168), .C(n1169) );
  CKBD0 U1052 ( .CLK(n1169), .C(n1170) );
  CKBD0 U1053 ( .CLK(n1170), .C(n1171) );
  CKBD0 U1054 ( .CLK(n1171), .C(n1172) );
  CKBD0 U1055 ( .CLK(n1172), .C(n1173) );
  CKBD0 U1056 ( .CLK(n1173), .C(n1174) );
  CKBD0 U1057 ( .CLK(n1174), .C(n1175) );
  CKBD0 U1058 ( .CLK(n1175), .C(n1176) );
  CKBD0 U1059 ( .CLK(n1176), .C(n1177) );
  CKBD0 U1060 ( .CLK(n1177), .C(n1178) );
  BUFFD0 U1061 ( .I(n1178), .Z(n1179) );
  CKBD0 U1062 ( .CLK(n1179), .C(n1180) );
  CKBD0 U1063 ( .CLK(n1180), .C(n1181) );
  CKBD0 U1064 ( .CLK(n1181), .C(n1182) );
  CKBD0 U1065 ( .CLK(n1182), .C(n1183) );
  CKBD0 U1066 ( .CLK(n1183), .C(n1184) );
  CKBD0 U1067 ( .CLK(n1184), .C(n1185) );
  CKBD0 U1068 ( .CLK(n1185), .C(n1186) );
  CKBD0 U1069 ( .CLK(n1186), .C(n1187) );
  CKBD0 U1070 ( .CLK(n1187), .C(n1188) );
  BUFFD0 U1071 ( .I(n1188), .Z(n1189) );
  CKBD0 U1072 ( .CLK(n1189), .C(n1190) );
  CKBD0 U1073 ( .CLK(n1190), .C(n1191) );
  CKBD0 U1074 ( .CLK(n1191), .C(n1192) );
  CKBD0 U1075 ( .CLK(n1192), .C(n1193) );
  CKBD0 U1076 ( .CLK(n1193), .C(n1194) );
  CKBD0 U1077 ( .CLK(n1194), .C(n1195) );
  CKBD0 U1078 ( .CLK(n1195), .C(n1196) );
  CKBD0 U1079 ( .CLK(n1196), .C(n1197) );
  CKBD0 U1080 ( .CLK(n1197), .C(n1198) );
  CKBD0 U1081 ( .CLK(n1198), .C(n1199) );
  BUFFD0 U1082 ( .I(n1199), .Z(n1200) );
  CKBD0 U1083 ( .CLK(n1200), .C(n1201) );
  CKBD0 U1084 ( .CLK(n1201), .C(n1202) );
  CKBD0 U1085 ( .CLK(n1202), .C(n1203) );
  CKBD0 U1086 ( .CLK(n1203), .C(n1204) );
  CKBD0 U1087 ( .CLK(n1204), .C(n1205) );
  CKBD0 U1088 ( .CLK(n1205), .C(n1206) );
  CKBD0 U1089 ( .CLK(n1206), .C(n1207) );
  CKBD0 U1090 ( .CLK(n1207), .C(n1208) );
  CKBD0 U1091 ( .CLK(n1208), .C(n1209) );
  CKBD0 U1092 ( .CLK(n1209), .C(n1210) );
  BUFFD0 U1093 ( .I(n1210), .Z(n1211) );
  CKBD0 U1094 ( .CLK(n1211), .C(n1212) );
  CKBD0 U1095 ( .CLK(n1212), .C(n1213) );
  CKBD0 U1096 ( .CLK(n1213), .C(n1214) );
  CKBD0 U1097 ( .CLK(n1214), .C(n1215) );
  CKBD0 U1098 ( .CLK(n1215), .C(n1216) );
  CKBD0 U1099 ( .CLK(n1216), .C(n1217) );
  CKBD0 U1100 ( .CLK(n1217), .C(n1218) );
  CKBD0 U1101 ( .CLK(n1218), .C(n1219) );
  CKBD0 U1102 ( .CLK(n1219), .C(n1220) );
  CKBD0 U1103 ( .CLK(n1220), .C(n1221) );
  BUFFD0 U1104 ( .I(n1221), .Z(n1222) );
  CKBD0 U1105 ( .CLK(n1222), .C(n1223) );
  CKBD0 U1106 ( .CLK(n1223), .C(n1224) );
  CKBD0 U1107 ( .CLK(n1224), .C(n1225) );
  CKBD0 U1108 ( .CLK(n1225), .C(n1226) );
  CKBD0 U1109 ( .CLK(n1226), .C(n1227) );
  CKBD0 U1110 ( .CLK(n1227), .C(n1228) );
  CKBD0 U1111 ( .CLK(n1228), .C(n1229) );
  CKBD0 U1112 ( .CLK(n1229), .C(n1230) );
  CKBD0 U1113 ( .CLK(n1230), .C(n1231) );
  CKBD0 U1114 ( .CLK(n1231), .C(n1232) );
  BUFFD0 U1115 ( .I(n1232), .Z(n1233) );
  CKBD0 U1116 ( .CLK(n1233), .C(n1234) );
  CKBD0 U1117 ( .CLK(n1234), .C(n1235) );
  CKBD0 U1118 ( .CLK(n1235), .C(n1236) );
  CKBD0 U1119 ( .CLK(n1236), .C(n1237) );
  CKBD0 U1120 ( .CLK(n1237), .C(n1238) );
  CKBD0 U1121 ( .CLK(n1238), .C(n1239) );
  CKBD0 U1122 ( .CLK(n1239), .C(n1240) );
  CKBD0 U1123 ( .CLK(n1240), .C(n1241) );
  CKBD0 U1124 ( .CLK(n1241), .C(n1242) );
  CKBD0 U1125 ( .CLK(n1242), .C(n1243) );
  BUFFD0 U1126 ( .I(n1243), .Z(n1244) );
  CKBD0 U1127 ( .CLK(n1244), .C(n1245) );
  CKBD0 U1128 ( .CLK(n1245), .C(n1246) );
  CKBD0 U1129 ( .CLK(n1246), .C(n1247) );
  CKBD0 U1130 ( .CLK(n1247), .C(n1248) );
  CKBD0 U1131 ( .CLK(n1248), .C(n1249) );
  CKBD0 U1132 ( .CLK(n1249), .C(n1250) );
  CKBD0 U1133 ( .CLK(n1250), .C(n1251) );
  CKBD0 U1134 ( .CLK(n1251), .C(n1252) );
  CKBD0 U1135 ( .CLK(n1252), .C(n1253) );
  CKBD0 U1136 ( .CLK(n1253), .C(n1254) );
  BUFFD0 U1137 ( .I(n1254), .Z(n1255) );
  CKBD0 U1138 ( .CLK(n1255), .C(n1256) );
  CKBD0 U1139 ( .CLK(n1256), .C(n1257) );
  CKBD0 U1140 ( .CLK(n1257), .C(n1258) );
  CKBD0 U1141 ( .CLK(n1258), .C(n1259) );
  CKBD0 U1142 ( .CLK(n1259), .C(n1260) );
  CKBD0 U1143 ( .CLK(n1260), .C(n1261) );
  CKBD0 U1144 ( .CLK(n1261), .C(n1262) );
  CKBD0 U1145 ( .CLK(n1262), .C(n1263) );
  BUFFD0 U1146 ( .I(n4781), .Z(n1264) );
  CKBD0 U1147 ( .CLK(FrameSR[40]), .C(n1265) );
  BUFFD0 U1148 ( .I(n4645), .Z(n1266) );
  CKBD0 U1149 ( .CLK(FrameSR[41]), .C(n1267) );
  BUFFD0 U1150 ( .I(n4509), .Z(n1268) );
  CKBD0 U1151 ( .CLK(FrameSR[42]), .C(n1269) );
  BUFFD0 U1152 ( .I(n4373), .Z(n1270) );
  CKBD0 U1153 ( .CLK(FrameSR[43]), .C(n1271) );
  BUFFD0 U1154 ( .I(n4236), .Z(n1272) );
  CKBD0 U1155 ( .CLK(FrameSR[44]), .C(n1273) );
  BUFFD0 U1156 ( .I(n4100), .Z(n1274) );
  CKBD0 U1157 ( .CLK(FrameSR[45]), .C(n1275) );
  BUFFD0 U1158 ( .I(n3964), .Z(n1276) );
  CKBD0 U1159 ( .CLK(FrameSR[46]), .C(n1277) );
  BUFFD0 U1160 ( .I(n8152), .Z(n1278) );
  CKBD0 U1161 ( .CLK(FrameSR[55]), .C(n1279) );
  CKBD0 U1162 ( .CLK(n1279), .C(n1280) );
  CKBD0 U1163 ( .CLK(n1280), .C(n1281) );
  CKBD0 U1164 ( .CLK(n1281), .C(n1282) );
  CKBD0 U1165 ( .CLK(n1282), .C(n1283) );
  CKBD0 U1166 ( .CLK(n1283), .C(n1284) );
  CKBD0 U1167 ( .CLK(n1284), .C(n1285) );
  CKBD0 U1168 ( .CLK(n1285), .C(n1286) );
  CKBD0 U1169 ( .CLK(n1286), .C(n1287) );
  BUFFD0 U1170 ( .I(n1287), .Z(n1288) );
  CKBD0 U1171 ( .CLK(n1288), .C(n1289) );
  CKBD0 U1172 ( .CLK(n1289), .C(n1290) );
  CKBD0 U1173 ( .CLK(n1290), .C(n1291) );
  CKBD0 U1174 ( .CLK(n1291), .C(n1292) );
  CKBD0 U1175 ( .CLK(n1292), .C(n1293) );
  CKBD0 U1176 ( .CLK(n1293), .C(n1294) );
  CKBD0 U1177 ( .CLK(n1294), .C(n1295) );
  CKBD0 U1178 ( .CLK(n1295), .C(n1296) );
  CKBD0 U1179 ( .CLK(n1296), .C(n1297) );
  CKBD0 U1180 ( .CLK(n1297), .C(n1298) );
  BUFFD0 U1181 ( .I(n1298), .Z(n1299) );
  CKBD0 U1182 ( .CLK(n1299), .C(n1300) );
  CKBD0 U1183 ( .CLK(n1300), .C(n1301) );
  CKBD0 U1184 ( .CLK(n1301), .C(n1302) );
  CKBD0 U1185 ( .CLK(n1302), .C(n1303) );
  CKBD0 U1186 ( .CLK(n1303), .C(n1304) );
  CKBD0 U1187 ( .CLK(n1304), .C(n1305) );
  CKBD0 U1188 ( .CLK(n1305), .C(n1306) );
  CKBD0 U1189 ( .CLK(n1306), .C(n1307) );
  CKBD0 U1190 ( .CLK(n1307), .C(n1308) );
  CKBD0 U1191 ( .CLK(n1308), .C(n1309) );
  BUFFD0 U1192 ( .I(n1309), .Z(n1310) );
  CKBD0 U1193 ( .CLK(n1310), .C(n1311) );
  CKBD0 U1194 ( .CLK(n1311), .C(n1312) );
  CKBD0 U1195 ( .CLK(n1312), .C(n1313) );
  CKBD0 U1196 ( .CLK(n1313), .C(n1314) );
  CKBD0 U1197 ( .CLK(n1314), .C(n1315) );
  CKBD0 U1198 ( .CLK(n1315), .C(n1316) );
  CKBD0 U1199 ( .CLK(n1316), .C(n1317) );
  CKBD0 U1200 ( .CLK(n1317), .C(n1318) );
  CKBD0 U1201 ( .CLK(n1318), .C(n1319) );
  BUFFD0 U1202 ( .I(n1319), .Z(n1320) );
  CKBD0 U1203 ( .CLK(n1320), .C(n1321) );
  CKBD0 U1204 ( .CLK(n1321), .C(n1322) );
  CKBD0 U1205 ( .CLK(n1322), .C(n1323) );
  CKBD0 U1206 ( .CLK(n1323), .C(n1324) );
  CKBD0 U1207 ( .CLK(n1324), .C(n1325) );
  CKBD0 U1208 ( .CLK(n1325), .C(n1326) );
  CKBD0 U1209 ( .CLK(n1326), .C(n1327) );
  CKBD0 U1210 ( .CLK(n1327), .C(n1328) );
  CKBD0 U1211 ( .CLK(n1328), .C(n1329) );
  CKBD0 U1212 ( .CLK(n1329), .C(n1330) );
  BUFFD0 U1213 ( .I(n1330), .Z(n1331) );
  CKBD0 U1214 ( .CLK(n1331), .C(n1332) );
  CKBD0 U1215 ( .CLK(n1332), .C(n1333) );
  CKBD0 U1216 ( .CLK(n1333), .C(n1334) );
  CKBD0 U1217 ( .CLK(n1334), .C(n1335) );
  CKBD0 U1218 ( .CLK(n1335), .C(n1336) );
  CKBD0 U1219 ( .CLK(n1336), .C(n1337) );
  CKBD0 U1220 ( .CLK(n1337), .C(n1338) );
  CKBD0 U1221 ( .CLK(n1338), .C(n1339) );
  CKBD0 U1222 ( .CLK(n1339), .C(n1340) );
  CKBD0 U1223 ( .CLK(n1340), .C(n1341) );
  BUFFD0 U1224 ( .I(n1341), .Z(n1342) );
  CKBD0 U1225 ( .CLK(n1342), .C(n1343) );
  CKBD0 U1226 ( .CLK(n1343), .C(n1344) );
  CKBD0 U1227 ( .CLK(n1344), .C(n1345) );
  CKBD0 U1228 ( .CLK(n1345), .C(n1346) );
  CKBD0 U1229 ( .CLK(n1346), .C(n1347) );
  CKBD0 U1230 ( .CLK(n1347), .C(n1348) );
  CKBD0 U1231 ( .CLK(n1348), .C(n1349) );
  CKBD0 U1232 ( .CLK(n1349), .C(n1350) );
  CKBD0 U1233 ( .CLK(n1350), .C(n1351) );
  CKBD0 U1234 ( .CLK(n1351), .C(n1352) );
  BUFFD0 U1235 ( .I(n1352), .Z(n1353) );
  CKBD0 U1236 ( .CLK(n1353), .C(n1354) );
  CKBD0 U1237 ( .CLK(n1354), .C(n1355) );
  CKBD0 U1238 ( .CLK(n1355), .C(n1356) );
  CKBD0 U1239 ( .CLK(n1356), .C(n1357) );
  CKBD0 U1240 ( .CLK(n1357), .C(n1358) );
  CKBD0 U1241 ( .CLK(n1358), .C(n1359) );
  CKBD0 U1242 ( .CLK(n1359), .C(n1360) );
  CKBD0 U1243 ( .CLK(n1360), .C(n1361) );
  CKBD0 U1244 ( .CLK(n1361), .C(n1362) );
  CKBD0 U1245 ( .CLK(n1362), .C(n1363) );
  BUFFD0 U1246 ( .I(n1363), .Z(n1364) );
  CKBD0 U1247 ( .CLK(n1364), .C(n1365) );
  CKBD0 U1248 ( .CLK(n1365), .C(n1366) );
  CKBD0 U1249 ( .CLK(n1366), .C(n1367) );
  CKBD0 U1250 ( .CLK(n1367), .C(n1368) );
  CKBD0 U1251 ( .CLK(n1368), .C(n1369) );
  CKBD0 U1252 ( .CLK(n1369), .C(n1370) );
  CKBD0 U1253 ( .CLK(n1370), .C(n1371) );
  CKBD0 U1254 ( .CLK(n1371), .C(n1372) );
  CKBD0 U1255 ( .CLK(n1372), .C(n1373) );
  CKBD0 U1256 ( .CLK(n1373), .C(n1374) );
  BUFFD0 U1257 ( .I(n1374), .Z(n1375) );
  CKBD0 U1258 ( .CLK(n1375), .C(n1376) );
  CKBD0 U1259 ( .CLK(n1376), .C(n1377) );
  BUFFD0 U1260 ( .I(n3692), .Z(n1378) );
  CKBD0 U1261 ( .CLK(FrameSR[56]), .C(n1379) );
  BUFFD0 U1262 ( .I(n3556), .Z(n1380) );
  CKBD0 U1263 ( .CLK(FrameSR[57]), .C(n1381) );
  BUFFD0 U1264 ( .I(n3420), .Z(n1382) );
  CKBD0 U1265 ( .CLK(FrameSR[58]), .C(n1383) );
  BUFFD0 U1266 ( .I(n3284), .Z(n1384) );
  CKBD0 U1267 ( .CLK(FrameSR[59]), .C(n1385) );
  BUFFD0 U1268 ( .I(n3148), .Z(n1386) );
  CKBD0 U1269 ( .CLK(FrameSR[60]), .C(n1387) );
  BUFFD0 U1270 ( .I(n3012), .Z(n1388) );
  CKBD0 U1271 ( .CLK(FrameSR[61]), .C(n1389) );
  BUFFD0 U1272 ( .I(n8888), .Z(n1390) );
  CKBD0 U1273 ( .CLK(FrameSR[3]), .C(n1391) );
  CKBD0 U1274 ( .CLK(n1391), .C(n1392) );
  BUFFD0 U1275 ( .I(n8172), .Z(n1393) );
  CKBD0 U1276 ( .CLK(FrameSR[19]), .C(n1394) );
  CKBD0 U1277 ( .CLK(n1394), .C(n1395) );
  CKBD0 U1278 ( .CLK(n1395), .C(n1396) );
  CKBD0 U1279 ( .CLK(n1396), .C(n1397) );
  CKBD0 U1280 ( .CLK(n1397), .C(n1398) );
  CKBD0 U1281 ( .CLK(n1398), .C(n1399) );
  CKBD0 U1282 ( .CLK(n1399), .C(n1400) );
  CKBD0 U1283 ( .CLK(n1400), .C(n1401) );
  CKBD0 U1284 ( .CLK(n1401), .C(n1402) );
  BUFFD0 U1285 ( .I(n1402), .Z(n1403) );
  CKBD0 U1286 ( .CLK(n1403), .C(n1404) );
  CKBD0 U1287 ( .CLK(n1404), .C(n1405) );
  CKBD0 U1288 ( .CLK(n1405), .C(n1406) );
  CKBD0 U1289 ( .CLK(n1406), .C(n1407) );
  CKBD0 U1290 ( .CLK(n1407), .C(n1408) );
  CKBD0 U1291 ( .CLK(n1408), .C(n1409) );
  CKBD0 U1292 ( .CLK(n1409), .C(n1410) );
  CKBD0 U1293 ( .CLK(n1410), .C(n1411) );
  CKBD0 U1294 ( .CLK(n1411), .C(n1412) );
  CKBD0 U1295 ( .CLK(n1412), .C(n1413) );
  BUFFD0 U1296 ( .I(n1413), .Z(n1414) );
  CKBD0 U1297 ( .CLK(n1414), .C(n1415) );
  CKBD0 U1298 ( .CLK(n1415), .C(n1416) );
  CKBD0 U1299 ( .CLK(n1416), .C(n1417) );
  CKBD0 U1300 ( .CLK(n1417), .C(n1418) );
  CKBD0 U1301 ( .CLK(n1418), .C(n1419) );
  CKBD0 U1302 ( .CLK(n1419), .C(n1420) );
  CKBD0 U1303 ( .CLK(n1420), .C(n1421) );
  CKBD0 U1304 ( .CLK(n1421), .C(n1422) );
  CKBD0 U1305 ( .CLK(n1422), .C(n1423) );
  BUFFD0 U1306 ( .I(n1423), .Z(n1424) );
  CKBD0 U1307 ( .CLK(n1424), .C(n1425) );
  CKBD0 U1308 ( .CLK(n1425), .C(n1426) );
  CKBD0 U1309 ( .CLK(n1426), .C(n1427) );
  CKBD0 U1310 ( .CLK(n1427), .C(n1428) );
  CKBD0 U1311 ( .CLK(n1428), .C(n1429) );
  CKBD0 U1312 ( .CLK(n1429), .C(n1430) );
  CKBD0 U1313 ( .CLK(n1430), .C(n1431) );
  CKBD0 U1314 ( .CLK(n1431), .C(n1432) );
  CKBD0 U1315 ( .CLK(n1432), .C(n1433) );
  CKBD0 U1316 ( .CLK(n1433), .C(n1434) );
  BUFFD0 U1317 ( .I(n1434), .Z(n1435) );
  CKBD0 U1318 ( .CLK(n1435), .C(n1436) );
  CKBD0 U1319 ( .CLK(n1436), .C(n1437) );
  CKBD0 U1320 ( .CLK(n1437), .C(n1438) );
  CKBD0 U1321 ( .CLK(n1438), .C(n1439) );
  CKBD0 U1322 ( .CLK(n1439), .C(n1440) );
  CKBD0 U1323 ( .CLK(n1440), .C(n1441) );
  CKBD0 U1324 ( .CLK(n1441), .C(n1442) );
  CKBD0 U1325 ( .CLK(n1442), .C(n1443) );
  CKBD0 U1326 ( .CLK(n1443), .C(n1444) );
  CKBD0 U1327 ( .CLK(n1444), .C(n1445) );
  BUFFD0 U1328 ( .I(n1445), .Z(n1446) );
  CKBD0 U1329 ( .CLK(n1446), .C(n1447) );
  CKBD0 U1330 ( .CLK(n1447), .C(n1448) );
  CKBD0 U1331 ( .CLK(n1448), .C(n1449) );
  CKBD0 U1332 ( .CLK(n1449), .C(n1450) );
  CKBD0 U1333 ( .CLK(n1450), .C(n1451) );
  CKBD0 U1334 ( .CLK(n1451), .C(n1452) );
  CKBD0 U1335 ( .CLK(n1452), .C(n1453) );
  CKBD0 U1336 ( .CLK(n1453), .C(n1454) );
  CKBD0 U1337 ( .CLK(n1454), .C(n1455) );
  CKBD0 U1338 ( .CLK(n1455), .C(n1456) );
  BUFFD0 U1339 ( .I(n1456), .Z(n1457) );
  CKBD0 U1340 ( .CLK(n1457), .C(n1458) );
  CKBD0 U1341 ( .CLK(n1458), .C(n1459) );
  CKBD0 U1342 ( .CLK(n1459), .C(n1460) );
  CKBD0 U1343 ( .CLK(n1460), .C(n1461) );
  CKBD0 U1344 ( .CLK(n1461), .C(n1462) );
  CKBD0 U1345 ( .CLK(n1462), .C(n1463) );
  CKBD0 U1346 ( .CLK(n1463), .C(n1464) );
  CKBD0 U1347 ( .CLK(n1464), .C(n1465) );
  CKBD0 U1348 ( .CLK(n1465), .C(n1466) );
  CKBD0 U1349 ( .CLK(n1466), .C(n1467) );
  BUFFD0 U1350 ( .I(n1467), .Z(n1468) );
  CKBD0 U1351 ( .CLK(n1468), .C(n1469) );
  CKBD0 U1352 ( .CLK(n1469), .C(n1470) );
  CKBD0 U1353 ( .CLK(n1470), .C(n1471) );
  CKBD0 U1354 ( .CLK(n1471), .C(n1472) );
  CKBD0 U1355 ( .CLK(n1472), .C(n1473) );
  CKBD0 U1356 ( .CLK(n1473), .C(n1474) );
  CKBD0 U1357 ( .CLK(n1474), .C(n1475) );
  CKBD0 U1358 ( .CLK(n1475), .C(n1476) );
  CKBD0 U1359 ( .CLK(n1476), .C(n1477) );
  CKBD0 U1360 ( .CLK(n1477), .C(n1478) );
  BUFFD0 U1361 ( .I(n1478), .Z(n1479) );
  CKBD0 U1362 ( .CLK(n1479), .C(n1480) );
  CKBD0 U1363 ( .CLK(n1480), .C(n1481) );
  CKBD0 U1364 ( .CLK(n1481), .C(n1482) );
  CKBD0 U1365 ( .CLK(n1482), .C(n1483) );
  CKBD0 U1366 ( .CLK(n1483), .C(n1484) );
  CKBD0 U1367 ( .CLK(n1484), .C(n1485) );
  CKBD0 U1368 ( .CLK(n1485), .C(n1486) );
  CKBD0 U1369 ( .CLK(n1486), .C(n1487) );
  CKBD0 U1370 ( .CLK(n1487), .C(n1488) );
  BUFFD0 U1371 ( .I(n1488), .Z(n1489) );
  CKBD0 U1372 ( .CLK(n1489), .C(n1490) );
  CKBD0 U1373 ( .CLK(n1490), .C(n1491) );
  BUFFD0 U1374 ( .I(n8266), .Z(n1492) );
  CKBD0 U1375 ( .CLK(FrameSR[33]), .C(n1493) );
  CKBD0 U1376 ( .CLK(n1493), .C(n1494) );
  CKBD0 U1377 ( .CLK(n1494), .C(n1495) );
  CKBD0 U1378 ( .CLK(n1495), .C(n1496) );
  CKBD0 U1379 ( .CLK(n1496), .C(n1497) );
  CKBD0 U1380 ( .CLK(n1497), .C(n1498) );
  CKBD0 U1381 ( .CLK(n1498), .C(n1499) );
  CKBD0 U1382 ( .CLK(n1499), .C(n1500) );
  BUFFD0 U1383 ( .I(n1500), .Z(n1501) );
  CKBD0 U1384 ( .CLK(n1501), .C(n1502) );
  CKBD0 U1385 ( .CLK(n1502), .C(n1503) );
  CKBD0 U1386 ( .CLK(n1503), .C(n1504) );
  CKBD0 U1387 ( .CLK(n1504), .C(n1505) );
  CKBD0 U1388 ( .CLK(n1505), .C(n1506) );
  CKBD0 U1389 ( .CLK(n1506), .C(n1507) );
  CKBD0 U1390 ( .CLK(n1507), .C(n1508) );
  CKBD0 U1391 ( .CLK(n1508), .C(n1509) );
  CKBD0 U1392 ( .CLK(n1509), .C(n1510) );
  CKBD0 U1393 ( .CLK(n1510), .C(n1511) );
  BUFFD0 U1394 ( .I(n1511), .Z(n1512) );
  CKBD0 U1395 ( .CLK(n1512), .C(n1513) );
  CKBD0 U1396 ( .CLK(n1513), .C(n1514) );
  CKBD0 U1397 ( .CLK(n1514), .C(n1515) );
  CKBD0 U1398 ( .CLK(n1515), .C(n1516) );
  CKBD0 U1399 ( .CLK(n1516), .C(n1517) );
  CKBD0 U1400 ( .CLK(n1517), .C(n1518) );
  CKBD0 U1401 ( .CLK(n1518), .C(n1519) );
  CKBD0 U1402 ( .CLK(n1519), .C(n1520) );
  CKBD0 U1403 ( .CLK(n1520), .C(n1521) );
  CKBD0 U1404 ( .CLK(n1521), .C(n1522) );
  BUFFD0 U1405 ( .I(n1522), .Z(n1523) );
  CKBD0 U1406 ( .CLK(n1523), .C(n1524) );
  CKBD0 U1407 ( .CLK(n1524), .C(n1525) );
  CKBD0 U1408 ( .CLK(n1525), .C(n1526) );
  CKBD0 U1409 ( .CLK(n1526), .C(n1527) );
  CKBD0 U1410 ( .CLK(n1527), .C(n1528) );
  CKBD0 U1411 ( .CLK(n1528), .C(n1529) );
  CKBD0 U1412 ( .CLK(n1529), .C(n1530) );
  CKBD0 U1413 ( .CLK(n1530), .C(n1531) );
  CKBD0 U1414 ( .CLK(n1531), .C(n1532) );
  CKBD0 U1415 ( .CLK(n1532), .C(n1533) );
  BUFFD0 U1416 ( .I(n1533), .Z(n1534) );
  CKBD0 U1417 ( .CLK(n1534), .C(n1535) );
  CKBD0 U1418 ( .CLK(n1535), .C(n1536) );
  CKBD0 U1419 ( .CLK(n1536), .C(n1537) );
  CKBD0 U1420 ( .CLK(n1537), .C(n1538) );
  CKBD0 U1421 ( .CLK(n1538), .C(n1539) );
  CKBD0 U1422 ( .CLK(n1539), .C(n1540) );
  CKBD0 U1423 ( .CLK(n1540), .C(n1541) );
  CKBD0 U1424 ( .CLK(n1541), .C(n1542) );
  CKBD0 U1425 ( .CLK(n1542), .C(n1543) );
  BUFFD0 U1426 ( .I(n1543), .Z(n1544) );
  CKBD0 U1427 ( .CLK(n1544), .C(n1545) );
  CKBD0 U1428 ( .CLK(n1545), .C(n1546) );
  CKBD0 U1429 ( .CLK(n1546), .C(n1547) );
  CKBD0 U1430 ( .CLK(n1547), .C(n1548) );
  CKBD0 U1431 ( .CLK(n1548), .C(n1549) );
  CKBD0 U1432 ( .CLK(n1549), .C(n1550) );
  CKBD0 U1433 ( .CLK(n1550), .C(n1551) );
  CKBD0 U1434 ( .CLK(n1551), .C(n1552) );
  CKBD0 U1435 ( .CLK(n1552), .C(n1553) );
  CKBD0 U1436 ( .CLK(n1553), .C(n1554) );
  BUFFD0 U1437 ( .I(n1554), .Z(n1555) );
  CKBD0 U1438 ( .CLK(n1555), .C(n1556) );
  CKBD0 U1439 ( .CLK(n1556), .C(n1557) );
  CKBD0 U1440 ( .CLK(n1557), .C(n1558) );
  CKBD0 U1441 ( .CLK(n1558), .C(n1559) );
  CKBD0 U1442 ( .CLK(n1559), .C(n1560) );
  CKBD0 U1443 ( .CLK(n1560), .C(n1561) );
  CKBD0 U1444 ( .CLK(n1561), .C(n1562) );
  CKBD0 U1445 ( .CLK(n1562), .C(n1563) );
  CKBD0 U1446 ( .CLK(n1563), .C(n1564) );
  CKBD0 U1447 ( .CLK(n1564), .C(n1565) );
  BUFFD0 U1448 ( .I(n1565), .Z(n1566) );
  CKBD0 U1449 ( .CLK(n1566), .C(n1567) );
  CKBD0 U1450 ( .CLK(n1567), .C(n1568) );
  CKBD0 U1451 ( .CLK(n1568), .C(n1569) );
  CKBD0 U1452 ( .CLK(n1569), .C(n1570) );
  CKBD0 U1453 ( .CLK(n1570), .C(n1571) );
  CKBD0 U1454 ( .CLK(n1571), .C(n1572) );
  CKBD0 U1455 ( .CLK(n1572), .C(n1573) );
  CKBD0 U1456 ( .CLK(n1573), .C(n1574) );
  CKBD0 U1457 ( .CLK(n1574), .C(n1575) );
  CKBD0 U1458 ( .CLK(n1575), .C(n1576) );
  BUFFD0 U1459 ( .I(n1576), .Z(n1577) );
  CKBD0 U1460 ( .CLK(n1577), .C(n1578) );
  CKBD0 U1461 ( .CLK(n1578), .C(n1579) );
  CKBD0 U1462 ( .CLK(n1579), .C(n1580) );
  CKBD0 U1463 ( .CLK(n1580), .C(n1581) );
  CKBD0 U1464 ( .CLK(n1581), .C(n1582) );
  CKBD0 U1465 ( .CLK(n1582), .C(n1583) );
  CKBD0 U1466 ( .CLK(n1583), .C(n1584) );
  CKBD0 U1467 ( .CLK(n1584), .C(n1585) );
  CKBD0 U1468 ( .CLK(n1585), .C(n1586) );
  CKBD0 U1469 ( .CLK(n1586), .C(n1587) );
  BUFFD0 U1470 ( .I(n1587), .Z(n1588) );
  CKBD0 U1471 ( .CLK(n1588), .C(n1589) );
  CKBD0 U1472 ( .CLK(n1589), .C(n1590) );
  BUFFD0 U1473 ( .I(n8996), .Z(n1591) );
  CKBD0 U1474 ( .CLK(FrameSR[48]), .C(n1592) );
  CKBD0 U1475 ( .CLK(n1592), .C(n1593) );
  BUFFD0 U1476 ( .I(n1593), .Z(n1594) );
  CKBD0 U1477 ( .CLK(n1594), .C(n1595) );
  CKBD0 U1478 ( .CLK(n1595), .C(n1596) );
  CKBD0 U1479 ( .CLK(n1596), .C(n1597) );
  CKBD0 U1480 ( .CLK(n1597), .C(n1598) );
  CKBD0 U1481 ( .CLK(n1598), .C(n1599) );
  CKBD0 U1482 ( .CLK(n1599), .C(n1600) );
  CKBD0 U1483 ( .CLK(n1600), .C(n1601) );
  CKBD0 U1484 ( .CLK(n1601), .C(n1602) );
  CKBD0 U1485 ( .CLK(n1602), .C(n1603) );
  CKBD0 U1486 ( .CLK(n1603), .C(n1604) );
  BUFFD0 U1487 ( .I(n1604), .Z(n1605) );
  CKBD0 U1488 ( .CLK(n1605), .C(n1606) );
  CKBD0 U1489 ( .CLK(n1606), .C(n1607) );
  CKBD0 U1490 ( .CLK(n1607), .C(n1608) );
  CKBD0 U1491 ( .CLK(n1608), .C(n1609) );
  CKBD0 U1492 ( .CLK(n1609), .C(n1610) );
  CKBD0 U1493 ( .CLK(n1610), .C(n1611) );
  CKBD0 U1494 ( .CLK(n1611), .C(n1612) );
  CKBD0 U1495 ( .CLK(n1612), .C(n1613) );
  CKBD0 U1496 ( .CLK(n1613), .C(n1614) );
  BUFFD0 U1497 ( .I(n1614), .Z(n1615) );
  CKBD0 U1498 ( .CLK(n1615), .C(n1616) );
  CKBD0 U1499 ( .CLK(n1616), .C(n1617) );
  CKBD0 U1500 ( .CLK(n1617), .C(n1618) );
  CKBD0 U1501 ( .CLK(n1618), .C(n1619) );
  CKBD0 U1502 ( .CLK(n1619), .C(n1620) );
  CKBD0 U1503 ( .CLK(n1620), .C(n1621) );
  CKBD0 U1504 ( .CLK(n1621), .C(n1622) );
  CKBD0 U1505 ( .CLK(n1622), .C(n1623) );
  CKBD0 U1506 ( .CLK(n1623), .C(n1624) );
  CKBD0 U1507 ( .CLK(n1624), .C(n1625) );
  BUFFD0 U1508 ( .I(n1625), .Z(n1626) );
  CKBD0 U1509 ( .CLK(n1626), .C(n1627) );
  CKBD0 U1510 ( .CLK(n1627), .C(n1628) );
  CKBD0 U1511 ( .CLK(n1628), .C(n1629) );
  CKBD0 U1512 ( .CLK(n1629), .C(n1630) );
  CKBD0 U1513 ( .CLK(n1630), .C(n1631) );
  CKBD0 U1514 ( .CLK(n1631), .C(n1632) );
  CKBD0 U1515 ( .CLK(n1632), .C(n1633) );
  CKBD0 U1516 ( .CLK(n1633), .C(n1634) );
  CKBD0 U1517 ( .CLK(n1634), .C(n1635) );
  CKBD0 U1518 ( .CLK(n1635), .C(n1636) );
  BUFFD0 U1519 ( .I(n1636), .Z(n1637) );
  CKBD0 U1520 ( .CLK(n1637), .C(n1638) );
  CKBD0 U1521 ( .CLK(n1638), .C(n1639) );
  CKBD0 U1522 ( .CLK(n1639), .C(n1640) );
  CKBD0 U1523 ( .CLK(n1640), .C(n1641) );
  CKBD0 U1524 ( .CLK(n1641), .C(n1642) );
  CKBD0 U1525 ( .CLK(n1642), .C(n1643) );
  CKBD0 U1526 ( .CLK(n1643), .C(n1644) );
  CKBD0 U1527 ( .CLK(n1644), .C(n1645) );
  CKBD0 U1528 ( .CLK(n1645), .C(n1646) );
  CKBD0 U1529 ( .CLK(n1646), .C(n1647) );
  BUFFD0 U1530 ( .I(n1647), .Z(n1648) );
  CKBD0 U1531 ( .CLK(n1648), .C(n1649) );
  CKBD0 U1532 ( .CLK(n1649), .C(n1650) );
  CKBD0 U1533 ( .CLK(n1650), .C(n1651) );
  CKBD0 U1534 ( .CLK(n1651), .C(n1652) );
  CKBD0 U1535 ( .CLK(n1652), .C(n1653) );
  CKBD0 U1536 ( .CLK(n1653), .C(n1654) );
  CKBD0 U1537 ( .CLK(n1654), .C(n1655) );
  CKBD0 U1538 ( .CLK(n1655), .C(n1656) );
  CKBD0 U1539 ( .CLK(n1656), .C(n1657) );
  CKBD0 U1540 ( .CLK(n1657), .C(n1658) );
  BUFFD0 U1541 ( .I(n1658), .Z(n1659) );
  CKBD0 U1542 ( .CLK(n1659), .C(n1660) );
  CKBD0 U1543 ( .CLK(n1660), .C(n1661) );
  CKBD0 U1544 ( .CLK(n1661), .C(n1662) );
  CKBD0 U1545 ( .CLK(n1662), .C(n1663) );
  CKBD0 U1546 ( .CLK(n1663), .C(n1664) );
  CKBD0 U1547 ( .CLK(n1664), .C(n1665) );
  CKBD0 U1548 ( .CLK(n1665), .C(n1666) );
  CKBD0 U1549 ( .CLK(n1666), .C(n1667) );
  CKBD0 U1550 ( .CLK(n1667), .C(n1668) );
  CKBD0 U1551 ( .CLK(n1668), .C(n1669) );
  BUFFD0 U1552 ( .I(n1669), .Z(n1670) );
  CKBD0 U1553 ( .CLK(n1670), .C(n1671) );
  CKBD0 U1554 ( .CLK(n1671), .C(n1672) );
  CKBD0 U1555 ( .CLK(n1672), .C(n1673) );
  CKBD0 U1556 ( .CLK(n1673), .C(n1674) );
  CKBD0 U1557 ( .CLK(n1674), .C(n1675) );
  CKBD0 U1558 ( .CLK(n1675), .C(n1676) );
  CKBD0 U1559 ( .CLK(n1676), .C(n1677) );
  CKBD0 U1560 ( .CLK(n1677), .C(n1678) );
  CKBD0 U1561 ( .CLK(n1678), .C(n1679) );
  CKBD0 U1562 ( .CLK(n1679), .C(n1680) );
  BUFFD0 U1563 ( .I(n1680), .Z(n1681) );
  CKBD0 U1564 ( .CLK(n1681), .C(n1682) );
  CKBD0 U1565 ( .CLK(n1682), .C(n1683) );
  CKBD0 U1566 ( .CLK(n1683), .C(n1684) );
  CKBD0 U1567 ( .CLK(n1684), .C(n1685) );
  CKBD0 U1568 ( .CLK(n1685), .C(n1686) );
  CKBD0 U1569 ( .CLK(n1686), .C(n1687) );
  CKBD0 U1570 ( .CLK(n1687), .C(n1688) );
  CKBD0 U1571 ( .CLK(n1688), .C(n1689) );
  BUFFD0 U1572 ( .I(n8904), .Z(n1690) );
  CKBD0 U1573 ( .CLK(FrameSR[1]), .C(n1691) );
  CKBD0 U1574 ( .CLK(n1691), .C(n1692) );
  BUFFD0 U1575 ( .I(n8882), .Z(n1693) );
  CKBD0 U1576 ( .CLK(FrameSR[5]), .C(n1694) );
  CKBD0 U1577 ( .CLK(n1694), .C(n1695) );
  CKBD0 U1578 ( .CLK(n1695), .C(n1696) );
  BUFFD0 U1579 ( .I(n8417), .Z(n1697) );
  CKBD0 U1580 ( .CLK(FrameSR[17]), .C(n1698) );
  CKBD0 U1581 ( .CLK(n1698), .C(n1699) );
  CKBD0 U1582 ( .CLK(n1699), .C(n1700) );
  CKBD0 U1583 ( .CLK(n1700), .C(n1701) );
  CKBD0 U1584 ( .CLK(n1701), .C(n1702) );
  CKBD0 U1585 ( .CLK(n1702), .C(n1703) );
  CKBD0 U1586 ( .CLK(n1703), .C(n1704) );
  CKBD0 U1587 ( .CLK(n1704), .C(n1705) );
  CKBD0 U1588 ( .CLK(n1705), .C(n1706) );
  CKBD0 U1589 ( .CLK(n1706), .C(n1707) );
  BUFFD0 U1590 ( .I(n1707), .Z(n1708) );
  CKBD0 U1591 ( .CLK(n1708), .C(n1709) );
  CKBD0 U1592 ( .CLK(n1709), .C(n1710) );
  CKBD0 U1593 ( .CLK(n1710), .C(n1711) );
  CKBD0 U1594 ( .CLK(n1711), .C(n1712) );
  CKBD0 U1595 ( .CLK(n1712), .C(n1713) );
  CKBD0 U1596 ( .CLK(n1713), .C(n1714) );
  CKBD0 U1597 ( .CLK(n1714), .C(n1715) );
  CKBD0 U1598 ( .CLK(n1715), .C(n1716) );
  CKBD0 U1599 ( .CLK(n1716), .C(n1717) );
  CKBD0 U1600 ( .CLK(n1717), .C(n1718) );
  BUFFD0 U1601 ( .I(n1718), .Z(n1719) );
  CKBD0 U1602 ( .CLK(n1719), .C(n1720) );
  CKBD0 U1603 ( .CLK(n1720), .C(n1721) );
  CKBD0 U1604 ( .CLK(n1721), .C(n1722) );
  CKBD0 U1605 ( .CLK(n1722), .C(n1723) );
  CKBD0 U1606 ( .CLK(n1723), .C(n1724) );
  CKBD0 U1607 ( .CLK(n1724), .C(n1725) );
  CKBD0 U1608 ( .CLK(n1725), .C(n1726) );
  CKBD0 U1609 ( .CLK(n1726), .C(n1727) );
  CKBD0 U1610 ( .CLK(n1727), .C(n1728) );
  BUFFD0 U1611 ( .I(n1728), .Z(n1729) );
  CKBD0 U1612 ( .CLK(n1729), .C(n1730) );
  CKBD0 U1613 ( .CLK(n1730), .C(n1731) );
  CKBD0 U1614 ( .CLK(n1731), .C(n1732) );
  CKBD0 U1615 ( .CLK(n1732), .C(n1733) );
  CKBD0 U1616 ( .CLK(n1733), .C(n1734) );
  CKBD0 U1617 ( .CLK(n1734), .C(n1735) );
  CKBD0 U1618 ( .CLK(n1735), .C(n1736) );
  CKBD0 U1619 ( .CLK(n1736), .C(n1737) );
  CKBD0 U1620 ( .CLK(n1737), .C(n1738) );
  CKBD0 U1621 ( .CLK(n1738), .C(n1739) );
  BUFFD0 U1622 ( .I(n1739), .Z(n1740) );
  CKBD0 U1623 ( .CLK(n1740), .C(n1741) );
  CKBD0 U1624 ( .CLK(n1741), .C(n1742) );
  CKBD0 U1625 ( .CLK(n1742), .C(n1743) );
  CKBD0 U1626 ( .CLK(n1743), .C(n1744) );
  CKBD0 U1627 ( .CLK(n1744), .C(n1745) );
  CKBD0 U1628 ( .CLK(n1745), .C(n1746) );
  CKBD0 U1629 ( .CLK(n1746), .C(n1747) );
  CKBD0 U1630 ( .CLK(n1747), .C(n1748) );
  CKBD0 U1631 ( .CLK(n1748), .C(n1749) );
  CKBD0 U1632 ( .CLK(n1749), .C(n1750) );
  BUFFD0 U1633 ( .I(n1750), .Z(n1751) );
  CKBD0 U1634 ( .CLK(n1751), .C(n1752) );
  CKBD0 U1635 ( .CLK(n1752), .C(n1753) );
  CKBD0 U1636 ( .CLK(n1753), .C(n1754) );
  CKBD0 U1637 ( .CLK(n1754), .C(n1755) );
  CKBD0 U1638 ( .CLK(n1755), .C(n1756) );
  CKBD0 U1639 ( .CLK(n1756), .C(n1757) );
  CKBD0 U1640 ( .CLK(n1757), .C(n1758) );
  CKBD0 U1641 ( .CLK(n1758), .C(n1759) );
  CKBD0 U1642 ( .CLK(n1759), .C(n1760) );
  CKBD0 U1643 ( .CLK(n1760), .C(n1761) );
  BUFFD0 U1644 ( .I(n1761), .Z(n1762) );
  CKBD0 U1645 ( .CLK(n1762), .C(n1763) );
  CKBD0 U1646 ( .CLK(n1763), .C(n1764) );
  CKBD0 U1647 ( .CLK(n1764), .C(n1765) );
  CKBD0 U1648 ( .CLK(n1765), .C(n1766) );
  CKBD0 U1649 ( .CLK(n1766), .C(n1767) );
  CKBD0 U1650 ( .CLK(n1767), .C(n1768) );
  CKBD0 U1651 ( .CLK(n1768), .C(n1769) );
  CKBD0 U1652 ( .CLK(n1769), .C(n1770) );
  CKBD0 U1653 ( .CLK(n1770), .C(n1771) );
  CKBD0 U1654 ( .CLK(n1771), .C(n1772) );
  BUFFD0 U1655 ( .I(n1772), .Z(n1773) );
  CKBD0 U1656 ( .CLK(n1773), .C(n1774) );
  CKBD0 U1657 ( .CLK(n1774), .C(n1775) );
  CKBD0 U1658 ( .CLK(n1775), .C(n1776) );
  CKBD0 U1659 ( .CLK(n1776), .C(n1777) );
  CKBD0 U1660 ( .CLK(n1777), .C(n1778) );
  CKBD0 U1661 ( .CLK(n1778), .C(n1779) );
  CKBD0 U1662 ( .CLK(n1779), .C(n1780) );
  CKBD0 U1663 ( .CLK(n1780), .C(n1781) );
  CKBD0 U1664 ( .CLK(n1781), .C(n1782) );
  CKBD0 U1665 ( .CLK(n1782), .C(n1783) );
  BUFFD0 U1666 ( .I(n1783), .Z(n1784) );
  CKBD0 U1667 ( .CLK(n1784), .C(n1785) );
  CKBD0 U1668 ( .CLK(n1785), .C(n1786) );
  CKBD0 U1669 ( .CLK(n1786), .C(n1787) );
  CKBD0 U1670 ( .CLK(n1787), .C(n1788) );
  CKBD0 U1671 ( .CLK(n1788), .C(n1789) );
  CKBD0 U1672 ( .CLK(n1789), .C(n1790) );
  CKBD0 U1673 ( .CLK(n1790), .C(n1791) );
  CKBD0 U1674 ( .CLK(n1791), .C(n1792) );
  CKBD0 U1675 ( .CLK(n1792), .C(n1793) );
  CKBD0 U1676 ( .CLK(n1793), .C(n1794) );
  CKBD0 U1677 ( .CLK(n1794), .C(n1795) );
  BUFFD0 U1678 ( .I(n8808), .Z(n1796) );
  CKBD0 U1679 ( .CLK(FrameSR[32]), .C(n1797) );
  CKBD0 U1680 ( .CLK(n1797), .C(n1798) );
  CKBD0 U1681 ( .CLK(n1798), .C(n1799) );
  CKBD0 U1682 ( .CLK(n1799), .C(n1800) );
  CKBD0 U1683 ( .CLK(n1800), .C(n1801) );
  BUFFD0 U1684 ( .I(n1801), .Z(n1802) );
  CKBD0 U1685 ( .CLK(n1802), .C(n1803) );
  CKBD0 U1686 ( .CLK(n1803), .C(n1804) );
  CKBD0 U1687 ( .CLK(n1804), .C(n1805) );
  CKBD0 U1688 ( .CLK(n1805), .C(n1806) );
  CKBD0 U1689 ( .CLK(n1806), .C(n1807) );
  CKBD0 U1690 ( .CLK(n1807), .C(n1808) );
  CKBD0 U1691 ( .CLK(n1808), .C(n1809) );
  CKBD0 U1692 ( .CLK(n1809), .C(n1810) );
  CKBD0 U1693 ( .CLK(n1810), .C(n1811) );
  CKBD0 U1694 ( .CLK(n1811), .C(n1812) );
  BUFFD0 U1695 ( .I(n1812), .Z(n1813) );
  CKBD0 U1696 ( .CLK(n1813), .C(n1814) );
  CKBD0 U1697 ( .CLK(n1814), .C(n1815) );
  CKBD0 U1698 ( .CLK(n1815), .C(n1816) );
  CKBD0 U1699 ( .CLK(n1816), .C(n1817) );
  CKBD0 U1700 ( .CLK(n1817), .C(n1818) );
  CKBD0 U1701 ( .CLK(n1818), .C(n1819) );
  CKBD0 U1702 ( .CLK(n1819), .C(n1820) );
  CKBD0 U1703 ( .CLK(n1820), .C(n1821) );
  CKBD0 U1704 ( .CLK(n1821), .C(n1822) );
  BUFFD0 U1705 ( .I(n1822), .Z(n1823) );
  CKBD0 U1706 ( .CLK(n1823), .C(n1824) );
  CKBD0 U1707 ( .CLK(n1824), .C(n1825) );
  CKBD0 U1708 ( .CLK(n1825), .C(n1826) );
  CKBD0 U1709 ( .CLK(n1826), .C(n1827) );
  CKBD0 U1710 ( .CLK(n1827), .C(n1828) );
  CKBD0 U1711 ( .CLK(n1828), .C(n1829) );
  CKBD0 U1712 ( .CLK(n1829), .C(n1830) );
  CKBD0 U1713 ( .CLK(n1830), .C(n1831) );
  CKBD0 U1714 ( .CLK(n1831), .C(n1832) );
  CKBD0 U1715 ( .CLK(n1832), .C(n1833) );
  BUFFD0 U1716 ( .I(n1833), .Z(n1834) );
  CKBD0 U1717 ( .CLK(n1834), .C(n1835) );
  CKBD0 U1718 ( .CLK(n1835), .C(n1836) );
  CKBD0 U1719 ( .CLK(n1836), .C(n1837) );
  CKBD0 U1720 ( .CLK(n1837), .C(n1838) );
  CKBD0 U1721 ( .CLK(n1838), .C(n1839) );
  CKBD0 U1722 ( .CLK(n1839), .C(n1840) );
  CKBD0 U1723 ( .CLK(n1840), .C(n1841) );
  CKBD0 U1724 ( .CLK(n1841), .C(n1842) );
  CKBD0 U1725 ( .CLK(n1842), .C(n1843) );
  CKBD0 U1726 ( .CLK(n1843), .C(n1844) );
  BUFFD0 U1727 ( .I(n1844), .Z(n1845) );
  CKBD0 U1728 ( .CLK(n1845), .C(n1846) );
  CKBD0 U1729 ( .CLK(n1846), .C(n1847) );
  CKBD0 U1730 ( .CLK(n1847), .C(n1848) );
  CKBD0 U1731 ( .CLK(n1848), .C(n1849) );
  CKBD0 U1732 ( .CLK(n1849), .C(n1850) );
  CKBD0 U1733 ( .CLK(n1850), .C(n1851) );
  CKBD0 U1734 ( .CLK(n1851), .C(n1852) );
  CKBD0 U1735 ( .CLK(n1852), .C(n1853) );
  CKBD0 U1736 ( .CLK(n1853), .C(n1854) );
  CKBD0 U1737 ( .CLK(n1854), .C(n1855) );
  BUFFD0 U1738 ( .I(n1855), .Z(n1856) );
  CKBD0 U1739 ( .CLK(n1856), .C(n1857) );
  CKBD0 U1740 ( .CLK(n1857), .C(n1858) );
  CKBD0 U1741 ( .CLK(n1858), .C(n1859) );
  CKBD0 U1742 ( .CLK(n1859), .C(n1860) );
  CKBD0 U1743 ( .CLK(n1860), .C(n1861) );
  CKBD0 U1744 ( .CLK(n1861), .C(n1862) );
  CKBD0 U1745 ( .CLK(n1862), .C(n1863) );
  CKBD0 U1746 ( .CLK(n1863), .C(n1864) );
  CKBD0 U1747 ( .CLK(n1864), .C(n1865) );
  CKBD0 U1748 ( .CLK(n1865), .C(n1866) );
  BUFFD0 U1749 ( .I(n1866), .Z(n1867) );
  CKBD0 U1750 ( .CLK(n1867), .C(n1868) );
  CKBD0 U1751 ( .CLK(n1868), .C(n1869) );
  CKBD0 U1752 ( .CLK(n1869), .C(n1870) );
  CKBD0 U1753 ( .CLK(n1870), .C(n1871) );
  CKBD0 U1754 ( .CLK(n1871), .C(n1872) );
  CKBD0 U1755 ( .CLK(n1872), .C(n1873) );
  CKBD0 U1756 ( .CLK(n1873), .C(n1874) );
  CKBD0 U1757 ( .CLK(n1874), .C(n1875) );
  CKBD0 U1758 ( .CLK(n1875), .C(n1876) );
  CKBD0 U1759 ( .CLK(n1876), .C(n1877) );
  BUFFD0 U1760 ( .I(n1877), .Z(n1878) );
  CKBD0 U1761 ( .CLK(n1878), .C(n1879) );
  CKBD0 U1762 ( .CLK(n1879), .C(n1880) );
  CKBD0 U1763 ( .CLK(n1880), .C(n1881) );
  CKBD0 U1764 ( .CLK(n1881), .C(n1882) );
  CKBD0 U1765 ( .CLK(n1882), .C(n1883) );
  CKBD0 U1766 ( .CLK(n1883), .C(n1884) );
  CKBD0 U1767 ( .CLK(n1884), .C(n1885) );
  CKBD0 U1768 ( .CLK(n1885), .C(n1886) );
  CKBD0 U1769 ( .CLK(n1886), .C(n1887) );
  CKBD0 U1770 ( .CLK(n1887), .C(n1888) );
  BUFFD0 U1771 ( .I(n1888), .Z(n1889) );
  CKBD0 U1772 ( .CLK(n1889), .C(n1890) );
  CKBD0 U1773 ( .CLK(n1890), .C(n1891) );
  CKBD0 U1774 ( .CLK(n1891), .C(n1892) );
  CKBD0 U1775 ( .CLK(n1892), .C(n1893) );
  CKBD0 U1776 ( .CLK(n1893), .C(n1894) );
  CKBD0 U1777 ( .CLK(n1894), .C(n1895) );
  BUFFD0 U1778 ( .I(n3828), .Z(n1896) );
  CKBD0 U1779 ( .CLK(FrameSR[47]), .C(n1897) );
  BUFFD0 U1780 ( .I(n8879), .Z(n1898) );
  CKBD0 U1781 ( .CLK(FrameSR[0]), .C(n1899) );
  CKBD0 U1782 ( .CLK(n1899), .C(n1900) );
  BUFFD0 U1783 ( .I(n8922), .Z(n1901) );
  CKBD0 U1784 ( .CLK(FrameSR[2]), .C(n1902) );
  CKBD0 U1785 ( .CLK(n1902), .C(n1903) );
  BUFFD0 U1786 ( .I(n8880), .Z(n1904) );
  CKBD0 U1787 ( .CLK(FrameSR[4]), .C(n1905) );
  CKBD0 U1788 ( .CLK(n1905), .C(n1906) );
  BUFFD0 U1789 ( .I(n8971), .Z(n1907) );
  CKBD0 U1790 ( .CLK(FrameSR[6]), .C(n1908) );
  CKBD0 U1791 ( .CLK(n1908), .C(n1909) );
  CKBD0 U1792 ( .CLK(n1909), .C(n1910) );
  BUFFD0 U1793 ( .I(n8182), .Z(n1911) );
  CKBD0 U1794 ( .CLK(FrameSR[20]), .C(n1912) );
  CKBD0 U1795 ( .CLK(n1912), .C(n1913) );
  CKBD0 U1796 ( .CLK(n1913), .C(n1914) );
  CKBD0 U1797 ( .CLK(n1914), .C(n1915) );
  CKBD0 U1798 ( .CLK(n1915), .C(n1916) );
  CKBD0 U1799 ( .CLK(n1916), .C(n1917) );
  BUFFD0 U1800 ( .I(n1917), .Z(n1918) );
  CKBD0 U1801 ( .CLK(n1918), .C(n1919) );
  CKBD0 U1802 ( .CLK(n1919), .C(n1920) );
  CKBD0 U1803 ( .CLK(n1920), .C(n1921) );
  CKBD0 U1804 ( .CLK(n1921), .C(n1922) );
  CKBD0 U1805 ( .CLK(n1922), .C(n1923) );
  CKBD0 U1806 ( .CLK(n1923), .C(n1924) );
  CKBD0 U1807 ( .CLK(n1924), .C(n1925) );
  CKBD0 U1808 ( .CLK(n1925), .C(n1926) );
  CKBD0 U1809 ( .CLK(n1926), .C(n1927) );
  CKBD0 U1810 ( .CLK(n1927), .C(n1928) );
  BUFFD0 U1811 ( .I(n1928), .Z(n1929) );
  CKBD0 U1812 ( .CLK(n1929), .C(n1930) );
  CKBD0 U1813 ( .CLK(n1930), .C(n1931) );
  CKBD0 U1814 ( .CLK(n1931), .C(n1932) );
  CKBD0 U1815 ( .CLK(n1932), .C(n1933) );
  CKBD0 U1816 ( .CLK(n1933), .C(n1934) );
  CKBD0 U1817 ( .CLK(n1934), .C(n1935) );
  CKBD0 U1818 ( .CLK(n1935), .C(n1936) );
  CKBD0 U1819 ( .CLK(n1936), .C(n1937) );
  CKBD0 U1820 ( .CLK(n1937), .C(n1938) );
  CKBD0 U1821 ( .CLK(n1938), .C(n1939) );
  BUFFD0 U1822 ( .I(n1939), .Z(n1940) );
  CKBD0 U1823 ( .CLK(n1940), .C(n1941) );
  CKBD0 U1824 ( .CLK(n1941), .C(n1942) );
  CKBD0 U1825 ( .CLK(n1942), .C(n1943) );
  CKBD0 U1826 ( .CLK(n1943), .C(n1944) );
  CKBD0 U1827 ( .CLK(n1944), .C(n1945) );
  CKBD0 U1828 ( .CLK(n1945), .C(n1946) );
  CKBD0 U1829 ( .CLK(n1946), .C(n1947) );
  CKBD0 U1830 ( .CLK(n1947), .C(n1948) );
  CKBD0 U1831 ( .CLK(n1948), .C(n1949) );
  CKBD0 U1832 ( .CLK(n1949), .C(n1950) );
  BUFFD0 U1833 ( .I(n1950), .Z(n1951) );
  CKBD0 U1834 ( .CLK(n1951), .C(n1952) );
  CKBD0 U1835 ( .CLK(n1952), .C(n1953) );
  CKBD0 U1836 ( .CLK(n1953), .C(n1954) );
  CKBD0 U1837 ( .CLK(n1954), .C(n1955) );
  CKBD0 U1838 ( .CLK(n1955), .C(n1956) );
  CKBD0 U1839 ( .CLK(n1956), .C(n1957) );
  CKBD0 U1840 ( .CLK(n1957), .C(n1958) );
  CKBD0 U1841 ( .CLK(n1958), .C(n1959) );
  CKBD0 U1842 ( .CLK(n1959), .C(n1960) );
  BUFFD0 U1843 ( .I(n1960), .Z(n1961) );
  CKBD0 U1844 ( .CLK(n1961), .C(n1962) );
  CKBD0 U1845 ( .CLK(n1962), .C(n1963) );
  CKBD0 U1846 ( .CLK(n1963), .C(n1964) );
  CKBD0 U1847 ( .CLK(n1964), .C(n1965) );
  CKBD0 U1848 ( .CLK(n1965), .C(n1966) );
  CKBD0 U1849 ( .CLK(n1966), .C(n1967) );
  CKBD0 U1850 ( .CLK(n1967), .C(n1968) );
  CKBD0 U1851 ( .CLK(n1968), .C(n1969) );
  CKBD0 U1852 ( .CLK(n1969), .C(n1970) );
  CKBD0 U1853 ( .CLK(n1970), .C(n1971) );
  BUFFD0 U1854 ( .I(n1971), .Z(n1972) );
  CKBD0 U1855 ( .CLK(n1972), .C(n1973) );
  CKBD0 U1856 ( .CLK(n1973), .C(n1974) );
  CKBD0 U1857 ( .CLK(n1974), .C(n1975) );
  CKBD0 U1858 ( .CLK(n1975), .C(n1976) );
  CKBD0 U1859 ( .CLK(n1976), .C(n1977) );
  CKBD0 U1860 ( .CLK(n1977), .C(n1978) );
  CKBD0 U1861 ( .CLK(n1978), .C(n1979) );
  CKBD0 U1862 ( .CLK(n1979), .C(n1980) );
  CKBD0 U1863 ( .CLK(n1980), .C(n1981) );
  CKBD0 U1864 ( .CLK(n1981), .C(n1982) );
  BUFFD0 U1865 ( .I(n1982), .Z(n1983) );
  CKBD0 U1866 ( .CLK(n1983), .C(n1984) );
  CKBD0 U1867 ( .CLK(n1984), .C(n1985) );
  CKBD0 U1868 ( .CLK(n1985), .C(n1986) );
  CKBD0 U1869 ( .CLK(n1986), .C(n1987) );
  CKBD0 U1870 ( .CLK(n1987), .C(n1988) );
  CKBD0 U1871 ( .CLK(n1988), .C(n1989) );
  CKBD0 U1872 ( .CLK(n1989), .C(n1990) );
  CKBD0 U1873 ( .CLK(n1990), .C(n1991) );
  CKBD0 U1874 ( .CLK(n1991), .C(n1992) );
  CKBD0 U1875 ( .CLK(n1992), .C(n1993) );
  BUFFD0 U1876 ( .I(n1993), .Z(n1994) );
  CKBD0 U1877 ( .CLK(n1994), .C(n1995) );
  CKBD0 U1878 ( .CLK(n1995), .C(n1996) );
  CKBD0 U1879 ( .CLK(n1996), .C(n1997) );
  CKBD0 U1880 ( .CLK(n1997), .C(n1998) );
  CKBD0 U1881 ( .CLK(n1998), .C(n1999) );
  CKBD0 U1882 ( .CLK(n1999), .C(n2000) );
  CKBD0 U1883 ( .CLK(n2000), .C(n2001) );
  CKBD0 U1884 ( .CLK(n2001), .C(n2002) );
  CKBD0 U1885 ( .CLK(n2002), .C(n2003) );
  CKBD0 U1886 ( .CLK(n2003), .C(n2004) );
  BUFFD0 U1887 ( .I(n2004), .Z(n2005) );
  CKBD0 U1888 ( .CLK(n2005), .C(n2006) );
  CKBD0 U1889 ( .CLK(n2006), .C(n2007) );
  CKBD0 U1890 ( .CLK(n2007), .C(n2008) );
  CKBD0 U1891 ( .CLK(n2008), .C(n2009) );
  BUFFD0 U1892 ( .I(n8444), .Z(n2010) );
  CKBD0 U1893 ( .CLK(FrameSR[34]), .C(n2011) );
  CKBD0 U1894 ( .CLK(n2011), .C(n2012) );
  CKBD0 U1895 ( .CLK(n2012), .C(n2013) );
  CKBD0 U1896 ( .CLK(n2013), .C(n2014) );
  BUFFD0 U1897 ( .I(n2014), .Z(n2015) );
  CKBD0 U1898 ( .CLK(n2015), .C(n2016) );
  CKBD0 U1899 ( .CLK(n2016), .C(n2017) );
  CKBD0 U1900 ( .CLK(n2017), .C(n2018) );
  CKBD0 U1901 ( .CLK(n2018), .C(n2019) );
  CKBD0 U1902 ( .CLK(n2019), .C(n2020) );
  CKBD0 U1903 ( .CLK(n2020), .C(n2021) );
  CKBD0 U1904 ( .CLK(n2021), .C(n2022) );
  CKBD0 U1905 ( .CLK(n2022), .C(n2023) );
  CKBD0 U1906 ( .CLK(n2023), .C(n2024) );
  CKBD0 U1907 ( .CLK(n2024), .C(n2025) );
  BUFFD0 U1908 ( .I(n2025), .Z(n2026) );
  CKBD0 U1909 ( .CLK(n2026), .C(n2027) );
  CKBD0 U1910 ( .CLK(n2027), .C(n2028) );
  CKBD0 U1911 ( .CLK(n2028), .C(n2029) );
  CKBD0 U1912 ( .CLK(n2029), .C(n2030) );
  CKBD0 U1913 ( .CLK(n2030), .C(n2031) );
  CKBD0 U1914 ( .CLK(n2031), .C(n2032) );
  CKBD0 U1915 ( .CLK(n2032), .C(n2033) );
  CKBD0 U1916 ( .CLK(n2033), .C(n2034) );
  CKBD0 U1917 ( .CLK(n2034), .C(n2035) );
  CKBD0 U1918 ( .CLK(n2035), .C(n2036) );
  BUFFD0 U1919 ( .I(n2036), .Z(n2037) );
  CKBD0 U1920 ( .CLK(n2037), .C(n2038) );
  CKBD0 U1921 ( .CLK(n2038), .C(n2039) );
  CKBD0 U1922 ( .CLK(n2039), .C(n2040) );
  CKBD0 U1923 ( .CLK(n2040), .C(n2041) );
  CKBD0 U1924 ( .CLK(n2041), .C(n2042) );
  CKBD0 U1925 ( .CLK(n2042), .C(n2043) );
  CKBD0 U1926 ( .CLK(n2043), .C(n2044) );
  CKBD0 U1927 ( .CLK(n2044), .C(n2045) );
  CKBD0 U1928 ( .CLK(n2045), .C(n2046) );
  BUFFD0 U1929 ( .I(n2046), .Z(n2047) );
  CKBD0 U1930 ( .CLK(n2047), .C(n2048) );
  CKBD0 U1931 ( .CLK(n2048), .C(n2049) );
  CKBD0 U1932 ( .CLK(n2049), .C(n2050) );
  CKBD0 U1933 ( .CLK(n2050), .C(n2051) );
  CKBD0 U1934 ( .CLK(n2051), .C(n2052) );
  CKBD0 U1935 ( .CLK(n2052), .C(n2053) );
  CKBD0 U1936 ( .CLK(n2053), .C(n2054) );
  CKBD0 U1937 ( .CLK(n2054), .C(n2055) );
  CKBD0 U1938 ( .CLK(n2055), .C(n2056) );
  CKBD0 U1939 ( .CLK(n2056), .C(n2057) );
  BUFFD0 U1940 ( .I(n2057), .Z(n2058) );
  CKBD0 U1941 ( .CLK(n2058), .C(n2059) );
  CKBD0 U1942 ( .CLK(n2059), .C(n2060) );
  CKBD0 U1943 ( .CLK(n2060), .C(n2061) );
  CKBD0 U1944 ( .CLK(n2061), .C(n2062) );
  CKBD0 U1945 ( .CLK(n2062), .C(n2063) );
  CKBD0 U1946 ( .CLK(n2063), .C(n2064) );
  CKBD0 U1947 ( .CLK(n2064), .C(n2065) );
  CKBD0 U1948 ( .CLK(n2065), .C(n2066) );
  CKBD0 U1949 ( .CLK(n2066), .C(n2067) );
  CKBD0 U1950 ( .CLK(n2067), .C(n2068) );
  BUFFD0 U1951 ( .I(n2068), .Z(n2069) );
  CKBD0 U1952 ( .CLK(n2069), .C(n2070) );
  CKBD0 U1953 ( .CLK(n2070), .C(n2071) );
  CKBD0 U1954 ( .CLK(n2071), .C(n2072) );
  CKBD0 U1955 ( .CLK(n2072), .C(n2073) );
  CKBD0 U1956 ( .CLK(n2073), .C(n2074) );
  CKBD0 U1957 ( .CLK(n2074), .C(n2075) );
  CKBD0 U1958 ( .CLK(n2075), .C(n2076) );
  CKBD0 U1959 ( .CLK(n2076), .C(n2077) );
  CKBD0 U1960 ( .CLK(n2077), .C(n2078) );
  CKBD0 U1961 ( .CLK(n2078), .C(n2079) );
  BUFFD0 U1962 ( .I(n2079), .Z(n2080) );
  CKBD0 U1963 ( .CLK(n2080), .C(n2081) );
  CKBD0 U1964 ( .CLK(n2081), .C(n2082) );
  CKBD0 U1965 ( .CLK(n2082), .C(n2083) );
  CKBD0 U1966 ( .CLK(n2083), .C(n2084) );
  CKBD0 U1967 ( .CLK(n2084), .C(n2085) );
  CKBD0 U1968 ( .CLK(n2085), .C(n2086) );
  CKBD0 U1969 ( .CLK(n2086), .C(n2087) );
  CKBD0 U1970 ( .CLK(n2087), .C(n2088) );
  CKBD0 U1971 ( .CLK(n2088), .C(n2089) );
  CKBD0 U1972 ( .CLK(n2089), .C(n2090) );
  BUFFD0 U1973 ( .I(n2090), .Z(n2091) );
  CKBD0 U1974 ( .CLK(n2091), .C(n2092) );
  CKBD0 U1975 ( .CLK(n2092), .C(n2093) );
  CKBD0 U1976 ( .CLK(n2093), .C(n2094) );
  CKBD0 U1977 ( .CLK(n2094), .C(n2095) );
  CKBD0 U1978 ( .CLK(n2095), .C(n2096) );
  CKBD0 U1979 ( .CLK(n2096), .C(n2097) );
  CKBD0 U1980 ( .CLK(n2097), .C(n2098) );
  CKBD0 U1981 ( .CLK(n2098), .C(n2099) );
  CKBD0 U1982 ( .CLK(n2099), .C(n2100) );
  CKBD0 U1983 ( .CLK(n2100), .C(n2101) );
  BUFFD0 U1984 ( .I(n2101), .Z(n2102) );
  CKBD0 U1985 ( .CLK(n2102), .C(n2103) );
  CKBD0 U1986 ( .CLK(n2103), .C(n2104) );
  CKBD0 U1987 ( .CLK(n2104), .C(n2105) );
  CKBD0 U1988 ( .CLK(n2105), .C(n2106) );
  CKBD0 U1989 ( .CLK(n2106), .C(n2107) );
  CKBD0 U1990 ( .CLK(n2107), .C(n2108) );
  BUFFD0 U1991 ( .I(n8330), .Z(n2109) );
  CKBD0 U1992 ( .CLK(FrameSR[49]), .C(n2110) );
  CKBD0 U1993 ( .CLK(n2110), .C(n2111) );
  CKBD0 U1994 ( .CLK(n2111), .C(n2112) );
  CKBD0 U1995 ( .CLK(n2112), .C(n2113) );
  CKBD0 U1996 ( .CLK(n2113), .C(n2114) );
  CKBD0 U1997 ( .CLK(n2114), .C(n2115) );
  BUFFD0 U1998 ( .I(n2115), .Z(n2116) );
  CKBD0 U1999 ( .CLK(n2116), .C(n2117) );
  CKBD0 U2000 ( .CLK(n2117), .C(n2118) );
  CKBD0 U2001 ( .CLK(n2118), .C(n2119) );
  CKBD0 U2002 ( .CLK(n2119), .C(n2120) );
  CKBD0 U2003 ( .CLK(n2120), .C(n2121) );
  CKBD0 U2004 ( .CLK(n2121), .C(n2122) );
  CKBD0 U2005 ( .CLK(n2122), .C(n2123) );
  CKBD0 U2006 ( .CLK(n2123), .C(n2124) );
  CKBD0 U2007 ( .CLK(n2124), .C(n2125) );
  CKBD0 U2008 ( .CLK(n2125), .C(n2126) );
  BUFFD0 U2009 ( .I(n2126), .Z(n2127) );
  CKBD0 U2010 ( .CLK(n2127), .C(n2128) );
  CKBD0 U2011 ( .CLK(n2128), .C(n2129) );
  CKBD0 U2012 ( .CLK(n2129), .C(n2130) );
  CKBD0 U2013 ( .CLK(n2130), .C(n2131) );
  CKBD0 U2014 ( .CLK(n2131), .C(n2132) );
  CKBD0 U2015 ( .CLK(n2132), .C(n2133) );
  CKBD0 U2016 ( .CLK(n2133), .C(n2134) );
  CKBD0 U2017 ( .CLK(n2134), .C(n2135) );
  CKBD0 U2018 ( .CLK(n2135), .C(n2136) );
  CKBD0 U2019 ( .CLK(n2136), .C(n2137) );
  BUFFD0 U2020 ( .I(n2137), .Z(n2138) );
  CKBD0 U2021 ( .CLK(n2138), .C(n2139) );
  CKBD0 U2022 ( .CLK(n2139), .C(n2140) );
  CKBD0 U2023 ( .CLK(n2140), .C(n2141) );
  CKBD0 U2024 ( .CLK(n2141), .C(n2142) );
  CKBD0 U2025 ( .CLK(n2142), .C(n2143) );
  CKBD0 U2026 ( .CLK(n2143), .C(n2144) );
  CKBD0 U2027 ( .CLK(n2144), .C(n2145) );
  CKBD0 U2028 ( .CLK(n2145), .C(n2146) );
  CKBD0 U2029 ( .CLK(n2146), .C(n2147) );
  CKBD0 U2030 ( .CLK(n2147), .C(n2148) );
  BUFFD0 U2031 ( .I(n2148), .Z(n2149) );
  CKBD0 U2032 ( .CLK(n2149), .C(n2150) );
  CKBD0 U2033 ( .CLK(n2150), .C(n2151) );
  CKBD0 U2034 ( .CLK(n2151), .C(n2152) );
  CKBD0 U2035 ( .CLK(n2152), .C(n2153) );
  CKBD0 U2036 ( .CLK(n2153), .C(n2154) );
  CKBD0 U2037 ( .CLK(n2154), .C(n2155) );
  CKBD0 U2038 ( .CLK(n2155), .C(n2156) );
  CKBD0 U2039 ( .CLK(n2156), .C(n2157) );
  CKBD0 U2040 ( .CLK(n2157), .C(n2158) );
  BUFFD0 U2041 ( .I(n2158), .Z(n2159) );
  CKBD0 U2042 ( .CLK(n2159), .C(n2160) );
  CKBD0 U2043 ( .CLK(n2160), .C(n2161) );
  CKBD0 U2044 ( .CLK(n2161), .C(n2162) );
  CKBD0 U2045 ( .CLK(n2162), .C(n2163) );
  CKBD0 U2046 ( .CLK(n2163), .C(n2164) );
  CKBD0 U2047 ( .CLK(n2164), .C(n2165) );
  CKBD0 U2048 ( .CLK(n2165), .C(n2166) );
  CKBD0 U2049 ( .CLK(n2166), .C(n2167) );
  CKBD0 U2050 ( .CLK(n2167), .C(n2168) );
  CKBD0 U2051 ( .CLK(n2168), .C(n2169) );
  BUFFD0 U2052 ( .I(n2169), .Z(n2170) );
  CKBD0 U2053 ( .CLK(n2170), .C(n2171) );
  CKBD0 U2054 ( .CLK(n2171), .C(n2172) );
  CKBD0 U2055 ( .CLK(n2172), .C(n2173) );
  CKBD0 U2056 ( .CLK(n2173), .C(n2174) );
  CKBD0 U2057 ( .CLK(n2174), .C(n2175) );
  CKBD0 U2058 ( .CLK(n2175), .C(n2176) );
  CKBD0 U2059 ( .CLK(n2176), .C(n2177) );
  CKBD0 U2060 ( .CLK(n2177), .C(n2178) );
  CKBD0 U2061 ( .CLK(n2178), .C(n2179) );
  CKBD0 U2062 ( .CLK(n2179), .C(n2180) );
  BUFFD0 U2063 ( .I(n2180), .Z(n2181) );
  CKBD0 U2064 ( .CLK(n2181), .C(n2182) );
  CKBD0 U2065 ( .CLK(n2182), .C(n2183) );
  CKBD0 U2066 ( .CLK(n2183), .C(n2184) );
  CKBD0 U2067 ( .CLK(n2184), .C(n2185) );
  CKBD0 U2068 ( .CLK(n2185), .C(n2186) );
  CKBD0 U2069 ( .CLK(n2186), .C(n2187) );
  CKBD0 U2070 ( .CLK(n2187), .C(n2188) );
  CKBD0 U2071 ( .CLK(n2188), .C(n2189) );
  CKBD0 U2072 ( .CLK(n2189), .C(n2190) );
  CKBD0 U2073 ( .CLK(n2190), .C(n2191) );
  BUFFD0 U2074 ( .I(n2191), .Z(n2192) );
  CKBD0 U2075 ( .CLK(n2192), .C(n2193) );
  CKBD0 U2076 ( .CLK(n2193), .C(n2194) );
  CKBD0 U2077 ( .CLK(n2194), .C(n2195) );
  CKBD0 U2078 ( .CLK(n2195), .C(n2196) );
  CKBD0 U2079 ( .CLK(n2196), .C(n2197) );
  CKBD0 U2080 ( .CLK(n2197), .C(n2198) );
  CKBD0 U2081 ( .CLK(n2198), .C(n2199) );
  CKBD0 U2082 ( .CLK(n2199), .C(n2200) );
  CKBD0 U2083 ( .CLK(n2200), .C(n2201) );
  CKBD0 U2084 ( .CLK(n2201), .C(n2202) );
  BUFFD0 U2085 ( .I(n2202), .Z(n2203) );
  CKBD0 U2086 ( .CLK(n2203), .C(n2204) );
  CKBD0 U2087 ( .CLK(n2204), .C(n2205) );
  CKBD0 U2088 ( .CLK(n2205), .C(n2206) );
  CKBD0 U2089 ( .CLK(n2206), .C(n2207) );
  BUFFD0 U2090 ( .I(n8140), .Z(n2208) );
  CKBD0 U2091 ( .CLK(FrameSR[50]), .C(n2209) );
  CKBD0 U2092 ( .CLK(n2209), .C(n2210) );
  CKBD0 U2093 ( .CLK(n2210), .C(n2211) );
  CKBD0 U2094 ( .CLK(n2211), .C(n2212) );
  BUFFD0 U2095 ( .I(n2212), .Z(n2213) );
  CKBD0 U2096 ( .CLK(n2213), .C(n2214) );
  CKBD0 U2097 ( .CLK(n2214), .C(n2215) );
  CKBD0 U2098 ( .CLK(n2215), .C(n2216) );
  CKBD0 U2099 ( .CLK(n2216), .C(n2217) );
  CKBD0 U2100 ( .CLK(n2217), .C(n2218) );
  CKBD0 U2101 ( .CLK(n2218), .C(n2219) );
  CKBD0 U2102 ( .CLK(n2219), .C(n2220) );
  CKBD0 U2103 ( .CLK(n2220), .C(n2221) );
  CKBD0 U2104 ( .CLK(n2221), .C(n2222) );
  CKBD0 U2105 ( .CLK(n2222), .C(n2223) );
  BUFFD0 U2106 ( .I(n2223), .Z(n2224) );
  CKBD0 U2107 ( .CLK(n2224), .C(n2225) );
  CKBD0 U2108 ( .CLK(n2225), .C(n2226) );
  CKBD0 U2109 ( .CLK(n2226), .C(n2227) );
  CKBD0 U2110 ( .CLK(n2227), .C(n2228) );
  CKBD0 U2111 ( .CLK(n2228), .C(n2229) );
  CKBD0 U2112 ( .CLK(n2229), .C(n2230) );
  CKBD0 U2113 ( .CLK(n2230), .C(n2231) );
  CKBD0 U2114 ( .CLK(n2231), .C(n2232) );
  CKBD0 U2115 ( .CLK(n2232), .C(n2233) );
  CKBD0 U2116 ( .CLK(n2233), .C(n2234) );
  BUFFD0 U2117 ( .I(n2234), .Z(n2235) );
  CKBD0 U2118 ( .CLK(n2235), .C(n2236) );
  CKBD0 U2119 ( .CLK(n2236), .C(n2237) );
  CKBD0 U2120 ( .CLK(n2237), .C(n2238) );
  CKBD0 U2121 ( .CLK(n2238), .C(n2239) );
  CKBD0 U2122 ( .CLK(n2239), .C(n2240) );
  CKBD0 U2123 ( .CLK(n2240), .C(n2241) );
  CKBD0 U2124 ( .CLK(n2241), .C(n2242) );
  CKBD0 U2125 ( .CLK(n2242), .C(n2243) );
  CKBD0 U2126 ( .CLK(n2243), .C(n2244) );
  BUFFD0 U2127 ( .I(n2244), .Z(n2245) );
  CKBD0 U2128 ( .CLK(n2245), .C(n2246) );
  CKBD0 U2129 ( .CLK(n2246), .C(n2247) );
  CKBD0 U2130 ( .CLK(n2247), .C(n2248) );
  CKBD0 U2131 ( .CLK(n2248), .C(n2249) );
  CKBD0 U2132 ( .CLK(n2249), .C(n2250) );
  CKBD0 U2133 ( .CLK(n2250), .C(n2251) );
  CKBD0 U2134 ( .CLK(n2251), .C(n2252) );
  CKBD0 U2135 ( .CLK(n2252), .C(n2253) );
  CKBD0 U2136 ( .CLK(n2253), .C(n2254) );
  CKBD0 U2137 ( .CLK(n2254), .C(n2255) );
  BUFFD0 U2138 ( .I(n2255), .Z(n2256) );
  CKBD0 U2139 ( .CLK(n2256), .C(n2257) );
  CKBD0 U2140 ( .CLK(n2257), .C(n2258) );
  CKBD0 U2141 ( .CLK(n2258), .C(n2259) );
  CKBD0 U2142 ( .CLK(n2259), .C(n2260) );
  CKBD0 U2143 ( .CLK(n2260), .C(n2261) );
  CKBD0 U2144 ( .CLK(n2261), .C(n2262) );
  CKBD0 U2145 ( .CLK(n2262), .C(n2263) );
  CKBD0 U2146 ( .CLK(n2263), .C(n2264) );
  CKBD0 U2147 ( .CLK(n2264), .C(n2265) );
  CKBD0 U2148 ( .CLK(n2265), .C(n2266) );
  BUFFD0 U2149 ( .I(n2266), .Z(n2267) );
  CKBD0 U2150 ( .CLK(n2267), .C(n2268) );
  CKBD0 U2151 ( .CLK(n2268), .C(n2269) );
  CKBD0 U2152 ( .CLK(n2269), .C(n2270) );
  CKBD0 U2153 ( .CLK(n2270), .C(n2271) );
  CKBD0 U2154 ( .CLK(n2271), .C(n2272) );
  CKBD0 U2155 ( .CLK(n2272), .C(n2273) );
  CKBD0 U2156 ( .CLK(n2273), .C(n2274) );
  CKBD0 U2157 ( .CLK(n2274), .C(n2275) );
  CKBD0 U2158 ( .CLK(n2275), .C(n2276) );
  CKBD0 U2159 ( .CLK(n2276), .C(n2277) );
  BUFFD0 U2160 ( .I(n2277), .Z(n2278) );
  CKBD0 U2161 ( .CLK(n2278), .C(n2279) );
  CKBD0 U2162 ( .CLK(n2279), .C(n2280) );
  CKBD0 U2163 ( .CLK(n2280), .C(n2281) );
  CKBD0 U2164 ( .CLK(n2281), .C(n2282) );
  CKBD0 U2165 ( .CLK(n2282), .C(n2283) );
  CKBD0 U2166 ( .CLK(n2283), .C(n2284) );
  CKBD0 U2167 ( .CLK(n2284), .C(n2285) );
  CKBD0 U2168 ( .CLK(n2285), .C(n2286) );
  CKBD0 U2169 ( .CLK(n2286), .C(n2287) );
  CKBD0 U2170 ( .CLK(n2287), .C(n2288) );
  BUFFD0 U2171 ( .I(n2288), .Z(n2289) );
  CKBD0 U2172 ( .CLK(n2289), .C(n2290) );
  CKBD0 U2173 ( .CLK(n2290), .C(n2291) );
  CKBD0 U2174 ( .CLK(n2291), .C(n2292) );
  CKBD0 U2175 ( .CLK(n2292), .C(n2293) );
  CKBD0 U2176 ( .CLK(n2293), .C(n2294) );
  CKBD0 U2177 ( .CLK(n2294), .C(n2295) );
  CKBD0 U2178 ( .CLK(n2295), .C(n2296) );
  CKBD0 U2179 ( .CLK(n2296), .C(n2297) );
  CKBD0 U2180 ( .CLK(n2297), .C(n2298) );
  CKBD0 U2181 ( .CLK(n2298), .C(n2299) );
  BUFFD0 U2182 ( .I(n2299), .Z(n2300) );
  CKBD0 U2183 ( .CLK(n2300), .C(n2301) );
  CKBD0 U2184 ( .CLK(n2301), .C(n2302) );
  CKBD0 U2185 ( .CLK(n2302), .C(n2303) );
  CKBD0 U2186 ( .CLK(n2303), .C(n2304) );
  CKBD0 U2187 ( .CLK(n2304), .C(n2305) );
  CKBD0 U2188 ( .CLK(n2305), .C(n2306) );
  BUFFD0 U2189 ( .I(n8335), .Z(n2307) );
  CKBD0 U2190 ( .CLK(FrameSR[35]), .C(n2308) );
  CKBD0 U2191 ( .CLK(n2308), .C(n2309) );
  CKBD0 U2192 ( .CLK(n2309), .C(n2310) );
  CKBD0 U2193 ( .CLK(n2310), .C(n2311) );
  CKBD0 U2194 ( .CLK(n2311), .C(n2312) );
  CKBD0 U2195 ( .CLK(n2312), .C(n2313) );
  BUFFD0 U2196 ( .I(n2313), .Z(n2314) );
  CKBD0 U2197 ( .CLK(n2314), .C(n2315) );
  CKBD0 U2198 ( .CLK(n2315), .C(n2316) );
  CKBD0 U2199 ( .CLK(n2316), .C(n2317) );
  CKBD0 U2200 ( .CLK(n2317), .C(n2318) );
  CKBD0 U2201 ( .CLK(n2318), .C(n2319) );
  CKBD0 U2202 ( .CLK(n2319), .C(n2320) );
  CKBD0 U2203 ( .CLK(n2320), .C(n2321) );
  CKBD0 U2204 ( .CLK(n2321), .C(n2322) );
  CKBD0 U2205 ( .CLK(n2322), .C(n2323) );
  CKBD0 U2206 ( .CLK(n2323), .C(n2324) );
  BUFFD0 U2207 ( .I(n2324), .Z(n2325) );
  CKBD0 U2208 ( .CLK(n2325), .C(n2326) );
  CKBD0 U2209 ( .CLK(n2326), .C(n2327) );
  CKBD0 U2210 ( .CLK(n2327), .C(n2328) );
  CKBD0 U2211 ( .CLK(n2328), .C(n2329) );
  CKBD0 U2212 ( .CLK(n2329), .C(n2330) );
  CKBD0 U2213 ( .CLK(n2330), .C(n2331) );
  CKBD0 U2214 ( .CLK(n2331), .C(n2332) );
  CKBD0 U2215 ( .CLK(n2332), .C(n2333) );
  CKBD0 U2216 ( .CLK(n2333), .C(n2334) );
  CKBD0 U2217 ( .CLK(n2334), .C(n2335) );
  BUFFD0 U2218 ( .I(n2335), .Z(n2336) );
  CKBD0 U2219 ( .CLK(n2336), .C(n2337) );
  CKBD0 U2220 ( .CLK(n2337), .C(n2338) );
  CKBD0 U2221 ( .CLK(n2338), .C(n2339) );
  CKBD0 U2222 ( .CLK(n2339), .C(n2340) );
  CKBD0 U2223 ( .CLK(n2340), .C(n2341) );
  CKBD0 U2224 ( .CLK(n2341), .C(n2342) );
  CKBD0 U2225 ( .CLK(n2342), .C(n2343) );
  CKBD0 U2226 ( .CLK(n2343), .C(n2344) );
  CKBD0 U2227 ( .CLK(n2344), .C(n2345) );
  CKBD0 U2228 ( .CLK(n2345), .C(n2346) );
  BUFFD0 U2229 ( .I(n2346), .Z(n2347) );
  CKBD0 U2230 ( .CLK(n2347), .C(n2348) );
  CKBD0 U2231 ( .CLK(n2348), .C(n2349) );
  CKBD0 U2232 ( .CLK(n2349), .C(n2350) );
  CKBD0 U2233 ( .CLK(n2350), .C(n2351) );
  CKBD0 U2234 ( .CLK(n2351), .C(n2352) );
  CKBD0 U2235 ( .CLK(n2352), .C(n2353) );
  CKBD0 U2236 ( .CLK(n2353), .C(n2354) );
  CKBD0 U2237 ( .CLK(n2354), .C(n2355) );
  CKBD0 U2238 ( .CLK(n2355), .C(n2356) );
  BUFFD0 U2239 ( .I(n2356), .Z(n2357) );
  CKBD0 U2240 ( .CLK(n2357), .C(n2358) );
  CKBD0 U2241 ( .CLK(n2358), .C(n2359) );
  CKBD0 U2242 ( .CLK(n2359), .C(n2360) );
  CKBD0 U2243 ( .CLK(n2360), .C(n2361) );
  CKBD0 U2244 ( .CLK(n2361), .C(n2362) );
  CKBD0 U2245 ( .CLK(n2362), .C(n2363) );
  CKBD0 U2246 ( .CLK(n2363), .C(n2364) );
  CKBD0 U2247 ( .CLK(n2364), .C(n2365) );
  CKBD0 U2248 ( .CLK(n2365), .C(n2366) );
  CKBD0 U2249 ( .CLK(n2366), .C(n2367) );
  BUFFD0 U2250 ( .I(n2367), .Z(n2368) );
  CKBD0 U2251 ( .CLK(n2368), .C(n2369) );
  CKBD0 U2252 ( .CLK(n2369), .C(n2370) );
  CKBD0 U2253 ( .CLK(n2370), .C(n2371) );
  CKBD0 U2254 ( .CLK(n2371), .C(n2372) );
  CKBD0 U2255 ( .CLK(n2372), .C(n2373) );
  CKBD0 U2256 ( .CLK(n2373), .C(n2374) );
  CKBD0 U2257 ( .CLK(n2374), .C(n2375) );
  CKBD0 U2258 ( .CLK(n2375), .C(n2376) );
  CKBD0 U2259 ( .CLK(n2376), .C(n2377) );
  CKBD0 U2260 ( .CLK(n2377), .C(n2378) );
  BUFFD0 U2261 ( .I(n2378), .Z(n2379) );
  CKBD0 U2262 ( .CLK(n2379), .C(n2380) );
  CKBD0 U2263 ( .CLK(n2380), .C(n2381) );
  CKBD0 U2264 ( .CLK(n2381), .C(n2382) );
  CKBD0 U2265 ( .CLK(n2382), .C(n2383) );
  CKBD0 U2266 ( .CLK(n2383), .C(n2384) );
  CKBD0 U2267 ( .CLK(n2384), .C(n2385) );
  CKBD0 U2268 ( .CLK(n2385), .C(n2386) );
  CKBD0 U2269 ( .CLK(n2386), .C(n2387) );
  CKBD0 U2270 ( .CLK(n2387), .C(n2388) );
  CKBD0 U2271 ( .CLK(n2388), .C(n2389) );
  BUFFD0 U2272 ( .I(n2389), .Z(n2390) );
  CKBD0 U2273 ( .CLK(n2390), .C(n2391) );
  CKBD0 U2274 ( .CLK(n2391), .C(n2392) );
  CKBD0 U2275 ( .CLK(n2392), .C(n2393) );
  CKBD0 U2276 ( .CLK(n2393), .C(n2394) );
  CKBD0 U2277 ( .CLK(n2394), .C(n2395) );
  CKBD0 U2278 ( .CLK(n2395), .C(n2396) );
  CKBD0 U2279 ( .CLK(n2396), .C(n2397) );
  CKBD0 U2280 ( .CLK(n2397), .C(n2398) );
  CKBD0 U2281 ( .CLK(n2398), .C(n2399) );
  CKBD0 U2282 ( .CLK(n2399), .C(n2400) );
  BUFFD0 U2283 ( .I(n2400), .Z(n2401) );
  CKBD0 U2284 ( .CLK(n2401), .C(n2402) );
  CKBD0 U2285 ( .CLK(n2402), .C(n2403) );
  CKBD0 U2286 ( .CLK(n2403), .C(n2404) );
  CKBD0 U2287 ( .CLK(n2404), .C(n2405) );
  BUFFD0 U2288 ( .I(n8234), .Z(n2406) );
  CKBD0 U2289 ( .CLK(FrameSR[51]), .C(n2407) );
  CKBD0 U2290 ( .CLK(n2407), .C(n2408) );
  CKBD0 U2291 ( .CLK(n2408), .C(n2409) );
  CKBD0 U2292 ( .CLK(n2409), .C(n2410) );
  CKBD0 U2293 ( .CLK(n2410), .C(n2411) );
  CKBD0 U2294 ( .CLK(n2411), .C(n2412) );
  CKBD0 U2295 ( .CLK(n2412), .C(n2413) );
  BUFFD0 U2296 ( .I(n2413), .Z(n2414) );
  CKBD0 U2297 ( .CLK(n2414), .C(n2415) );
  CKBD0 U2298 ( .CLK(n2415), .C(n2416) );
  CKBD0 U2299 ( .CLK(n2416), .C(n2417) );
  CKBD0 U2300 ( .CLK(n2417), .C(n2418) );
  CKBD0 U2301 ( .CLK(n2418), .C(n2419) );
  CKBD0 U2302 ( .CLK(n2419), .C(n2420) );
  CKBD0 U2303 ( .CLK(n2420), .C(n2421) );
  CKBD0 U2304 ( .CLK(n2421), .C(n2422) );
  CKBD0 U2305 ( .CLK(n2422), .C(n2423) );
  CKBD0 U2306 ( .CLK(n2423), .C(n2424) );
  BUFFD0 U2307 ( .I(n2424), .Z(n2425) );
  CKBD0 U2308 ( .CLK(n2425), .C(n2426) );
  CKBD0 U2309 ( .CLK(n2426), .C(n2427) );
  CKBD0 U2310 ( .CLK(n2427), .C(n2428) );
  CKBD0 U2311 ( .CLK(n2428), .C(n2429) );
  CKBD0 U2312 ( .CLK(n2429), .C(n2430) );
  CKBD0 U2313 ( .CLK(n2430), .C(n2431) );
  CKBD0 U2314 ( .CLK(n2431), .C(n2432) );
  CKBD0 U2315 ( .CLK(n2432), .C(n2433) );
  CKBD0 U2316 ( .CLK(n2433), .C(n2434) );
  CKBD0 U2317 ( .CLK(n2434), .C(n2435) );
  BUFFD0 U2318 ( .I(n2435), .Z(n2436) );
  CKBD0 U2319 ( .CLK(n2436), .C(n2437) );
  CKBD0 U2320 ( .CLK(n2437), .C(n2438) );
  CKBD0 U2321 ( .CLK(n2438), .C(n2439) );
  CKBD0 U2322 ( .CLK(n2439), .C(n2440) );
  CKBD0 U2323 ( .CLK(n2440), .C(n2441) );
  CKBD0 U2324 ( .CLK(n2441), .C(n2442) );
  CKBD0 U2325 ( .CLK(n2442), .C(n2443) );
  CKBD0 U2326 ( .CLK(n2443), .C(n2444) );
  CKBD0 U2327 ( .CLK(n2444), .C(n2445) );
  CKBD0 U2328 ( .CLK(n2445), .C(n2446) );
  BUFFD0 U2329 ( .I(n2446), .Z(n2447) );
  CKBD0 U2330 ( .CLK(n2447), .C(n2448) );
  CKBD0 U2331 ( .CLK(n2448), .C(n2449) );
  CKBD0 U2332 ( .CLK(n2449), .C(n2450) );
  CKBD0 U2333 ( .CLK(n2450), .C(n2451) );
  CKBD0 U2334 ( .CLK(n2451), .C(n2452) );
  CKBD0 U2335 ( .CLK(n2452), .C(n2453) );
  CKBD0 U2336 ( .CLK(n2453), .C(n2454) );
  CKBD0 U2337 ( .CLK(n2454), .C(n2455) );
  CKBD0 U2338 ( .CLK(n2455), .C(n2456) );
  BUFFD0 U2339 ( .I(n2456), .Z(n2457) );
  CKBD0 U2340 ( .CLK(n2457), .C(n2458) );
  CKBD0 U2341 ( .CLK(n2458), .C(n2459) );
  CKBD0 U2342 ( .CLK(n2459), .C(n2460) );
  CKBD0 U2343 ( .CLK(n2460), .C(n2461) );
  CKBD0 U2344 ( .CLK(n2461), .C(n2462) );
  CKBD0 U2345 ( .CLK(n2462), .C(n2463) );
  CKBD0 U2346 ( .CLK(n2463), .C(n2464) );
  CKBD0 U2347 ( .CLK(n2464), .C(n2465) );
  CKBD0 U2348 ( .CLK(n2465), .C(n2466) );
  CKBD0 U2349 ( .CLK(n2466), .C(n2467) );
  BUFFD0 U2350 ( .I(n2467), .Z(n2468) );
  CKBD0 U2351 ( .CLK(n2468), .C(n2469) );
  CKBD0 U2352 ( .CLK(n2469), .C(n2470) );
  CKBD0 U2353 ( .CLK(n2470), .C(n2471) );
  CKBD0 U2354 ( .CLK(n2471), .C(n2472) );
  CKBD0 U2355 ( .CLK(n2472), .C(n2473) );
  CKBD0 U2356 ( .CLK(n2473), .C(n2474) );
  CKBD0 U2357 ( .CLK(n2474), .C(n2475) );
  CKBD0 U2358 ( .CLK(n2475), .C(n2476) );
  CKBD0 U2359 ( .CLK(n2476), .C(n2477) );
  CKBD0 U2360 ( .CLK(n2477), .C(n2478) );
  BUFFD0 U2361 ( .I(n2478), .Z(n2479) );
  CKBD0 U2362 ( .CLK(n2479), .C(n2480) );
  CKBD0 U2363 ( .CLK(n2480), .C(n2481) );
  CKBD0 U2364 ( .CLK(n2481), .C(n2482) );
  CKBD0 U2365 ( .CLK(n2482), .C(n2483) );
  CKBD0 U2366 ( .CLK(n2483), .C(n2484) );
  CKBD0 U2367 ( .CLK(n2484), .C(n2485) );
  CKBD0 U2368 ( .CLK(n2485), .C(n2486) );
  CKBD0 U2369 ( .CLK(n2486), .C(n2487) );
  CKBD0 U2370 ( .CLK(n2487), .C(n2488) );
  CKBD0 U2371 ( .CLK(n2488), .C(n2489) );
  BUFFD0 U2372 ( .I(n2489), .Z(n2490) );
  CKBD0 U2373 ( .CLK(n2490), .C(n2491) );
  CKBD0 U2374 ( .CLK(n2491), .C(n2492) );
  CKBD0 U2375 ( .CLK(n2492), .C(n2493) );
  CKBD0 U2376 ( .CLK(n2493), .C(n2494) );
  CKBD0 U2377 ( .CLK(n2494), .C(n2495) );
  CKBD0 U2378 ( .CLK(n2495), .C(n2496) );
  CKBD0 U2379 ( .CLK(n2496), .C(n2497) );
  CKBD0 U2380 ( .CLK(n2497), .C(n2498) );
  CKBD0 U2381 ( .CLK(n2498), .C(n2499) );
  CKBD0 U2382 ( .CLK(n2499), .C(n2500) );
  BUFFD0 U2383 ( .I(n2500), .Z(n2501) );
  CKBD0 U2384 ( .CLK(n2501), .C(n2502) );
  CKBD0 U2385 ( .CLK(n2502), .C(n2503) );
  CKBD0 U2386 ( .CLK(n2503), .C(n2504) );
  BUFFD0 U2387 ( .I(n8223), .Z(n2505) );
  CKBD0 U2388 ( .CLK(FrameSR[16]), .C(n2506) );
  CKBD0 U2389 ( .CLK(n2506), .C(n2507) );
  CKBD0 U2390 ( .CLK(n2507), .C(n2508) );
  CKBD0 U2391 ( .CLK(n2508), .C(n2509) );
  CKBD0 U2392 ( .CLK(n2509), .C(n2510) );
  CKBD0 U2393 ( .CLK(n2510), .C(n2511) );
  CKBD0 U2394 ( .CLK(n2511), .C(n2512) );
  CKBD0 U2395 ( .CLK(n2512), .C(n2513) );
  CKBD0 U2396 ( .CLK(n2513), .C(n2514) );
  BUFFD0 U2397 ( .I(n2514), .Z(n2515) );
  CKBD0 U2398 ( .CLK(n2515), .C(n2516) );
  CKBD0 U2399 ( .CLK(n2516), .C(n2517) );
  CKBD0 U2400 ( .CLK(n2517), .C(n2518) );
  CKBD0 U2401 ( .CLK(n2518), .C(n2519) );
  CKBD0 U2402 ( .CLK(n2519), .C(n2520) );
  CKBD0 U2403 ( .CLK(n2520), .C(n2521) );
  CKBD0 U2404 ( .CLK(n2521), .C(n2522) );
  CKBD0 U2405 ( .CLK(n2522), .C(n2523) );
  CKBD0 U2406 ( .CLK(n2523), .C(n2524) );
  CKBD0 U2407 ( .CLK(n2524), .C(n2525) );
  BUFFD0 U2408 ( .I(n2525), .Z(n2526) );
  CKBD0 U2409 ( .CLK(n2526), .C(n2527) );
  CKBD0 U2410 ( .CLK(n2527), .C(n2528) );
  CKBD0 U2411 ( .CLK(n2528), .C(n2529) );
  CKBD0 U2412 ( .CLK(n2529), .C(n2530) );
  CKBD0 U2413 ( .CLK(n2530), .C(n2531) );
  CKBD0 U2414 ( .CLK(n2531), .C(n2532) );
  CKBD0 U2415 ( .CLK(n2532), .C(n2533) );
  CKBD0 U2416 ( .CLK(n2533), .C(n2534) );
  CKBD0 U2417 ( .CLK(n2534), .C(n2535) );
  CKBD0 U2418 ( .CLK(n2535), .C(n2536) );
  BUFFD0 U2419 ( .I(n2536), .Z(n2537) );
  CKBD0 U2420 ( .CLK(n2537), .C(n2538) );
  CKBD0 U2421 ( .CLK(n2538), .C(n2539) );
  CKBD0 U2422 ( .CLK(n2539), .C(n2540) );
  CKBD0 U2423 ( .CLK(n2540), .C(n2541) );
  CKBD0 U2424 ( .CLK(n2541), .C(n2542) );
  CKBD0 U2425 ( .CLK(n2542), .C(n2543) );
  CKBD0 U2426 ( .CLK(n2543), .C(n2544) );
  CKBD0 U2427 ( .CLK(n2544), .C(n2545) );
  CKBD0 U2428 ( .CLK(n2545), .C(n2546) );
  CKBD0 U2429 ( .CLK(n2546), .C(n2547) );
  BUFFD0 U2430 ( .I(n2547), .Z(n2548) );
  CKBD0 U2431 ( .CLK(n2548), .C(n2549) );
  CKBD0 U2432 ( .CLK(n2549), .C(n2550) );
  CKBD0 U2433 ( .CLK(n2550), .C(n2551) );
  CKBD0 U2434 ( .CLK(n2551), .C(n2552) );
  CKBD0 U2435 ( .CLK(n2552), .C(n2553) );
  CKBD0 U2436 ( .CLK(n2553), .C(n2554) );
  CKBD0 U2437 ( .CLK(n2554), .C(n2555) );
  CKBD0 U2438 ( .CLK(n2555), .C(n2556) );
  CKBD0 U2439 ( .CLK(n2556), .C(n2557) );
  CKBD0 U2440 ( .CLK(n2557), .C(n2558) );
  BUFFD0 U2441 ( .I(n2558), .Z(n2559) );
  CKBD0 U2442 ( .CLK(n2559), .C(n2560) );
  CKBD0 U2443 ( .CLK(n2560), .C(n2561) );
  CKBD0 U2444 ( .CLK(n2561), .C(n2562) );
  CKBD0 U2445 ( .CLK(n2562), .C(n2563) );
  CKBD0 U2446 ( .CLK(n2563), .C(n2564) );
  CKBD0 U2447 ( .CLK(n2564), .C(n2565) );
  CKBD0 U2448 ( .CLK(n2565), .C(n2566) );
  CKBD0 U2449 ( .CLK(n2566), .C(n2567) );
  CKBD0 U2450 ( .CLK(n2567), .C(n2568) );
  CKBD0 U2451 ( .CLK(n2568), .C(n2569) );
  BUFFD0 U2452 ( .I(n2569), .Z(n2570) );
  CKBD0 U2453 ( .CLK(n2570), .C(n2571) );
  CKBD0 U2454 ( .CLK(n2571), .C(n2572) );
  CKBD0 U2455 ( .CLK(n2572), .C(n2573) );
  CKBD0 U2456 ( .CLK(n2573), .C(n2574) );
  CKBD0 U2457 ( .CLK(n2574), .C(n2575) );
  CKBD0 U2458 ( .CLK(n2575), .C(n2576) );
  CKBD0 U2459 ( .CLK(n2576), .C(n2577) );
  CKBD0 U2460 ( .CLK(n2577), .C(n2578) );
  CKBD0 U2461 ( .CLK(n2578), .C(n2579) );
  BUFFD0 U2462 ( .I(n2579), .Z(n2580) );
  CKBD0 U2463 ( .CLK(n2580), .C(n2581) );
  CKBD0 U2464 ( .CLK(n2581), .C(n2582) );
  CKBD0 U2465 ( .CLK(n2582), .C(n2583) );
  CKBD0 U2466 ( .CLK(n2583), .C(n2584) );
  CKBD0 U2467 ( .CLK(n2584), .C(n2585) );
  CKBD0 U2468 ( .CLK(n2585), .C(n2586) );
  CKBD0 U2469 ( .CLK(n2586), .C(n2587) );
  CKBD0 U2470 ( .CLK(n2587), .C(n2588) );
  CKBD0 U2471 ( .CLK(n2588), .C(n2589) );
  CKBD0 U2472 ( .CLK(n2589), .C(n2590) );
  BUFFD0 U2473 ( .I(n2590), .Z(n2591) );
  CKBD0 U2474 ( .CLK(n2591), .C(n2592) );
  CKBD0 U2475 ( .CLK(n2592), .C(n2593) );
  CKBD0 U2476 ( .CLK(n2593), .C(n2594) );
  CKBD0 U2477 ( .CLK(n2594), .C(n2595) );
  CKBD0 U2478 ( .CLK(n2595), .C(n2596) );
  CKBD0 U2479 ( .CLK(n2596), .C(n2597) );
  CKBD0 U2480 ( .CLK(n2597), .C(n2598) );
  CKBD0 U2481 ( .CLK(n2598), .C(n2599) );
  CKBD0 U2482 ( .CLK(n2599), .C(n2600) );
  CKBD0 U2483 ( .CLK(n2600), .C(n2601) );
  CKBD0 U2484 ( .CLK(n2601), .C(n2602) );
  CKBD0 U2485 ( .CLK(n2602), .C(n2603) );
  BUFFD0 U2486 ( .I(n6006), .Z(n2604) );
  CKBD0 U2487 ( .CLK(FrameSR[15]), .C(n2605) );
  BUFFD0 U2488 ( .I(N42), .Z(n2606) );
  BUFFD0 U2489 ( .I(n2738), .Z(n2607) );
  CKBD0 U2490 ( .CLK(FrameSR[63]), .C(n2608) );
  CKBD0 U2491 ( .CLK(n2608), .C(n2609) );
  CKBD0 U2492 ( .CLK(n2609), .C(n2610) );
  CKBD0 U2493 ( .CLK(n2610), .C(n2611) );
  CKBD0 U2494 ( .CLK(n2611), .C(n2612) );
  CKBD0 U2495 ( .CLK(n2612), .C(n2613) );
  CKBD0 U2496 ( .CLK(n2613), .C(n2614) );
  CKBD0 U2497 ( .CLK(n2614), .C(n2615) );
  CKBD0 U2498 ( .CLK(n2615), .C(n2616) );
  CKBD0 U2499 ( .CLK(n2616), .C(n2617) );
  BUFFD0 U2500 ( .I(n2617), .Z(n2618) );
  CKBD0 U2501 ( .CLK(n2618), .C(n2619) );
  CKBD0 U2502 ( .CLK(n2619), .C(n2620) );
  CKBD0 U2503 ( .CLK(n2620), .C(n2621) );
  CKBD0 U2504 ( .CLK(n2621), .C(n2622) );
  CKBD0 U2505 ( .CLK(n2622), .C(n2623) );
  CKBD0 U2506 ( .CLK(n2623), .C(n2624) );
  CKBD0 U2507 ( .CLK(n2624), .C(n2625) );
  CKBD0 U2508 ( .CLK(n2625), .C(n2626) );
  CKBD0 U2509 ( .CLK(n2626), .C(n2627) );
  CKBD0 U2510 ( .CLK(n2627), .C(n2628) );
  BUFFD0 U2511 ( .I(n2628), .Z(n2629) );
  CKBD0 U2512 ( .CLK(n2629), .C(n2630) );
  CKBD0 U2513 ( .CLK(n2630), .C(n2631) );
  CKBD0 U2514 ( .CLK(n2631), .C(n2632) );
  CKBD0 U2515 ( .CLK(n2632), .C(n2633) );
  CKBD0 U2516 ( .CLK(n2633), .C(n2634) );
  CKBD0 U2517 ( .CLK(n2634), .C(n2635) );
  CKBD0 U2518 ( .CLK(n2635), .C(n2636) );
  CKBD0 U2519 ( .CLK(n2636), .C(n2637) );
  CKBD0 U2520 ( .CLK(n2637), .C(n2638) );
  CKBD0 U2521 ( .CLK(n2638), .C(n2639) );
  BUFFD0 U2522 ( .I(n2639), .Z(n2640) );
  CKBD0 U2523 ( .CLK(n2640), .C(n2641) );
  CKBD0 U2524 ( .CLK(n2641), .C(n2642) );
  CKBD0 U2525 ( .CLK(n2642), .C(n2643) );
  CKBD0 U2526 ( .CLK(n2643), .C(n2644) );
  CKBD0 U2527 ( .CLK(n2644), .C(n2645) );
  CKBD0 U2528 ( .CLK(n2645), .C(n2646) );
  CKBD0 U2529 ( .CLK(n2646), .C(n2647) );
  CKBD0 U2530 ( .CLK(n2647), .C(n2648) );
  CKBD0 U2531 ( .CLK(n2648), .C(n2649) );
  CKBD0 U2532 ( .CLK(n2649), .C(n2650) );
  BUFFD0 U2533 ( .I(n2650), .Z(n2651) );
  CKBD0 U2534 ( .CLK(n2651), .C(n2652) );
  CKBD0 U2535 ( .CLK(n2652), .C(n2653) );
  CKBD0 U2536 ( .CLK(n2653), .C(n2654) );
  CKBD0 U2537 ( .CLK(n2654), .C(n2655) );
  CKBD0 U2538 ( .CLK(n2655), .C(n2656) );
  CKBD0 U2539 ( .CLK(n2656), .C(n2657) );
  CKBD0 U2540 ( .CLK(n2657), .C(n2658) );
  CKBD0 U2541 ( .CLK(n2658), .C(n2659) );
  CKBD0 U2542 ( .CLK(n2659), .C(n2660) );
  CKBD0 U2543 ( .CLK(n2660), .C(n2661) );
  BUFFD0 U2544 ( .I(n2661), .Z(n2662) );
  CKBD0 U2545 ( .CLK(n2662), .C(n2663) );
  CKBD0 U2546 ( .CLK(n2663), .C(n2664) );
  CKBD0 U2547 ( .CLK(n2664), .C(n2665) );
  CKBD0 U2548 ( .CLK(n2665), .C(n2666) );
  CKBD0 U2549 ( .CLK(n2666), .C(n2667) );
  CKBD0 U2550 ( .CLK(n2667), .C(n2668) );
  CKBD0 U2551 ( .CLK(n2668), .C(n2669) );
  CKBD0 U2552 ( .CLK(n2669), .C(n2670) );
  CKBD0 U2553 ( .CLK(n2670), .C(n2671) );
  CKBD0 U2554 ( .CLK(n2671), .C(n2672) );
  BUFFD0 U2555 ( .I(n2672), .Z(n2673) );
  CKBD0 U2556 ( .CLK(n2673), .C(n2674) );
  CKBD0 U2557 ( .CLK(n2674), .C(n2675) );
  CKBD0 U2558 ( .CLK(n2675), .C(n2676) );
  CKBD0 U2559 ( .CLK(n2676), .C(n2677) );
  CKBD0 U2560 ( .CLK(n2677), .C(n2678) );
  CKBD0 U2561 ( .CLK(n2678), .C(n2679) );
  CKBD0 U2562 ( .CLK(n2679), .C(n2680) );
  CKBD0 U2563 ( .CLK(n2680), .C(n2681) );
  CKBD0 U2564 ( .CLK(n2681), .C(n2682) );
  BUFFD0 U2565 ( .I(n2682), .Z(n2683) );
  CKBD0 U2566 ( .CLK(n2683), .C(n2684) );
  CKBD0 U2567 ( .CLK(n2684), .C(n2685) );
  CKBD0 U2568 ( .CLK(n2685), .C(n2686) );
  CKBD0 U2569 ( .CLK(n2686), .C(n2687) );
  CKBD0 U2570 ( .CLK(n2687), .C(n2688) );
  CKBD0 U2571 ( .CLK(n2688), .C(n2689) );
  CKBD0 U2572 ( .CLK(n2689), .C(n2690) );
  CKBD0 U2573 ( .CLK(n2690), .C(n2691) );
  CKBD0 U2574 ( .CLK(n2691), .C(n2692) );
  CKBD0 U2575 ( .CLK(n2692), .C(n2693) );
  BUFFD0 U2576 ( .I(n2693), .Z(n2694) );
  CKBD0 U2577 ( .CLK(n2694), .C(n2695) );
  CKBD0 U2578 ( .CLK(n2695), .C(n2696) );
  CKBD0 U2579 ( .CLK(n2696), .C(n2697) );
  CKBD0 U2580 ( .CLK(n2697), .C(n2698) );
  CKBD0 U2581 ( .CLK(n2698), .C(n2699) );
  CKBD0 U2582 ( .CLK(n2699), .C(n2700) );
  CKBD0 U2583 ( .CLK(n2700), .C(n2701) );
  CKBD0 U2584 ( .CLK(n2701), .C(n2702) );
  CKBD0 U2585 ( .CLK(n2702), .C(n2703) );
  CKBD0 U2586 ( .CLK(n2703), .C(n2704) );
  BUFFD0 U2587 ( .I(n2704), .Z(n2705) );
  CKBD0 U2588 ( .CLK(n2705), .C(n2706) );
  CKBD0 U2589 ( .CLK(n2706), .C(n2707) );
  CKBD0 U2590 ( .CLK(n2707), .C(n2708) );
  CKBD0 U2591 ( .CLK(n2708), .C(n2709) );
  BUFFD0 U2592 ( .I(n2709), .Z(n2710) );
  CKBD0 U2593 ( .CLK(n2710), .C(n2711) );
  BUFFD0 U2594 ( .I(n2711), .Z(n2712) );
  CKBD0 U2595 ( .CLK(n2712), .C(n2713) );
  BUFFD0 U2596 ( .I(n2713), .Z(n2714) );
  CKBD0 U2597 ( .CLK(n2714), .C(n2715) );
  BUFFD0 U2598 ( .I(n2715), .Z(n2716) );
  CKBD0 U2599 ( .CLK(n2716), .C(n2717) );
  BUFFD0 U2600 ( .I(n2717), .Z(n2718) );
  CKBD0 U2601 ( .CLK(n2718), .C(n2719) );
  BUFFD0 U2602 ( .I(n2719), .Z(n2720) );
  CKBD0 U2603 ( .CLK(n2720), .C(n2721) );
  BUFFD0 U2604 ( .I(n2721), .Z(n2722) );
  CKBD0 U2605 ( .CLK(n2722), .C(n2723) );
  BUFFD0 U2606 ( .I(n2723), .Z(n2724) );
  CKBD0 U2607 ( .CLK(n2724), .C(n2725) );
  BUFFD0 U2608 ( .I(n2725), .Z(n2726) );
  CKBD0 U2609 ( .CLK(n2726), .C(n2727) );
  BUFFD0 U2610 ( .I(n2727), .Z(n2728) );
  CKBD0 U2611 ( .CLK(n2728), .C(n2729) );
  BUFFD0 U2612 ( .I(n2729), .Z(n2730) );
  CKBD0 U2613 ( .CLK(n2730), .C(n2731) );
  BUFFD0 U2614 ( .I(n2731), .Z(n2732) );
  CKBD0 U2615 ( .CLK(n2732), .C(n2733) );
  BUFFD0 U2616 ( .I(n2733), .Z(n2734) );
  CKBD0 U2617 ( .CLK(n2734), .C(n2735) );
  BUFFD0 U2618 ( .I(n2735), .Z(n2736) );
  CKBD0 U2619 ( .CLK(n2736), .C(n2737) );
  BUFFD0 U2620 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2621 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2622 ( .I(n9168), .Z(n2740) );
  BUFFD0 U2623 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2624 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2625 ( .I(n9169), .Z(n2743) );
  CKBD0 U2626 ( .CLK(n5), .C(n2744) );
  CKBD0 U2627 ( .CLK(n2744), .C(n2745) );
  CKBD0 U2628 ( .CLK(n2745), .C(n2746) );
  BUFFD0 U2629 ( .I(n2746), .Z(n2747) );
  CKBD0 U2630 ( .CLK(n2747), .C(n2748) );
  CKBD0 U2631 ( .CLK(n2748), .C(n2749) );
  CKBD0 U2632 ( .CLK(n2749), .C(n2750) );
  CKBD0 U2633 ( .CLK(n2750), .C(n2751) );
  CKBD0 U2634 ( .CLK(n2751), .C(n2752) );
  CKBD0 U2635 ( .CLK(n2752), .C(n2753) );
  CKBD0 U2636 ( .CLK(n2753), .C(n2754) );
  CKBD0 U2637 ( .CLK(n2754), .C(n2755) );
  CKBD0 U2638 ( .CLK(n2755), .C(n2756) );
  CKBD0 U2639 ( .CLK(n2756), .C(n2757) );
  BUFFD0 U2640 ( .I(n2757), .Z(n2758) );
  CKBD0 U2641 ( .CLK(n2758), .C(n2759) );
  CKBD0 U2642 ( .CLK(n2759), .C(n2760) );
  CKBD0 U2643 ( .CLK(n2760), .C(n2761) );
  CKBD0 U2644 ( .CLK(n2761), .C(n2762) );
  CKBD0 U2645 ( .CLK(n2762), .C(n2763) );
  CKBD0 U2646 ( .CLK(n2763), .C(n2764) );
  CKBD0 U2647 ( .CLK(n2764), .C(n2765) );
  CKBD0 U2648 ( .CLK(n2765), .C(n2766) );
  CKBD0 U2649 ( .CLK(n2766), .C(n2767) );
  CKBD0 U2650 ( .CLK(n2767), .C(n2768) );
  BUFFD0 U2651 ( .I(n2768), .Z(n2769) );
  CKBD0 U2652 ( .CLK(n2769), .C(n2770) );
  CKBD0 U2653 ( .CLK(n2770), .C(n2771) );
  CKBD0 U2654 ( .CLK(n2771), .C(n2772) );
  CKBD0 U2655 ( .CLK(n2772), .C(n2773) );
  CKBD0 U2656 ( .CLK(n2773), .C(n2774) );
  CKBD0 U2657 ( .CLK(n2774), .C(n2775) );
  CKBD0 U2658 ( .CLK(n2775), .C(n2776) );
  CKBD0 U2659 ( .CLK(n2776), .C(n2777) );
  CKBD0 U2660 ( .CLK(n2777), .C(n2778) );
  CKBD0 U2661 ( .CLK(n2778), .C(n2779) );
  BUFFD0 U2662 ( .I(n2779), .Z(n2780) );
  CKBD0 U2663 ( .CLK(n2780), .C(n2781) );
  CKBD0 U2664 ( .CLK(n2781), .C(n2782) );
  CKBD0 U2665 ( .CLK(n2782), .C(n2783) );
  CKBD0 U2666 ( .CLK(n2783), .C(n2784) );
  CKBD0 U2667 ( .CLK(n2784), .C(n2785) );
  CKBD0 U2668 ( .CLK(n2785), .C(n2786) );
  CKBD0 U2669 ( .CLK(n2786), .C(n2787) );
  CKBD0 U2670 ( .CLK(n2787), .C(n2788) );
  CKBD0 U2671 ( .CLK(n2788), .C(n2789) );
  BUFFD0 U2672 ( .I(n2789), .Z(n2790) );
  CKBD0 U2673 ( .CLK(n2790), .C(n2791) );
  CKBD0 U2674 ( .CLK(n2791), .C(n2792) );
  CKBD0 U2675 ( .CLK(n2792), .C(n2793) );
  CKBD0 U2676 ( .CLK(n2793), .C(n2794) );
  CKBD0 U2677 ( .CLK(n2794), .C(n2795) );
  CKBD0 U2678 ( .CLK(n2795), .C(n2796) );
  CKBD0 U2679 ( .CLK(n2796), .C(n2797) );
  CKBD0 U2680 ( .CLK(n2797), .C(n2798) );
  CKBD0 U2681 ( .CLK(n2798), .C(n2799) );
  CKBD0 U2682 ( .CLK(n2799), .C(n2800) );
  CKBD0 U2683 ( .CLK(n2800), .C(n2801) );
  BUFFD0 U2684 ( .I(n2801), .Z(n2802) );
  CKBD0 U2685 ( .CLK(n2802), .C(n2803) );
  CKBD0 U2686 ( .CLK(n2803), .C(n2804) );
  CKBD0 U2687 ( .CLK(n2804), .C(n2805) );
  CKBD0 U2688 ( .CLK(n2805), .C(n2806) );
  CKBD0 U2689 ( .CLK(n2806), .C(n2807) );
  CKBD0 U2690 ( .CLK(n2807), .C(n2808) );
  CKBD0 U2691 ( .CLK(n2808), .C(n2809) );
  CKBD0 U2692 ( .CLK(n2809), .C(n2810) );
  CKBD0 U2693 ( .CLK(n2810), .C(n2811) );
  BUFFD0 U2694 ( .I(n2811), .Z(n2812) );
  CKBD0 U2695 ( .CLK(n2812), .C(n2813) );
  CKBD0 U2696 ( .CLK(n2813), .C(n2814) );
  CKBD0 U2697 ( .CLK(n2814), .C(n2815) );
  CKBD0 U2698 ( .CLK(n2815), .C(n2816) );
  CKBD0 U2699 ( .CLK(n2816), .C(n2817) );
  CKBD0 U2700 ( .CLK(n2817), .C(n2818) );
  CKBD0 U2701 ( .CLK(n2818), .C(n2819) );
  CKBD0 U2702 ( .CLK(n2819), .C(n2820) );
  CKBD0 U2703 ( .CLK(n2820), .C(n2821) );
  CKBD0 U2704 ( .CLK(n2821), .C(n2822) );
  BUFFD0 U2705 ( .I(n2822), .Z(n2823) );
  CKBD0 U2706 ( .CLK(n2823), .C(n2824) );
  CKBD0 U2707 ( .CLK(n2824), .C(n2825) );
  CKBD0 U2708 ( .CLK(n2825), .C(n2826) );
  CKBD0 U2709 ( .CLK(n2826), .C(n2827) );
  CKBD0 U2710 ( .CLK(n2827), .C(n2828) );
  CKBD0 U2711 ( .CLK(n2828), .C(n2829) );
  CKBD0 U2712 ( .CLK(n2829), .C(n2830) );
  CKBD0 U2713 ( .CLK(n2830), .C(n2831) );
  CKBD0 U2714 ( .CLK(n2831), .C(n2832) );
  CKBD0 U2715 ( .CLK(n2832), .C(n2833) );
  BUFFD0 U2716 ( .I(n2833), .Z(n2834) );
  CKBD0 U2717 ( .CLK(n2834), .C(n2835) );
  CKBD0 U2718 ( .CLK(n2835), .C(n2836) );
  CKBD0 U2719 ( .CLK(n2836), .C(n2837) );
  CKBD0 U2720 ( .CLK(n2837), .C(n2838) );
  CKBD0 U2721 ( .CLK(n2838), .C(n2839) );
  CKBD0 U2722 ( .CLK(n2839), .C(n2840) );
  CKBD0 U2723 ( .CLK(n2840), .C(n2841) );
  CKBD0 U2724 ( .CLK(n2841), .C(n2842) );
  CKBD0 U2725 ( .CLK(n2842), .C(n2843) );
  CKBD0 U2726 ( .CLK(n2843), .C(n2844) );
  BUFFD0 U2727 ( .I(n2844), .Z(n2845) );
  CKBD0 U2728 ( .CLK(n2845), .C(n2846) );
  CKBD0 U2729 ( .CLK(n2846), .C(n2847) );
  CKBD0 U2730 ( .CLK(n2847), .C(n2848) );
  CKBD0 U2731 ( .CLK(n2848), .C(n2849) );
  CKBD0 U2732 ( .CLK(n2849), .C(n2850) );
  CKBD0 U2733 ( .CLK(n2850), .C(n2851) );
  CKBD0 U2734 ( .CLK(n2851), .C(n2852) );
  CKBD0 U2735 ( .CLK(n2852), .C(n2853) );
  CKBD0 U2736 ( .CLK(n2853), .C(n2854) );
  BUFFD0 U2737 ( .I(n2854), .Z(n2855) );
  CKBD0 U2738 ( .CLK(n2855), .C(n2856) );
  CKBD0 U2739 ( .CLK(n2856), .C(n2857) );
  CKBD0 U2740 ( .CLK(n2857), .C(n2858) );
  CKBD0 U2741 ( .CLK(n2858), .C(n2859) );
  CKBD0 U2742 ( .CLK(n2859), .C(n2860) );
  CKBD0 U2743 ( .CLK(n2860), .C(n2861) );
  BUFFD0 U2744 ( .I(n2861), .Z(n2862) );
  CKBD0 U2745 ( .CLK(n2862), .C(n2863) );
  BUFFD0 U2746 ( .I(n2863), .Z(n2864) );
  CKBD0 U2747 ( .CLK(n2864), .C(n2865) );
  BUFFD0 U2748 ( .I(n2865), .Z(n2866) );
  CKBD0 U2749 ( .CLK(n2866), .C(n2867) );
  BUFFD0 U2750 ( .I(n2867), .Z(n2868) );
  CKBD0 U2751 ( .CLK(n2868), .C(n2869) );
  BUFFD0 U2752 ( .I(n2869), .Z(n2870) );
  CKBD0 U2753 ( .CLK(n2870), .C(n2871) );
  BUFFD0 U2754 ( .I(n2871), .Z(n2872) );
  CKBD0 U2755 ( .CLK(n2872), .C(n2873) );
  BUFFD0 U2756 ( .I(n2873), .Z(n2874) );
  CKBD0 U2757 ( .CLK(n2874), .C(n2875) );
  BUFFD0 U2758 ( .I(n2875), .Z(n2876) );
  BUFFD0 U2759 ( .I(n2878), .Z(n2877) );
  BUFFD0 U2760 ( .I(n2879), .Z(n2878) );
  BUFFD0 U2761 ( .I(n9170), .Z(n2879) );
  CKBD0 U2762 ( .CLK(n1389), .C(n2880) );
  CKBD0 U2763 ( .CLK(n2880), .C(n2881) );
  CKBD0 U2764 ( .CLK(n2881), .C(n2882) );
  BUFFD0 U2765 ( .I(n2882), .Z(n2883) );
  CKBD0 U2766 ( .CLK(n2883), .C(n2884) );
  CKBD0 U2767 ( .CLK(n2884), .C(n2885) );
  CKBD0 U2768 ( .CLK(n2885), .C(n2886) );
  CKBD0 U2769 ( .CLK(n2886), .C(n2887) );
  CKBD0 U2770 ( .CLK(n2887), .C(n2888) );
  CKBD0 U2771 ( .CLK(n2888), .C(n2889) );
  CKBD0 U2772 ( .CLK(n2889), .C(n2890) );
  CKBD0 U2773 ( .CLK(n2890), .C(n2891) );
  CKBD0 U2774 ( .CLK(n2891), .C(n2892) );
  CKBD0 U2775 ( .CLK(n2892), .C(n2893) );
  BUFFD0 U2776 ( .I(n2893), .Z(n2894) );
  CKBD0 U2777 ( .CLK(n2894), .C(n2895) );
  CKBD0 U2778 ( .CLK(n2895), .C(n2896) );
  CKBD0 U2779 ( .CLK(n2896), .C(n2897) );
  CKBD0 U2780 ( .CLK(n2897), .C(n2898) );
  CKBD0 U2781 ( .CLK(n2898), .C(n2899) );
  CKBD0 U2782 ( .CLK(n2899), .C(n2900) );
  CKBD0 U2783 ( .CLK(n2900), .C(n2901) );
  CKBD0 U2784 ( .CLK(n2901), .C(n2902) );
  CKBD0 U2785 ( .CLK(n2902), .C(n2903) );
  CKBD0 U2786 ( .CLK(n2903), .C(n2904) );
  BUFFD0 U2787 ( .I(n2904), .Z(n2905) );
  CKBD0 U2788 ( .CLK(n2905), .C(n2906) );
  CKBD0 U2789 ( .CLK(n2906), .C(n2907) );
  CKBD0 U2790 ( .CLK(n2907), .C(n2908) );
  CKBD0 U2791 ( .CLK(n2908), .C(n2909) );
  CKBD0 U2792 ( .CLK(n2909), .C(n2910) );
  CKBD0 U2793 ( .CLK(n2910), .C(n2911) );
  CKBD0 U2794 ( .CLK(n2911), .C(n2912) );
  CKBD0 U2795 ( .CLK(n2912), .C(n2913) );
  CKBD0 U2796 ( .CLK(n2913), .C(n2914) );
  CKBD0 U2797 ( .CLK(n2914), .C(n2915) );
  BUFFD0 U2798 ( .I(n2915), .Z(n2916) );
  CKBD0 U2799 ( .CLK(n2916), .C(n2917) );
  CKBD0 U2800 ( .CLK(n2917), .C(n2918) );
  CKBD0 U2801 ( .CLK(n2918), .C(n2919) );
  CKBD0 U2802 ( .CLK(n2919), .C(n2920) );
  CKBD0 U2803 ( .CLK(n2920), .C(n2921) );
  CKBD0 U2804 ( .CLK(n2921), .C(n2922) );
  CKBD0 U2805 ( .CLK(n2922), .C(n2923) );
  CKBD0 U2806 ( .CLK(n2923), .C(n2924) );
  CKBD0 U2807 ( .CLK(n2924), .C(n2925) );
  BUFFD0 U2808 ( .I(n2925), .Z(n2926) );
  CKBD0 U2809 ( .CLK(n2926), .C(n2927) );
  CKBD0 U2810 ( .CLK(n2927), .C(n2928) );
  CKBD0 U2811 ( .CLK(n2928), .C(n2929) );
  CKBD0 U2812 ( .CLK(n2929), .C(n2930) );
  CKBD0 U2813 ( .CLK(n2930), .C(n2931) );
  CKBD0 U2814 ( .CLK(n2931), .C(n2932) );
  CKBD0 U2815 ( .CLK(n2932), .C(n2933) );
  CKBD0 U2816 ( .CLK(n2933), .C(n2934) );
  CKBD0 U2817 ( .CLK(n2934), .C(n2935) );
  CKBD0 U2818 ( .CLK(n2935), .C(n2936) );
  CKBD0 U2819 ( .CLK(n2936), .C(n2937) );
  BUFFD0 U2820 ( .I(n2937), .Z(n2938) );
  CKBD0 U2821 ( .CLK(n2938), .C(n2939) );
  CKBD0 U2822 ( .CLK(n2939), .C(n2940) );
  CKBD0 U2823 ( .CLK(n2940), .C(n2941) );
  CKBD0 U2824 ( .CLK(n2941), .C(n2942) );
  CKBD0 U2825 ( .CLK(n2942), .C(n2943) );
  CKBD0 U2826 ( .CLK(n2943), .C(n2944) );
  CKBD0 U2827 ( .CLK(n2944), .C(n2945) );
  CKBD0 U2828 ( .CLK(n2945), .C(n2946) );
  CKBD0 U2829 ( .CLK(n2946), .C(n2947) );
  BUFFD0 U2830 ( .I(n2947), .Z(n2948) );
  CKBD0 U2831 ( .CLK(n2948), .C(n2949) );
  CKBD0 U2832 ( .CLK(n2949), .C(n2950) );
  CKBD0 U2833 ( .CLK(n2950), .C(n2951) );
  CKBD0 U2834 ( .CLK(n2951), .C(n2952) );
  CKBD0 U2835 ( .CLK(n2952), .C(n2953) );
  CKBD0 U2836 ( .CLK(n2953), .C(n2954) );
  CKBD0 U2837 ( .CLK(n2954), .C(n2955) );
  CKBD0 U2838 ( .CLK(n2955), .C(n2956) );
  CKBD0 U2839 ( .CLK(n2956), .C(n2957) );
  CKBD0 U2840 ( .CLK(n2957), .C(n2958) );
  BUFFD0 U2841 ( .I(n2958), .Z(n2959) );
  CKBD0 U2842 ( .CLK(n2959), .C(n2960) );
  CKBD0 U2843 ( .CLK(n2960), .C(n2961) );
  CKBD0 U2844 ( .CLK(n2961), .C(n2962) );
  CKBD0 U2845 ( .CLK(n2962), .C(n2963) );
  CKBD0 U2846 ( .CLK(n2963), .C(n2964) );
  CKBD0 U2847 ( .CLK(n2964), .C(n2965) );
  CKBD0 U2848 ( .CLK(n2965), .C(n2966) );
  CKBD0 U2849 ( .CLK(n2966), .C(n2967) );
  CKBD0 U2850 ( .CLK(n2967), .C(n2968) );
  CKBD0 U2851 ( .CLK(n2968), .C(n2969) );
  BUFFD0 U2852 ( .I(n2969), .Z(n2970) );
  CKBD0 U2853 ( .CLK(n2970), .C(n2971) );
  CKBD0 U2854 ( .CLK(n2971), .C(n2972) );
  CKBD0 U2855 ( .CLK(n2972), .C(n2973) );
  CKBD0 U2856 ( .CLK(n2973), .C(n2974) );
  CKBD0 U2857 ( .CLK(n2974), .C(n2975) );
  CKBD0 U2858 ( .CLK(n2975), .C(n2976) );
  CKBD0 U2859 ( .CLK(n2976), .C(n2977) );
  CKBD0 U2860 ( .CLK(n2977), .C(n2978) );
  CKBD0 U2861 ( .CLK(n2978), .C(n2979) );
  CKBD0 U2862 ( .CLK(n2979), .C(n2980) );
  BUFFD0 U2863 ( .I(n2980), .Z(n2981) );
  CKBD0 U2864 ( .CLK(n2981), .C(n2982) );
  CKBD0 U2865 ( .CLK(n2982), .C(n2983) );
  CKBD0 U2866 ( .CLK(n2983), .C(n2984) );
  CKBD0 U2867 ( .CLK(n2984), .C(n2985) );
  CKBD0 U2868 ( .CLK(n2985), .C(n2986) );
  CKBD0 U2869 ( .CLK(n2986), .C(n2987) );
  CKBD0 U2870 ( .CLK(n2987), .C(n2988) );
  CKBD0 U2871 ( .CLK(n2988), .C(n2989) );
  CKBD0 U2872 ( .CLK(n2989), .C(n2990) );
  CKBD0 U2873 ( .CLK(n2990), .C(n2991) );
  BUFFD0 U2874 ( .I(n2991), .Z(n2992) );
  CKBD0 U2875 ( .CLK(n2992), .C(n2993) );
  CKBD0 U2876 ( .CLK(n2993), .C(n2994) );
  CKBD0 U2877 ( .CLK(n2994), .C(n2995) );
  CKBD0 U2878 ( .CLK(n2995), .C(n2996) );
  CKBD0 U2879 ( .CLK(n2996), .C(n2997) );
  BUFFD0 U2880 ( .I(n2997), .Z(n2998) );
  CKBD0 U2881 ( .CLK(n2998), .C(n2999) );
  BUFFD0 U2882 ( .I(n2999), .Z(n3000) );
  CKBD0 U2883 ( .CLK(n3000), .C(n3001) );
  BUFFD0 U2884 ( .I(n3001), .Z(n3002) );
  CKBD0 U2885 ( .CLK(n3002), .C(n3003) );
  BUFFD0 U2886 ( .I(n3003), .Z(n3004) );
  CKBD0 U2887 ( .CLK(n3004), .C(n3005) );
  BUFFD0 U2888 ( .I(n3005), .Z(n3006) );
  CKBD0 U2889 ( .CLK(n3006), .C(n3007) );
  BUFFD0 U2890 ( .I(n3007), .Z(n3008) );
  CKBD0 U2891 ( .CLK(n3008), .C(n3009) );
  BUFFD0 U2892 ( .I(n3009), .Z(n3010) );
  CKBD0 U2893 ( .CLK(n3010), .C(n3011) );
  BUFFD0 U2894 ( .I(n3011), .Z(n3012) );
  BUFFD0 U2895 ( .I(n3014), .Z(n3013) );
  BUFFD0 U2896 ( .I(n3015), .Z(n3014) );
  BUFFD0 U2897 ( .I(n9171), .Z(n3015) );
  CKBD0 U2898 ( .CLK(n1387), .C(n3016) );
  CKBD0 U2899 ( .CLK(n3016), .C(n3017) );
  CKBD0 U2900 ( .CLK(n3017), .C(n3018) );
  BUFFD0 U2901 ( .I(n3018), .Z(n3019) );
  CKBD0 U2902 ( .CLK(n3019), .C(n3020) );
  CKBD0 U2903 ( .CLK(n3020), .C(n3021) );
  CKBD0 U2904 ( .CLK(n3021), .C(n3022) );
  CKBD0 U2905 ( .CLK(n3022), .C(n3023) );
  CKBD0 U2906 ( .CLK(n3023), .C(n3024) );
  CKBD0 U2907 ( .CLK(n3024), .C(n3025) );
  CKBD0 U2908 ( .CLK(n3025), .C(n3026) );
  CKBD0 U2909 ( .CLK(n3026), .C(n3027) );
  CKBD0 U2910 ( .CLK(n3027), .C(n3028) );
  CKBD0 U2911 ( .CLK(n3028), .C(n3029) );
  BUFFD0 U2912 ( .I(n3029), .Z(n3030) );
  CKBD0 U2913 ( .CLK(n3030), .C(n3031) );
  CKBD0 U2914 ( .CLK(n3031), .C(n3032) );
  CKBD0 U2915 ( .CLK(n3032), .C(n3033) );
  CKBD0 U2916 ( .CLK(n3033), .C(n3034) );
  CKBD0 U2917 ( .CLK(n3034), .C(n3035) );
  CKBD0 U2918 ( .CLK(n3035), .C(n3036) );
  CKBD0 U2919 ( .CLK(n3036), .C(n3037) );
  CKBD0 U2920 ( .CLK(n3037), .C(n3038) );
  CKBD0 U2921 ( .CLK(n3038), .C(n3039) );
  CKBD0 U2922 ( .CLK(n3039), .C(n3040) );
  BUFFD0 U2923 ( .I(n3040), .Z(n3041) );
  CKBD0 U2924 ( .CLK(n3041), .C(n3042) );
  CKBD0 U2925 ( .CLK(n3042), .C(n3043) );
  CKBD0 U2926 ( .CLK(n3043), .C(n3044) );
  CKBD0 U2927 ( .CLK(n3044), .C(n3045) );
  CKBD0 U2928 ( .CLK(n3045), .C(n3046) );
  CKBD0 U2929 ( .CLK(n3046), .C(n3047) );
  CKBD0 U2930 ( .CLK(n3047), .C(n3048) );
  CKBD0 U2931 ( .CLK(n3048), .C(n3049) );
  CKBD0 U2932 ( .CLK(n3049), .C(n3050) );
  BUFFD0 U2933 ( .I(n3050), .Z(n3051) );
  CKBD0 U2934 ( .CLK(n3051), .C(n3052) );
  CKBD0 U2935 ( .CLK(n3052), .C(n3053) );
  CKBD0 U2936 ( .CLK(n3053), .C(n3054) );
  CKBD0 U2937 ( .CLK(n3054), .C(n3055) );
  CKBD0 U2938 ( .CLK(n3055), .C(n3056) );
  CKBD0 U2939 ( .CLK(n3056), .C(n3057) );
  CKBD0 U2940 ( .CLK(n3057), .C(n3058) );
  CKBD0 U2941 ( .CLK(n3058), .C(n3059) );
  CKBD0 U2942 ( .CLK(n3059), .C(n3060) );
  CKBD0 U2943 ( .CLK(n3060), .C(n3061) );
  CKBD0 U2944 ( .CLK(n3061), .C(n3062) );
  BUFFD0 U2945 ( .I(n3062), .Z(n3063) );
  CKBD0 U2946 ( .CLK(n3063), .C(n3064) );
  CKBD0 U2947 ( .CLK(n3064), .C(n3065) );
  CKBD0 U2948 ( .CLK(n3065), .C(n3066) );
  CKBD0 U2949 ( .CLK(n3066), .C(n3067) );
  CKBD0 U2950 ( .CLK(n3067), .C(n3068) );
  CKBD0 U2951 ( .CLK(n3068), .C(n3069) );
  CKBD0 U2952 ( .CLK(n3069), .C(n3070) );
  CKBD0 U2953 ( .CLK(n3070), .C(n3071) );
  CKBD0 U2954 ( .CLK(n3071), .C(n3072) );
  CKBD0 U2955 ( .CLK(n3072), .C(n3073) );
  BUFFD0 U2956 ( .I(n3073), .Z(n3074) );
  CKBD0 U2957 ( .CLK(n3074), .C(n3075) );
  CKBD0 U2958 ( .CLK(n3075), .C(n3076) );
  CKBD0 U2959 ( .CLK(n3076), .C(n3077) );
  CKBD0 U2960 ( .CLK(n3077), .C(n3078) );
  CKBD0 U2961 ( .CLK(n3078), .C(n3079) );
  CKBD0 U2962 ( .CLK(n3079), .C(n3080) );
  CKBD0 U2963 ( .CLK(n3080), .C(n3081) );
  CKBD0 U2964 ( .CLK(n3081), .C(n3082) );
  CKBD0 U2965 ( .CLK(n3082), .C(n3083) );
  BUFFD0 U2966 ( .I(n3083), .Z(n3084) );
  CKBD0 U2967 ( .CLK(n3084), .C(n3085) );
  CKBD0 U2968 ( .CLK(n3085), .C(n3086) );
  CKBD0 U2969 ( .CLK(n3086), .C(n3087) );
  CKBD0 U2970 ( .CLK(n3087), .C(n3088) );
  CKBD0 U2971 ( .CLK(n3088), .C(n3089) );
  CKBD0 U2972 ( .CLK(n3089), .C(n3090) );
  CKBD0 U2973 ( .CLK(n3090), .C(n3091) );
  CKBD0 U2974 ( .CLK(n3091), .C(n3092) );
  CKBD0 U2975 ( .CLK(n3092), .C(n3093) );
  CKBD0 U2976 ( .CLK(n3093), .C(n3094) );
  CKBD0 U2977 ( .CLK(n3094), .C(n3095) );
  BUFFD0 U2978 ( .I(n3095), .Z(n3096) );
  CKBD0 U2979 ( .CLK(n3096), .C(n3097) );
  CKBD0 U2980 ( .CLK(n3097), .C(n3098) );
  CKBD0 U2981 ( .CLK(n3098), .C(n3099) );
  CKBD0 U2982 ( .CLK(n3099), .C(n3100) );
  CKBD0 U2983 ( .CLK(n3100), .C(n3101) );
  CKBD0 U2984 ( .CLK(n3101), .C(n3102) );
  CKBD0 U2985 ( .CLK(n3102), .C(n3103) );
  CKBD0 U2986 ( .CLK(n3103), .C(n3104) );
  CKBD0 U2987 ( .CLK(n3104), .C(n3105) );
  BUFFD0 U2988 ( .I(n3105), .Z(n3106) );
  CKBD0 U2989 ( .CLK(n3106), .C(n3107) );
  CKBD0 U2990 ( .CLK(n3107), .C(n3108) );
  CKBD0 U2991 ( .CLK(n3108), .C(n3109) );
  CKBD0 U2992 ( .CLK(n3109), .C(n3110) );
  CKBD0 U2993 ( .CLK(n3110), .C(n3111) );
  CKBD0 U2994 ( .CLK(n3111), .C(n3112) );
  CKBD0 U2995 ( .CLK(n3112), .C(n3113) );
  CKBD0 U2996 ( .CLK(n3113), .C(n3114) );
  CKBD0 U2997 ( .CLK(n3114), .C(n3115) );
  BUFFD0 U2998 ( .I(n3115), .Z(n3116) );
  CKBD0 U2999 ( .CLK(n3116), .C(n3117) );
  CKBD0 U3000 ( .CLK(n3117), .C(n3118) );
  CKBD0 U3001 ( .CLK(n3118), .C(n3119) );
  CKBD0 U3002 ( .CLK(n3119), .C(n3120) );
  CKBD0 U3003 ( .CLK(n3120), .C(n3121) );
  CKBD0 U3004 ( .CLK(n3121), .C(n3122) );
  CKBD0 U3005 ( .CLK(n3122), .C(n3123) );
  CKBD0 U3006 ( .CLK(n3123), .C(n3124) );
  CKBD0 U3007 ( .CLK(n3124), .C(n3125) );
  CKBD0 U3008 ( .CLK(n3125), .C(n3126) );
  CKBD0 U3009 ( .CLK(n3126), .C(n3127) );
  BUFFD0 U3010 ( .I(n3127), .Z(n3128) );
  CKBD0 U3011 ( .CLK(n3128), .C(n3129) );
  CKBD0 U3012 ( .CLK(n3129), .C(n3130) );
  CKBD0 U3013 ( .CLK(n3130), .C(n3131) );
  CKBD0 U3014 ( .CLK(n3131), .C(n3132) );
  CKBD0 U3015 ( .CLK(n3132), .C(n3133) );
  BUFFD0 U3016 ( .I(n3133), .Z(n3134) );
  CKBD0 U3017 ( .CLK(n3134), .C(n3135) );
  BUFFD0 U3018 ( .I(n3135), .Z(n3136) );
  CKBD0 U3019 ( .CLK(n3136), .C(n3137) );
  BUFFD0 U3020 ( .I(n3137), .Z(n3138) );
  CKBD0 U3021 ( .CLK(n3138), .C(n3139) );
  BUFFD0 U3022 ( .I(n3139), .Z(n3140) );
  CKBD0 U3023 ( .CLK(n3140), .C(n3141) );
  BUFFD0 U3024 ( .I(n3141), .Z(n3142) );
  CKBD0 U3025 ( .CLK(n3142), .C(n3143) );
  BUFFD0 U3026 ( .I(n3143), .Z(n3144) );
  CKBD0 U3027 ( .CLK(n3144), .C(n3145) );
  BUFFD0 U3028 ( .I(n3145), .Z(n3146) );
  CKBD0 U3029 ( .CLK(n3146), .C(n3147) );
  BUFFD0 U3030 ( .I(n3147), .Z(n3148) );
  BUFFD0 U3031 ( .I(n3150), .Z(n3149) );
  BUFFD0 U3032 ( .I(n3151), .Z(n3150) );
  BUFFD0 U3033 ( .I(n9172), .Z(n3151) );
  CKBD0 U3034 ( .CLK(n1385), .C(n3152) );
  CKBD0 U3035 ( .CLK(n3152), .C(n3153) );
  CKBD0 U3036 ( .CLK(n3153), .C(n3154) );
  BUFFD0 U3037 ( .I(n3154), .Z(n3155) );
  CKBD0 U3038 ( .CLK(n3155), .C(n3156) );
  CKBD0 U3039 ( .CLK(n3156), .C(n3157) );
  CKBD0 U3040 ( .CLK(n3157), .C(n3158) );
  CKBD0 U3041 ( .CLK(n3158), .C(n3159) );
  CKBD0 U3042 ( .CLK(n3159), .C(n3160) );
  CKBD0 U3043 ( .CLK(n3160), .C(n3161) );
  CKBD0 U3044 ( .CLK(n3161), .C(n3162) );
  CKBD0 U3045 ( .CLK(n3162), .C(n3163) );
  CKBD0 U3046 ( .CLK(n3163), .C(n3164) );
  CKBD0 U3047 ( .CLK(n3164), .C(n3165) );
  BUFFD0 U3048 ( .I(n3165), .Z(n3166) );
  CKBD0 U3049 ( .CLK(n3166), .C(n3167) );
  CKBD0 U3050 ( .CLK(n3167), .C(n3168) );
  CKBD0 U3051 ( .CLK(n3168), .C(n3169) );
  CKBD0 U3052 ( .CLK(n3169), .C(n3170) );
  CKBD0 U3053 ( .CLK(n3170), .C(n3171) );
  CKBD0 U3054 ( .CLK(n3171), .C(n3172) );
  CKBD0 U3055 ( .CLK(n3172), .C(n3173) );
  CKBD0 U3056 ( .CLK(n3173), .C(n3174) );
  CKBD0 U3057 ( .CLK(n3174), .C(n3175) );
  CKBD0 U3058 ( .CLK(n3175), .C(n3176) );
  BUFFD0 U3059 ( .I(n3176), .Z(n3177) );
  CKBD0 U3060 ( .CLK(n3177), .C(n3178) );
  CKBD0 U3061 ( .CLK(n3178), .C(n3179) );
  CKBD0 U3062 ( .CLK(n3179), .C(n3180) );
  CKBD0 U3063 ( .CLK(n3180), .C(n3181) );
  CKBD0 U3064 ( .CLK(n3181), .C(n3182) );
  CKBD0 U3065 ( .CLK(n3182), .C(n3183) );
  CKBD0 U3066 ( .CLK(n3183), .C(n3184) );
  CKBD0 U3067 ( .CLK(n3184), .C(n3185) );
  CKBD0 U3068 ( .CLK(n3185), .C(n3186) );
  BUFFD0 U3069 ( .I(n3186), .Z(n3187) );
  CKBD0 U3070 ( .CLK(n3187), .C(n3188) );
  CKBD0 U3071 ( .CLK(n3188), .C(n3189) );
  CKBD0 U3072 ( .CLK(n3189), .C(n3190) );
  CKBD0 U3073 ( .CLK(n3190), .C(n3191) );
  CKBD0 U3074 ( .CLK(n3191), .C(n3192) );
  CKBD0 U3075 ( .CLK(n3192), .C(n3193) );
  CKBD0 U3076 ( .CLK(n3193), .C(n3194) );
  CKBD0 U3077 ( .CLK(n3194), .C(n3195) );
  CKBD0 U3078 ( .CLK(n3195), .C(n3196) );
  CKBD0 U3079 ( .CLK(n3196), .C(n3197) );
  CKBD0 U3080 ( .CLK(n3197), .C(n3198) );
  BUFFD0 U3081 ( .I(n3198), .Z(n3199) );
  CKBD0 U3082 ( .CLK(n3199), .C(n3200) );
  CKBD0 U3083 ( .CLK(n3200), .C(n3201) );
  CKBD0 U3084 ( .CLK(n3201), .C(n3202) );
  CKBD0 U3085 ( .CLK(n3202), .C(n3203) );
  CKBD0 U3086 ( .CLK(n3203), .C(n3204) );
  CKBD0 U3087 ( .CLK(n3204), .C(n3205) );
  CKBD0 U3088 ( .CLK(n3205), .C(n3206) );
  CKBD0 U3089 ( .CLK(n3206), .C(n3207) );
  CKBD0 U3090 ( .CLK(n3207), .C(n3208) );
  BUFFD0 U3091 ( .I(n3208), .Z(n3209) );
  CKBD0 U3092 ( .CLK(n3209), .C(n3210) );
  CKBD0 U3093 ( .CLK(n3210), .C(n3211) );
  CKBD0 U3094 ( .CLK(n3211), .C(n3212) );
  CKBD0 U3095 ( .CLK(n3212), .C(n3213) );
  CKBD0 U3096 ( .CLK(n3213), .C(n3214) );
  CKBD0 U3097 ( .CLK(n3214), .C(n3215) );
  CKBD0 U3098 ( .CLK(n3215), .C(n3216) );
  CKBD0 U3099 ( .CLK(n3216), .C(n3217) );
  CKBD0 U3100 ( .CLK(n3217), .C(n3218) );
  CKBD0 U3101 ( .CLK(n3218), .C(n3219) );
  BUFFD0 U3102 ( .I(n3219), .Z(n3220) );
  CKBD0 U3103 ( .CLK(n3220), .C(n3221) );
  CKBD0 U3104 ( .CLK(n3221), .C(n3222) );
  CKBD0 U3105 ( .CLK(n3222), .C(n3223) );
  CKBD0 U3106 ( .CLK(n3223), .C(n3224) );
  CKBD0 U3107 ( .CLK(n3224), .C(n3225) );
  CKBD0 U3108 ( .CLK(n3225), .C(n3226) );
  CKBD0 U3109 ( .CLK(n3226), .C(n3227) );
  CKBD0 U3110 ( .CLK(n3227), .C(n3228) );
  CKBD0 U3111 ( .CLK(n3228), .C(n3229) );
  CKBD0 U3112 ( .CLK(n3229), .C(n3230) );
  BUFFD0 U3113 ( .I(n3230), .Z(n3231) );
  CKBD0 U3114 ( .CLK(n3231), .C(n3232) );
  CKBD0 U3115 ( .CLK(n3232), .C(n3233) );
  CKBD0 U3116 ( .CLK(n3233), .C(n3234) );
  CKBD0 U3117 ( .CLK(n3234), .C(n3235) );
  CKBD0 U3118 ( .CLK(n3235), .C(n3236) );
  CKBD0 U3119 ( .CLK(n3236), .C(n3237) );
  CKBD0 U3120 ( .CLK(n3237), .C(n3238) );
  CKBD0 U3121 ( .CLK(n3238), .C(n3239) );
  CKBD0 U3122 ( .CLK(n3239), .C(n3240) );
  CKBD0 U3123 ( .CLK(n3240), .C(n3241) );
  BUFFD0 U3124 ( .I(n3241), .Z(n3242) );
  CKBD0 U3125 ( .CLK(n3242), .C(n3243) );
  CKBD0 U3126 ( .CLK(n3243), .C(n3244) );
  CKBD0 U3127 ( .CLK(n3244), .C(n3245) );
  CKBD0 U3128 ( .CLK(n3245), .C(n3246) );
  CKBD0 U3129 ( .CLK(n3246), .C(n3247) );
  CKBD0 U3130 ( .CLK(n3247), .C(n3248) );
  CKBD0 U3131 ( .CLK(n3248), .C(n3249) );
  CKBD0 U3132 ( .CLK(n3249), .C(n3250) );
  CKBD0 U3133 ( .CLK(n3250), .C(n3251) );
  CKBD0 U3134 ( .CLK(n3251), .C(n3252) );
  BUFFD0 U3135 ( .I(n3252), .Z(n3253) );
  CKBD0 U3136 ( .CLK(n3253), .C(n3254) );
  CKBD0 U3137 ( .CLK(n3254), .C(n3255) );
  CKBD0 U3138 ( .CLK(n3255), .C(n3256) );
  CKBD0 U3139 ( .CLK(n3256), .C(n3257) );
  CKBD0 U3140 ( .CLK(n3257), .C(n3258) );
  CKBD0 U3141 ( .CLK(n3258), .C(n3259) );
  CKBD0 U3142 ( .CLK(n3259), .C(n3260) );
  CKBD0 U3143 ( .CLK(n3260), .C(n3261) );
  CKBD0 U3144 ( .CLK(n3261), .C(n3262) );
  CKBD0 U3145 ( .CLK(n3262), .C(n3263) );
  BUFFD0 U3146 ( .I(n3263), .Z(n3264) );
  CKBD0 U3147 ( .CLK(n3264), .C(n3265) );
  CKBD0 U3148 ( .CLK(n3265), .C(n3266) );
  CKBD0 U3149 ( .CLK(n3266), .C(n3267) );
  CKBD0 U3150 ( .CLK(n3267), .C(n3268) );
  CKBD0 U3151 ( .CLK(n3268), .C(n3269) );
  BUFFD0 U3152 ( .I(n3269), .Z(n3270) );
  CKBD0 U3153 ( .CLK(n3270), .C(n3271) );
  BUFFD0 U3154 ( .I(n3271), .Z(n3272) );
  CKBD0 U3155 ( .CLK(n3272), .C(n3273) );
  BUFFD0 U3156 ( .I(n3273), .Z(n3274) );
  CKBD0 U3157 ( .CLK(n3274), .C(n3275) );
  BUFFD0 U3158 ( .I(n3275), .Z(n3276) );
  CKBD0 U3159 ( .CLK(n3276), .C(n3277) );
  BUFFD0 U3160 ( .I(n3277), .Z(n3278) );
  CKBD0 U3161 ( .CLK(n3278), .C(n3279) );
  BUFFD0 U3162 ( .I(n3279), .Z(n3280) );
  CKBD0 U3163 ( .CLK(n3280), .C(n3281) );
  BUFFD0 U3164 ( .I(n3281), .Z(n3282) );
  CKBD0 U3165 ( .CLK(n3282), .C(n3283) );
  BUFFD0 U3166 ( .I(n3283), .Z(n3284) );
  BUFFD0 U3167 ( .I(n3286), .Z(n3285) );
  BUFFD0 U3168 ( .I(n3287), .Z(n3286) );
  BUFFD0 U3169 ( .I(n9173), .Z(n3287) );
  CKBD0 U3170 ( .CLK(n1383), .C(n3288) );
  CKBD0 U3171 ( .CLK(n3288), .C(n3289) );
  CKBD0 U3172 ( .CLK(n3289), .C(n3290) );
  BUFFD0 U3173 ( .I(n3290), .Z(n3291) );
  CKBD0 U3174 ( .CLK(n3291), .C(n3292) );
  CKBD0 U3175 ( .CLK(n3292), .C(n3293) );
  CKBD0 U3176 ( .CLK(n3293), .C(n3294) );
  CKBD0 U3177 ( .CLK(n3294), .C(n3295) );
  CKBD0 U3178 ( .CLK(n3295), .C(n3296) );
  CKBD0 U3179 ( .CLK(n3296), .C(n3297) );
  CKBD0 U3180 ( .CLK(n3297), .C(n3298) );
  CKBD0 U3181 ( .CLK(n3298), .C(n3299) );
  CKBD0 U3182 ( .CLK(n3299), .C(n3300) );
  CKBD0 U3183 ( .CLK(n3300), .C(n3301) );
  BUFFD0 U3184 ( .I(n3301), .Z(n3302) );
  CKBD0 U3185 ( .CLK(n3302), .C(n3303) );
  CKBD0 U3186 ( .CLK(n3303), .C(n3304) );
  CKBD0 U3187 ( .CLK(n3304), .C(n3305) );
  CKBD0 U3188 ( .CLK(n3305), .C(n3306) );
  CKBD0 U3189 ( .CLK(n3306), .C(n3307) );
  CKBD0 U3190 ( .CLK(n3307), .C(n3308) );
  CKBD0 U3191 ( .CLK(n3308), .C(n3309) );
  CKBD0 U3192 ( .CLK(n3309), .C(n3310) );
  CKBD0 U3193 ( .CLK(n3310), .C(n3311) );
  CKBD0 U3194 ( .CLK(n3311), .C(n3312) );
  BUFFD0 U3195 ( .I(n3312), .Z(n3313) );
  CKBD0 U3196 ( .CLK(n3313), .C(n3314) );
  CKBD0 U3197 ( .CLK(n3314), .C(n3315) );
  CKBD0 U3198 ( .CLK(n3315), .C(n3316) );
  CKBD0 U3199 ( .CLK(n3316), .C(n3317) );
  CKBD0 U3200 ( .CLK(n3317), .C(n3318) );
  CKBD0 U3201 ( .CLK(n3318), .C(n3319) );
  CKBD0 U3202 ( .CLK(n3319), .C(n3320) );
  CKBD0 U3203 ( .CLK(n3320), .C(n3321) );
  CKBD0 U3204 ( .CLK(n3321), .C(n3322) );
  CKBD0 U3205 ( .CLK(n3322), .C(n3323) );
  BUFFD0 U3206 ( .I(n3323), .Z(n3324) );
  CKBD0 U3207 ( .CLK(n3324), .C(n3325) );
  CKBD0 U3208 ( .CLK(n3325), .C(n3326) );
  CKBD0 U3209 ( .CLK(n3326), .C(n3327) );
  CKBD0 U3210 ( .CLK(n3327), .C(n3328) );
  CKBD0 U3211 ( .CLK(n3328), .C(n3329) );
  CKBD0 U3212 ( .CLK(n3329), .C(n3330) );
  CKBD0 U3213 ( .CLK(n3330), .C(n3331) );
  CKBD0 U3214 ( .CLK(n3331), .C(n3332) );
  CKBD0 U3215 ( .CLK(n3332), .C(n3333) );
  CKBD0 U3216 ( .CLK(n3333), .C(n3334) );
  BUFFD0 U3217 ( .I(n3334), .Z(n3335) );
  CKBD0 U3218 ( .CLK(n3335), .C(n3336) );
  CKBD0 U3219 ( .CLK(n3336), .C(n3337) );
  CKBD0 U3220 ( .CLK(n3337), .C(n3338) );
  CKBD0 U3221 ( .CLK(n3338), .C(n3339) );
  CKBD0 U3222 ( .CLK(n3339), .C(n3340) );
  CKBD0 U3223 ( .CLK(n3340), .C(n3341) );
  CKBD0 U3224 ( .CLK(n3341), .C(n3342) );
  CKBD0 U3225 ( .CLK(n3342), .C(n3343) );
  CKBD0 U3226 ( .CLK(n3343), .C(n3344) );
  BUFFD0 U3227 ( .I(n3344), .Z(n3345) );
  CKBD0 U3228 ( .CLK(n3345), .C(n3346) );
  CKBD0 U3229 ( .CLK(n3346), .C(n3347) );
  CKBD0 U3230 ( .CLK(n3347), .C(n3348) );
  CKBD0 U3231 ( .CLK(n3348), .C(n3349) );
  CKBD0 U3232 ( .CLK(n3349), .C(n3350) );
  CKBD0 U3233 ( .CLK(n3350), .C(n3351) );
  CKBD0 U3234 ( .CLK(n3351), .C(n3352) );
  CKBD0 U3235 ( .CLK(n3352), .C(n3353) );
  CKBD0 U3236 ( .CLK(n3353), .C(n3354) );
  CKBD0 U3237 ( .CLK(n3354), .C(n3355) );
  CKBD0 U3238 ( .CLK(n3355), .C(n3356) );
  BUFFD0 U3239 ( .I(n3356), .Z(n3357) );
  CKBD0 U3240 ( .CLK(n3357), .C(n3358) );
  CKBD0 U3241 ( .CLK(n3358), .C(n3359) );
  CKBD0 U3242 ( .CLK(n3359), .C(n3360) );
  CKBD0 U3243 ( .CLK(n3360), .C(n3361) );
  CKBD0 U3244 ( .CLK(n3361), .C(n3362) );
  CKBD0 U3245 ( .CLK(n3362), .C(n3363) );
  CKBD0 U3246 ( .CLK(n3363), .C(n3364) );
  CKBD0 U3247 ( .CLK(n3364), .C(n3365) );
  CKBD0 U3248 ( .CLK(n3365), .C(n3366) );
  BUFFD0 U3249 ( .I(n3366), .Z(n3367) );
  CKBD0 U3250 ( .CLK(n3367), .C(n3368) );
  CKBD0 U3251 ( .CLK(n3368), .C(n3369) );
  CKBD0 U3252 ( .CLK(n3369), .C(n3370) );
  CKBD0 U3253 ( .CLK(n3370), .C(n3371) );
  CKBD0 U3254 ( .CLK(n3371), .C(n3372) );
  CKBD0 U3255 ( .CLK(n3372), .C(n3373) );
  CKBD0 U3256 ( .CLK(n3373), .C(n3374) );
  CKBD0 U3257 ( .CLK(n3374), .C(n3375) );
  CKBD0 U3258 ( .CLK(n3375), .C(n3376) );
  CKBD0 U3259 ( .CLK(n3376), .C(n3377) );
  BUFFD0 U3260 ( .I(n3377), .Z(n3378) );
  CKBD0 U3261 ( .CLK(n3378), .C(n3379) );
  CKBD0 U3262 ( .CLK(n3379), .C(n3380) );
  CKBD0 U3263 ( .CLK(n3380), .C(n3381) );
  CKBD0 U3264 ( .CLK(n3381), .C(n3382) );
  CKBD0 U3265 ( .CLK(n3382), .C(n3383) );
  CKBD0 U3266 ( .CLK(n3383), .C(n3384) );
  CKBD0 U3267 ( .CLK(n3384), .C(n3385) );
  CKBD0 U3268 ( .CLK(n3385), .C(n3386) );
  CKBD0 U3269 ( .CLK(n3386), .C(n3387) );
  CKBD0 U3270 ( .CLK(n3387), .C(n3388) );
  BUFFD0 U3271 ( .I(n3388), .Z(n3389) );
  CKBD0 U3272 ( .CLK(n3389), .C(n3390) );
  CKBD0 U3273 ( .CLK(n3390), .C(n3391) );
  CKBD0 U3274 ( .CLK(n3391), .C(n3392) );
  CKBD0 U3275 ( .CLK(n3392), .C(n3393) );
  CKBD0 U3276 ( .CLK(n3393), .C(n3394) );
  CKBD0 U3277 ( .CLK(n3394), .C(n3395) );
  CKBD0 U3278 ( .CLK(n3395), .C(n3396) );
  CKBD0 U3279 ( .CLK(n3396), .C(n3397) );
  CKBD0 U3280 ( .CLK(n3397), .C(n3398) );
  CKBD0 U3281 ( .CLK(n3398), .C(n3399) );
  BUFFD0 U3282 ( .I(n3399), .Z(n3400) );
  CKBD0 U3283 ( .CLK(n3400), .C(n3401) );
  CKBD0 U3284 ( .CLK(n3401), .C(n3402) );
  CKBD0 U3285 ( .CLK(n3402), .C(n3403) );
  CKBD0 U3286 ( .CLK(n3403), .C(n3404) );
  CKBD0 U3287 ( .CLK(n3404), .C(n3405) );
  BUFFD0 U3288 ( .I(n3405), .Z(n3406) );
  CKBD0 U3289 ( .CLK(n3406), .C(n3407) );
  BUFFD0 U3290 ( .I(n3407), .Z(n3408) );
  CKBD0 U3291 ( .CLK(n3408), .C(n3409) );
  BUFFD0 U3292 ( .I(n3409), .Z(n3410) );
  CKBD0 U3293 ( .CLK(n3410), .C(n3411) );
  BUFFD0 U3294 ( .I(n3411), .Z(n3412) );
  CKBD0 U3295 ( .CLK(n3412), .C(n3413) );
  BUFFD0 U3296 ( .I(n3413), .Z(n3414) );
  CKBD0 U3297 ( .CLK(n3414), .C(n3415) );
  BUFFD0 U3298 ( .I(n3415), .Z(n3416) );
  CKBD0 U3299 ( .CLK(n3416), .C(n3417) );
  BUFFD0 U3300 ( .I(n3417), .Z(n3418) );
  CKBD0 U3301 ( .CLK(n3418), .C(n3419) );
  BUFFD0 U3302 ( .I(n3419), .Z(n3420) );
  BUFFD0 U3303 ( .I(n3422), .Z(n3421) );
  BUFFD0 U3304 ( .I(n3423), .Z(n3422) );
  BUFFD0 U3305 ( .I(n9174), .Z(n3423) );
  CKBD0 U3306 ( .CLK(n1381), .C(n3424) );
  CKBD0 U3307 ( .CLK(n3424), .C(n3425) );
  CKBD0 U3308 ( .CLK(n3425), .C(n3426) );
  CKBD0 U3309 ( .CLK(n3426), .C(n3427) );
  BUFFD0 U3310 ( .I(n3427), .Z(n3428) );
  CKBD0 U3311 ( .CLK(n3428), .C(n3429) );
  CKBD0 U3312 ( .CLK(n3429), .C(n3430) );
  CKBD0 U3313 ( .CLK(n3430), .C(n3431) );
  CKBD0 U3314 ( .CLK(n3431), .C(n3432) );
  CKBD0 U3315 ( .CLK(n3432), .C(n3433) );
  CKBD0 U3316 ( .CLK(n3433), .C(n3434) );
  CKBD0 U3317 ( .CLK(n3434), .C(n3435) );
  CKBD0 U3318 ( .CLK(n3435), .C(n3436) );
  CKBD0 U3319 ( .CLK(n3436), .C(n3437) );
  BUFFD0 U3320 ( .I(n3437), .Z(n3438) );
  CKBD0 U3321 ( .CLK(n3438), .C(n3439) );
  CKBD0 U3322 ( .CLK(n3439), .C(n3440) );
  CKBD0 U3323 ( .CLK(n3440), .C(n3441) );
  CKBD0 U3324 ( .CLK(n3441), .C(n3442) );
  CKBD0 U3325 ( .CLK(n3442), .C(n3443) );
  CKBD0 U3326 ( .CLK(n3443), .C(n3444) );
  CKBD0 U3327 ( .CLK(n3444), .C(n3445) );
  CKBD0 U3328 ( .CLK(n3445), .C(n3446) );
  CKBD0 U3329 ( .CLK(n3446), .C(n3447) );
  BUFFD0 U3330 ( .I(n3447), .Z(n3448) );
  CKBD0 U3331 ( .CLK(n3448), .C(n3449) );
  CKBD0 U3332 ( .CLK(n3449), .C(n3450) );
  CKBD0 U3333 ( .CLK(n3450), .C(n3451) );
  CKBD0 U3334 ( .CLK(n3451), .C(n3452) );
  CKBD0 U3335 ( .CLK(n3452), .C(n3453) );
  CKBD0 U3336 ( .CLK(n3453), .C(n3454) );
  CKBD0 U3337 ( .CLK(n3454), .C(n3455) );
  CKBD0 U3338 ( .CLK(n3455), .C(n3456) );
  CKBD0 U3339 ( .CLK(n3456), .C(n3457) );
  CKBD0 U3340 ( .CLK(n3457), .C(n3458) );
  CKBD0 U3341 ( .CLK(n3458), .C(n3459) );
  BUFFD0 U3342 ( .I(n3459), .Z(n3460) );
  CKBD0 U3343 ( .CLK(n3460), .C(n3461) );
  CKBD0 U3344 ( .CLK(n3461), .C(n3462) );
  CKBD0 U3345 ( .CLK(n3462), .C(n3463) );
  CKBD0 U3346 ( .CLK(n3463), .C(n3464) );
  CKBD0 U3347 ( .CLK(n3464), .C(n3465) );
  CKBD0 U3348 ( .CLK(n3465), .C(n3466) );
  CKBD0 U3349 ( .CLK(n3466), .C(n3467) );
  CKBD0 U3350 ( .CLK(n3467), .C(n3468) );
  CKBD0 U3351 ( .CLK(n3468), .C(n3469) );
  CKBD0 U3352 ( .CLK(n3469), .C(n3470) );
  BUFFD0 U3353 ( .I(n3470), .Z(n3471) );
  CKBD0 U3354 ( .CLK(n3471), .C(n3472) );
  CKBD0 U3355 ( .CLK(n3472), .C(n3473) );
  CKBD0 U3356 ( .CLK(n3473), .C(n3474) );
  CKBD0 U3357 ( .CLK(n3474), .C(n3475) );
  CKBD0 U3358 ( .CLK(n3475), .C(n3476) );
  CKBD0 U3359 ( .CLK(n3476), .C(n3477) );
  CKBD0 U3360 ( .CLK(n3477), .C(n3478) );
  CKBD0 U3361 ( .CLK(n3478), .C(n3479) );
  CKBD0 U3362 ( .CLK(n3479), .C(n3480) );
  BUFFD0 U3363 ( .I(n3480), .Z(n3481) );
  CKBD0 U3364 ( .CLK(n3481), .C(n3482) );
  CKBD0 U3365 ( .CLK(n3482), .C(n3483) );
  CKBD0 U3366 ( .CLK(n3483), .C(n3484) );
  CKBD0 U3367 ( .CLK(n3484), .C(n3485) );
  CKBD0 U3368 ( .CLK(n3485), .C(n3486) );
  CKBD0 U3369 ( .CLK(n3486), .C(n3487) );
  CKBD0 U3370 ( .CLK(n3487), .C(n3488) );
  CKBD0 U3371 ( .CLK(n3488), .C(n3489) );
  CKBD0 U3372 ( .CLK(n3489), .C(n3490) );
  CKBD0 U3373 ( .CLK(n3490), .C(n3491) );
  CKBD0 U3374 ( .CLK(n3491), .C(n3492) );
  BUFFD0 U3375 ( .I(n3492), .Z(n3493) );
  CKBD0 U3376 ( .CLK(n3493), .C(n3494) );
  CKBD0 U3377 ( .CLK(n3494), .C(n3495) );
  CKBD0 U3378 ( .CLK(n3495), .C(n3496) );
  CKBD0 U3379 ( .CLK(n3496), .C(n3497) );
  CKBD0 U3380 ( .CLK(n3497), .C(n3498) );
  CKBD0 U3381 ( .CLK(n3498), .C(n3499) );
  CKBD0 U3382 ( .CLK(n3499), .C(n3500) );
  CKBD0 U3383 ( .CLK(n3500), .C(n3501) );
  CKBD0 U3384 ( .CLK(n3501), .C(n3502) );
  BUFFD0 U3385 ( .I(n3502), .Z(n3503) );
  CKBD0 U3386 ( .CLK(n3503), .C(n3504) );
  CKBD0 U3387 ( .CLK(n3504), .C(n3505) );
  CKBD0 U3388 ( .CLK(n3505), .C(n3506) );
  CKBD0 U3389 ( .CLK(n3506), .C(n3507) );
  CKBD0 U3390 ( .CLK(n3507), .C(n3508) );
  CKBD0 U3391 ( .CLK(n3508), .C(n3509) );
  CKBD0 U3392 ( .CLK(n3509), .C(n3510) );
  CKBD0 U3393 ( .CLK(n3510), .C(n3511) );
  CKBD0 U3394 ( .CLK(n3511), .C(n3512) );
  CKBD0 U3395 ( .CLK(n3512), .C(n3513) );
  BUFFD0 U3396 ( .I(n3513), .Z(n3514) );
  CKBD0 U3397 ( .CLK(n3514), .C(n3515) );
  CKBD0 U3398 ( .CLK(n3515), .C(n3516) );
  CKBD0 U3399 ( .CLK(n3516), .C(n3517) );
  CKBD0 U3400 ( .CLK(n3517), .C(n3518) );
  CKBD0 U3401 ( .CLK(n3518), .C(n3519) );
  CKBD0 U3402 ( .CLK(n3519), .C(n3520) );
  CKBD0 U3403 ( .CLK(n3520), .C(n3521) );
  CKBD0 U3404 ( .CLK(n3521), .C(n3522) );
  CKBD0 U3405 ( .CLK(n3522), .C(n3523) );
  CKBD0 U3406 ( .CLK(n3523), .C(n3524) );
  BUFFD0 U3407 ( .I(n3524), .Z(n3525) );
  CKBD0 U3408 ( .CLK(n3525), .C(n3526) );
  CKBD0 U3409 ( .CLK(n3526), .C(n3527) );
  CKBD0 U3410 ( .CLK(n3527), .C(n3528) );
  CKBD0 U3411 ( .CLK(n3528), .C(n3529) );
  CKBD0 U3412 ( .CLK(n3529), .C(n3530) );
  CKBD0 U3413 ( .CLK(n3530), .C(n3531) );
  CKBD0 U3414 ( .CLK(n3531), .C(n3532) );
  CKBD0 U3415 ( .CLK(n3532), .C(n3533) );
  CKBD0 U3416 ( .CLK(n3533), .C(n3534) );
  BUFFD0 U3417 ( .I(n3534), .Z(n3535) );
  CKBD0 U3418 ( .CLK(n3535), .C(n3536) );
  CKBD0 U3419 ( .CLK(n3536), .C(n3537) );
  CKBD0 U3420 ( .CLK(n3537), .C(n3538) );
  CKBD0 U3421 ( .CLK(n3538), .C(n3539) );
  CKBD0 U3422 ( .CLK(n3539), .C(n3540) );
  CKBD0 U3423 ( .CLK(n3540), .C(n3541) );
  BUFFD0 U3424 ( .I(n3541), .Z(n3542) );
  CKBD0 U3425 ( .CLK(n3542), .C(n3543) );
  BUFFD0 U3426 ( .I(n3543), .Z(n3544) );
  CKBD0 U3427 ( .CLK(n3544), .C(n3545) );
  BUFFD0 U3428 ( .I(n3545), .Z(n3546) );
  CKBD0 U3429 ( .CLK(n3546), .C(n3547) );
  BUFFD0 U3430 ( .I(n3547), .Z(n3548) );
  CKBD0 U3431 ( .CLK(n3548), .C(n3549) );
  BUFFD0 U3432 ( .I(n3549), .Z(n3550) );
  CKBD0 U3433 ( .CLK(n3550), .C(n3551) );
  BUFFD0 U3434 ( .I(n3551), .Z(n3552) );
  CKBD0 U3435 ( .CLK(n3552), .C(n3553) );
  BUFFD0 U3436 ( .I(n3553), .Z(n3554) );
  CKBD0 U3437 ( .CLK(n3554), .C(n3555) );
  BUFFD0 U3438 ( .I(n3555), .Z(n3556) );
  BUFFD0 U3439 ( .I(n3558), .Z(n3557) );
  BUFFD0 U3440 ( .I(n3559), .Z(n3558) );
  BUFFD0 U3441 ( .I(n9175), .Z(n3559) );
  CKBD0 U3442 ( .CLK(n1379), .C(n3560) );
  CKBD0 U3443 ( .CLK(n3560), .C(n3561) );
  CKBD0 U3444 ( .CLK(n3561), .C(n3562) );
  BUFFD0 U3445 ( .I(n3562), .Z(n3563) );
  CKBD0 U3446 ( .CLK(n3563), .C(n3564) );
  CKBD0 U3447 ( .CLK(n3564), .C(n3565) );
  CKBD0 U3448 ( .CLK(n3565), .C(n3566) );
  CKBD0 U3449 ( .CLK(n3566), .C(n3567) );
  CKBD0 U3450 ( .CLK(n3567), .C(n3568) );
  CKBD0 U3451 ( .CLK(n3568), .C(n3569) );
  CKBD0 U3452 ( .CLK(n3569), .C(n3570) );
  CKBD0 U3453 ( .CLK(n3570), .C(n3571) );
  CKBD0 U3454 ( .CLK(n3571), .C(n3572) );
  CKBD0 U3455 ( .CLK(n3572), .C(n3573) );
  BUFFD0 U3456 ( .I(n3573), .Z(n3574) );
  CKBD0 U3457 ( .CLK(n3574), .C(n3575) );
  CKBD0 U3458 ( .CLK(n3575), .C(n3576) );
  CKBD0 U3459 ( .CLK(n3576), .C(n3577) );
  CKBD0 U3460 ( .CLK(n3577), .C(n3578) );
  CKBD0 U3461 ( .CLK(n3578), .C(n3579) );
  CKBD0 U3462 ( .CLK(n3579), .C(n3580) );
  CKBD0 U3463 ( .CLK(n3580), .C(n3581) );
  CKBD0 U3464 ( .CLK(n3581), .C(n3582) );
  CKBD0 U3465 ( .CLK(n3582), .C(n3583) );
  CKBD0 U3466 ( .CLK(n3583), .C(n3584) );
  BUFFD0 U3467 ( .I(n3584), .Z(n3585) );
  CKBD0 U3468 ( .CLK(n3585), .C(n3586) );
  CKBD0 U3469 ( .CLK(n3586), .C(n3587) );
  CKBD0 U3470 ( .CLK(n3587), .C(n3588) );
  CKBD0 U3471 ( .CLK(n3588), .C(n3589) );
  CKBD0 U3472 ( .CLK(n3589), .C(n3590) );
  CKBD0 U3473 ( .CLK(n3590), .C(n3591) );
  CKBD0 U3474 ( .CLK(n3591), .C(n3592) );
  CKBD0 U3475 ( .CLK(n3592), .C(n3593) );
  CKBD0 U3476 ( .CLK(n3593), .C(n3594) );
  CKBD0 U3477 ( .CLK(n3594), .C(n3595) );
  BUFFD0 U3478 ( .I(n3595), .Z(n3596) );
  CKBD0 U3479 ( .CLK(n3596), .C(n3597) );
  CKBD0 U3480 ( .CLK(n3597), .C(n3598) );
  CKBD0 U3481 ( .CLK(n3598), .C(n3599) );
  CKBD0 U3482 ( .CLK(n3599), .C(n3600) );
  CKBD0 U3483 ( .CLK(n3600), .C(n3601) );
  CKBD0 U3484 ( .CLK(n3601), .C(n3602) );
  CKBD0 U3485 ( .CLK(n3602), .C(n3603) );
  CKBD0 U3486 ( .CLK(n3603), .C(n3604) );
  CKBD0 U3487 ( .CLK(n3604), .C(n3605) );
  BUFFD0 U3488 ( .I(n3605), .Z(n3606) );
  CKBD0 U3489 ( .CLK(n3606), .C(n3607) );
  CKBD0 U3490 ( .CLK(n3607), .C(n3608) );
  CKBD0 U3491 ( .CLK(n3608), .C(n3609) );
  CKBD0 U3492 ( .CLK(n3609), .C(n3610) );
  CKBD0 U3493 ( .CLK(n3610), .C(n3611) );
  CKBD0 U3494 ( .CLK(n3611), .C(n3612) );
  CKBD0 U3495 ( .CLK(n3612), .C(n3613) );
  CKBD0 U3496 ( .CLK(n3613), .C(n3614) );
  CKBD0 U3497 ( .CLK(n3614), .C(n3615) );
  CKBD0 U3498 ( .CLK(n3615), .C(n3616) );
  CKBD0 U3499 ( .CLK(n3616), .C(n3617) );
  BUFFD0 U3500 ( .I(n3617), .Z(n3618) );
  CKBD0 U3501 ( .CLK(n3618), .C(n3619) );
  CKBD0 U3502 ( .CLK(n3619), .C(n3620) );
  CKBD0 U3503 ( .CLK(n3620), .C(n3621) );
  CKBD0 U3504 ( .CLK(n3621), .C(n3622) );
  CKBD0 U3505 ( .CLK(n3622), .C(n3623) );
  CKBD0 U3506 ( .CLK(n3623), .C(n3624) );
  CKBD0 U3507 ( .CLK(n3624), .C(n3625) );
  CKBD0 U3508 ( .CLK(n3625), .C(n3626) );
  CKBD0 U3509 ( .CLK(n3626), .C(n3627) );
  BUFFD0 U3510 ( .I(n3627), .Z(n3628) );
  CKBD0 U3511 ( .CLK(n3628), .C(n3629) );
  CKBD0 U3512 ( .CLK(n3629), .C(n3630) );
  CKBD0 U3513 ( .CLK(n3630), .C(n3631) );
  CKBD0 U3514 ( .CLK(n3631), .C(n3632) );
  CKBD0 U3515 ( .CLK(n3632), .C(n3633) );
  CKBD0 U3516 ( .CLK(n3633), .C(n3634) );
  CKBD0 U3517 ( .CLK(n3634), .C(n3635) );
  CKBD0 U3518 ( .CLK(n3635), .C(n3636) );
  CKBD0 U3519 ( .CLK(n3636), .C(n3637) );
  CKBD0 U3520 ( .CLK(n3637), .C(n3638) );
  BUFFD0 U3521 ( .I(n3638), .Z(n3639) );
  CKBD0 U3522 ( .CLK(n3639), .C(n3640) );
  CKBD0 U3523 ( .CLK(n3640), .C(n3641) );
  CKBD0 U3524 ( .CLK(n3641), .C(n3642) );
  CKBD0 U3525 ( .CLK(n3642), .C(n3643) );
  CKBD0 U3526 ( .CLK(n3643), .C(n3644) );
  CKBD0 U3527 ( .CLK(n3644), .C(n3645) );
  CKBD0 U3528 ( .CLK(n3645), .C(n3646) );
  CKBD0 U3529 ( .CLK(n3646), .C(n3647) );
  CKBD0 U3530 ( .CLK(n3647), .C(n3648) );
  CKBD0 U3531 ( .CLK(n3648), .C(n3649) );
  BUFFD0 U3532 ( .I(n3649), .Z(n3650) );
  CKBD0 U3533 ( .CLK(n3650), .C(n3651) );
  CKBD0 U3534 ( .CLK(n3651), .C(n3652) );
  CKBD0 U3535 ( .CLK(n3652), .C(n3653) );
  CKBD0 U3536 ( .CLK(n3653), .C(n3654) );
  CKBD0 U3537 ( .CLK(n3654), .C(n3655) );
  CKBD0 U3538 ( .CLK(n3655), .C(n3656) );
  CKBD0 U3539 ( .CLK(n3656), .C(n3657) );
  CKBD0 U3540 ( .CLK(n3657), .C(n3658) );
  CKBD0 U3541 ( .CLK(n3658), .C(n3659) );
  CKBD0 U3542 ( .CLK(n3659), .C(n3660) );
  BUFFD0 U3543 ( .I(n3660), .Z(n3661) );
  CKBD0 U3544 ( .CLK(n3661), .C(n3662) );
  CKBD0 U3545 ( .CLK(n3662), .C(n3663) );
  CKBD0 U3546 ( .CLK(n3663), .C(n3664) );
  CKBD0 U3547 ( .CLK(n3664), .C(n3665) );
  CKBD0 U3548 ( .CLK(n3665), .C(n3666) );
  CKBD0 U3549 ( .CLK(n3666), .C(n3667) );
  CKBD0 U3550 ( .CLK(n3667), .C(n3668) );
  CKBD0 U3551 ( .CLK(n3668), .C(n3669) );
  CKBD0 U3552 ( .CLK(n3669), .C(n3670) );
  BUFFD0 U3553 ( .I(n3670), .Z(n3671) );
  CKBD0 U3554 ( .CLK(n3671), .C(n3672) );
  CKBD0 U3555 ( .CLK(n3672), .C(n3673) );
  CKBD0 U3556 ( .CLK(n3673), .C(n3674) );
  CKBD0 U3557 ( .CLK(n3674), .C(n3675) );
  CKBD0 U3558 ( .CLK(n3675), .C(n3676) );
  CKBD0 U3559 ( .CLK(n3676), .C(n3677) );
  BUFFD0 U3560 ( .I(n3677), .Z(n3678) );
  CKBD0 U3561 ( .CLK(n3678), .C(n3679) );
  BUFFD0 U3562 ( .I(n3679), .Z(n3680) );
  CKBD0 U3563 ( .CLK(n3680), .C(n3681) );
  BUFFD0 U3564 ( .I(n3681), .Z(n3682) );
  CKBD0 U3565 ( .CLK(n3682), .C(n3683) );
  BUFFD0 U3566 ( .I(n3683), .Z(n3684) );
  CKBD0 U3567 ( .CLK(n3684), .C(n3685) );
  BUFFD0 U3568 ( .I(n3685), .Z(n3686) );
  CKBD0 U3569 ( .CLK(n3686), .C(n3687) );
  BUFFD0 U3570 ( .I(n3687), .Z(n3688) );
  CKBD0 U3571 ( .CLK(n3688), .C(n3689) );
  BUFFD0 U3572 ( .I(n3689), .Z(n3690) );
  CKBD0 U3573 ( .CLK(n3690), .C(n3691) );
  BUFFD0 U3574 ( .I(n3691), .Z(n3692) );
  BUFFD0 U3575 ( .I(n3694), .Z(n3693) );
  BUFFD0 U3576 ( .I(n3695), .Z(n3694) );
  BUFFD0 U3577 ( .I(n9176), .Z(n3695) );
  CKBD0 U3578 ( .CLK(n1897), .C(n3696) );
  CKBD0 U3579 ( .CLK(n3696), .C(n3697) );
  CKBD0 U3580 ( .CLK(n3697), .C(n3698) );
  BUFFD0 U3581 ( .I(n3698), .Z(n3699) );
  CKBD0 U3582 ( .CLK(n3699), .C(n3700) );
  CKBD0 U3583 ( .CLK(n3700), .C(n3701) );
  CKBD0 U3584 ( .CLK(n3701), .C(n3702) );
  CKBD0 U3585 ( .CLK(n3702), .C(n3703) );
  CKBD0 U3586 ( .CLK(n3703), .C(n3704) );
  CKBD0 U3587 ( .CLK(n3704), .C(n3705) );
  CKBD0 U3588 ( .CLK(n3705), .C(n3706) );
  CKBD0 U3589 ( .CLK(n3706), .C(n3707) );
  CKBD0 U3590 ( .CLK(n3707), .C(n3708) );
  CKBD0 U3591 ( .CLK(n3708), .C(n3709) );
  BUFFD0 U3592 ( .I(n3709), .Z(n3710) );
  CKBD0 U3593 ( .CLK(n3710), .C(n3711) );
  CKBD0 U3594 ( .CLK(n3711), .C(n3712) );
  CKBD0 U3595 ( .CLK(n3712), .C(n3713) );
  CKBD0 U3596 ( .CLK(n3713), .C(n3714) );
  CKBD0 U3597 ( .CLK(n3714), .C(n3715) );
  CKBD0 U3598 ( .CLK(n3715), .C(n3716) );
  CKBD0 U3599 ( .CLK(n3716), .C(n3717) );
  CKBD0 U3600 ( .CLK(n3717), .C(n3718) );
  CKBD0 U3601 ( .CLK(n3718), .C(n3719) );
  CKBD0 U3602 ( .CLK(n3719), .C(n3720) );
  BUFFD0 U3603 ( .I(n3720), .Z(n3721) );
  CKBD0 U3604 ( .CLK(n3721), .C(n3722) );
  CKBD0 U3605 ( .CLK(n3722), .C(n3723) );
  CKBD0 U3606 ( .CLK(n3723), .C(n3724) );
  CKBD0 U3607 ( .CLK(n3724), .C(n3725) );
  CKBD0 U3608 ( .CLK(n3725), .C(n3726) );
  CKBD0 U3609 ( .CLK(n3726), .C(n3727) );
  CKBD0 U3610 ( .CLK(n3727), .C(n3728) );
  CKBD0 U3611 ( .CLK(n3728), .C(n3729) );
  CKBD0 U3612 ( .CLK(n3729), .C(n3730) );
  CKBD0 U3613 ( .CLK(n3730), .C(n3731) );
  BUFFD0 U3614 ( .I(n3731), .Z(n3732) );
  CKBD0 U3615 ( .CLK(n3732), .C(n3733) );
  CKBD0 U3616 ( .CLK(n3733), .C(n3734) );
  CKBD0 U3617 ( .CLK(n3734), .C(n3735) );
  CKBD0 U3618 ( .CLK(n3735), .C(n3736) );
  CKBD0 U3619 ( .CLK(n3736), .C(n3737) );
  CKBD0 U3620 ( .CLK(n3737), .C(n3738) );
  CKBD0 U3621 ( .CLK(n3738), .C(n3739) );
  CKBD0 U3622 ( .CLK(n3739), .C(n3740) );
  CKBD0 U3623 ( .CLK(n3740), .C(n3741) );
  BUFFD0 U3624 ( .I(n3741), .Z(n3742) );
  CKBD0 U3625 ( .CLK(n3742), .C(n3743) );
  CKBD0 U3626 ( .CLK(n3743), .C(n3744) );
  CKBD0 U3627 ( .CLK(n3744), .C(n3745) );
  CKBD0 U3628 ( .CLK(n3745), .C(n3746) );
  CKBD0 U3629 ( .CLK(n3746), .C(n3747) );
  CKBD0 U3630 ( .CLK(n3747), .C(n3748) );
  CKBD0 U3631 ( .CLK(n3748), .C(n3749) );
  CKBD0 U3632 ( .CLK(n3749), .C(n3750) );
  CKBD0 U3633 ( .CLK(n3750), .C(n3751) );
  CKBD0 U3634 ( .CLK(n3751), .C(n3752) );
  CKBD0 U3635 ( .CLK(n3752), .C(n3753) );
  BUFFD0 U3636 ( .I(n3753), .Z(n3754) );
  CKBD0 U3637 ( .CLK(n3754), .C(n3755) );
  CKBD0 U3638 ( .CLK(n3755), .C(n3756) );
  CKBD0 U3639 ( .CLK(n3756), .C(n3757) );
  CKBD0 U3640 ( .CLK(n3757), .C(n3758) );
  CKBD0 U3641 ( .CLK(n3758), .C(n3759) );
  CKBD0 U3642 ( .CLK(n3759), .C(n3760) );
  CKBD0 U3643 ( .CLK(n3760), .C(n3761) );
  CKBD0 U3644 ( .CLK(n3761), .C(n3762) );
  CKBD0 U3645 ( .CLK(n3762), .C(n3763) );
  BUFFD0 U3646 ( .I(n3763), .Z(n3764) );
  CKBD0 U3647 ( .CLK(n3764), .C(n3765) );
  CKBD0 U3648 ( .CLK(n3765), .C(n3766) );
  CKBD0 U3649 ( .CLK(n3766), .C(n3767) );
  CKBD0 U3650 ( .CLK(n3767), .C(n3768) );
  CKBD0 U3651 ( .CLK(n3768), .C(n3769) );
  CKBD0 U3652 ( .CLK(n3769), .C(n3770) );
  CKBD0 U3653 ( .CLK(n3770), .C(n3771) );
  CKBD0 U3654 ( .CLK(n3771), .C(n3772) );
  CKBD0 U3655 ( .CLK(n3772), .C(n3773) );
  CKBD0 U3656 ( .CLK(n3773), .C(n3774) );
  BUFFD0 U3657 ( .I(n3774), .Z(n3775) );
  CKBD0 U3658 ( .CLK(n3775), .C(n3776) );
  CKBD0 U3659 ( .CLK(n3776), .C(n3777) );
  CKBD0 U3660 ( .CLK(n3777), .C(n3778) );
  CKBD0 U3661 ( .CLK(n3778), .C(n3779) );
  CKBD0 U3662 ( .CLK(n3779), .C(n3780) );
  CKBD0 U3663 ( .CLK(n3780), .C(n3781) );
  CKBD0 U3664 ( .CLK(n3781), .C(n3782) );
  CKBD0 U3665 ( .CLK(n3782), .C(n3783) );
  CKBD0 U3666 ( .CLK(n3783), .C(n3784) );
  CKBD0 U3667 ( .CLK(n3784), .C(n3785) );
  BUFFD0 U3668 ( .I(n3785), .Z(n3786) );
  CKBD0 U3669 ( .CLK(n3786), .C(n3787) );
  CKBD0 U3670 ( .CLK(n3787), .C(n3788) );
  CKBD0 U3671 ( .CLK(n3788), .C(n3789) );
  CKBD0 U3672 ( .CLK(n3789), .C(n3790) );
  CKBD0 U3673 ( .CLK(n3790), .C(n3791) );
  CKBD0 U3674 ( .CLK(n3791), .C(n3792) );
  CKBD0 U3675 ( .CLK(n3792), .C(n3793) );
  CKBD0 U3676 ( .CLK(n3793), .C(n3794) );
  CKBD0 U3677 ( .CLK(n3794), .C(n3795) );
  CKBD0 U3678 ( .CLK(n3795), .C(n3796) );
  BUFFD0 U3679 ( .I(n3796), .Z(n3797) );
  CKBD0 U3680 ( .CLK(n3797), .C(n3798) );
  CKBD0 U3681 ( .CLK(n3798), .C(n3799) );
  CKBD0 U3682 ( .CLK(n3799), .C(n3800) );
  CKBD0 U3683 ( .CLK(n3800), .C(n3801) );
  CKBD0 U3684 ( .CLK(n3801), .C(n3802) );
  CKBD0 U3685 ( .CLK(n3802), .C(n3803) );
  CKBD0 U3686 ( .CLK(n3803), .C(n3804) );
  CKBD0 U3687 ( .CLK(n3804), .C(n3805) );
  CKBD0 U3688 ( .CLK(n3805), .C(n3806) );
  CKBD0 U3689 ( .CLK(n3806), .C(n3807) );
  BUFFD0 U3690 ( .I(n3807), .Z(n3808) );
  CKBD0 U3691 ( .CLK(n3808), .C(n3809) );
  CKBD0 U3692 ( .CLK(n3809), .C(n3810) );
  CKBD0 U3693 ( .CLK(n3810), .C(n3811) );
  CKBD0 U3694 ( .CLK(n3811), .C(n3812) );
  CKBD0 U3695 ( .CLK(n3812), .C(n3813) );
  BUFFD0 U3696 ( .I(n3813), .Z(n3814) );
  CKBD0 U3697 ( .CLK(n3814), .C(n3815) );
  BUFFD0 U3698 ( .I(n3815), .Z(n3816) );
  CKBD0 U3699 ( .CLK(n3816), .C(n3817) );
  BUFFD0 U3700 ( .I(n3817), .Z(n3818) );
  CKBD0 U3701 ( .CLK(n3818), .C(n3819) );
  BUFFD0 U3702 ( .I(n3819), .Z(n3820) );
  CKBD0 U3703 ( .CLK(n3820), .C(n3821) );
  BUFFD0 U3704 ( .I(n3821), .Z(n3822) );
  CKBD0 U3705 ( .CLK(n3822), .C(n3823) );
  BUFFD0 U3706 ( .I(n3823), .Z(n3824) );
  CKBD0 U3707 ( .CLK(n3824), .C(n3825) );
  BUFFD0 U3708 ( .I(n3825), .Z(n3826) );
  CKBD0 U3709 ( .CLK(n3826), .C(n3827) );
  BUFFD0 U3710 ( .I(n3827), .Z(n3828) );
  BUFFD0 U3711 ( .I(n3830), .Z(n3829) );
  BUFFD0 U3712 ( .I(n3831), .Z(n3830) );
  BUFFD0 U3713 ( .I(n9177), .Z(n3831) );
  CKBD0 U3714 ( .CLK(n1277), .C(n3832) );
  CKBD0 U3715 ( .CLK(n3832), .C(n3833) );
  CKBD0 U3716 ( .CLK(n3833), .C(n3834) );
  BUFFD0 U3717 ( .I(n3834), .Z(n3835) );
  CKBD0 U3718 ( .CLK(n3835), .C(n3836) );
  CKBD0 U3719 ( .CLK(n3836), .C(n3837) );
  CKBD0 U3720 ( .CLK(n3837), .C(n3838) );
  CKBD0 U3721 ( .CLK(n3838), .C(n3839) );
  CKBD0 U3722 ( .CLK(n3839), .C(n3840) );
  CKBD0 U3723 ( .CLK(n3840), .C(n3841) );
  CKBD0 U3724 ( .CLK(n3841), .C(n3842) );
  CKBD0 U3725 ( .CLK(n3842), .C(n3843) );
  CKBD0 U3726 ( .CLK(n3843), .C(n3844) );
  CKBD0 U3727 ( .CLK(n3844), .C(n3845) );
  BUFFD0 U3728 ( .I(n3845), .Z(n3846) );
  CKBD0 U3729 ( .CLK(n3846), .C(n3847) );
  CKBD0 U3730 ( .CLK(n3847), .C(n3848) );
  CKBD0 U3731 ( .CLK(n3848), .C(n3849) );
  CKBD0 U3732 ( .CLK(n3849), .C(n3850) );
  CKBD0 U3733 ( .CLK(n3850), .C(n3851) );
  CKBD0 U3734 ( .CLK(n3851), .C(n3852) );
  CKBD0 U3735 ( .CLK(n3852), .C(n3853) );
  CKBD0 U3736 ( .CLK(n3853), .C(n3854) );
  CKBD0 U3737 ( .CLK(n3854), .C(n3855) );
  CKBD0 U3738 ( .CLK(n3855), .C(n3856) );
  BUFFD0 U3739 ( .I(n3856), .Z(n3857) );
  CKBD0 U3740 ( .CLK(n3857), .C(n3858) );
  CKBD0 U3741 ( .CLK(n3858), .C(n3859) );
  CKBD0 U3742 ( .CLK(n3859), .C(n3860) );
  CKBD0 U3743 ( .CLK(n3860), .C(n3861) );
  CKBD0 U3744 ( .CLK(n3861), .C(n3862) );
  CKBD0 U3745 ( .CLK(n3862), .C(n3863) );
  CKBD0 U3746 ( .CLK(n3863), .C(n3864) );
  CKBD0 U3747 ( .CLK(n3864), .C(n3865) );
  CKBD0 U3748 ( .CLK(n3865), .C(n3866) );
  CKBD0 U3749 ( .CLK(n3866), .C(n3867) );
  BUFFD0 U3750 ( .I(n3867), .Z(n3868) );
  CKBD0 U3751 ( .CLK(n3868), .C(n3869) );
  CKBD0 U3752 ( .CLK(n3869), .C(n3870) );
  CKBD0 U3753 ( .CLK(n3870), .C(n3871) );
  CKBD0 U3754 ( .CLK(n3871), .C(n3872) );
  CKBD0 U3755 ( .CLK(n3872), .C(n3873) );
  CKBD0 U3756 ( .CLK(n3873), .C(n3874) );
  CKBD0 U3757 ( .CLK(n3874), .C(n3875) );
  CKBD0 U3758 ( .CLK(n3875), .C(n3876) );
  CKBD0 U3759 ( .CLK(n3876), .C(n3877) );
  CKBD0 U3760 ( .CLK(n3877), .C(n3878) );
  BUFFD0 U3761 ( .I(n3878), .Z(n3879) );
  CKBD0 U3762 ( .CLK(n3879), .C(n3880) );
  CKBD0 U3763 ( .CLK(n3880), .C(n3881) );
  CKBD0 U3764 ( .CLK(n3881), .C(n3882) );
  CKBD0 U3765 ( .CLK(n3882), .C(n3883) );
  CKBD0 U3766 ( .CLK(n3883), .C(n3884) );
  CKBD0 U3767 ( .CLK(n3884), .C(n3885) );
  CKBD0 U3768 ( .CLK(n3885), .C(n3886) );
  CKBD0 U3769 ( .CLK(n3886), .C(n3887) );
  CKBD0 U3770 ( .CLK(n3887), .C(n3888) );
  CKBD0 U3771 ( .CLK(n3888), .C(n3889) );
  BUFFD0 U3772 ( .I(n3889), .Z(n3890) );
  CKBD0 U3773 ( .CLK(n3890), .C(n3891) );
  CKBD0 U3774 ( .CLK(n3891), .C(n3892) );
  CKBD0 U3775 ( .CLK(n3892), .C(n3893) );
  CKBD0 U3776 ( .CLK(n3893), .C(n3894) );
  CKBD0 U3777 ( .CLK(n3894), .C(n3895) );
  CKBD0 U3778 ( .CLK(n3895), .C(n3896) );
  CKBD0 U3779 ( .CLK(n3896), .C(n3897) );
  CKBD0 U3780 ( .CLK(n3897), .C(n3898) );
  CKBD0 U3781 ( .CLK(n3898), .C(n3899) );
  BUFFD0 U3782 ( .I(n3899), .Z(n3900) );
  CKBD0 U3783 ( .CLK(n3900), .C(n3901) );
  CKBD0 U3784 ( .CLK(n3901), .C(n3902) );
  CKBD0 U3785 ( .CLK(n3902), .C(n3903) );
  CKBD0 U3786 ( .CLK(n3903), .C(n3904) );
  CKBD0 U3787 ( .CLK(n3904), .C(n3905) );
  CKBD0 U3788 ( .CLK(n3905), .C(n3906) );
  CKBD0 U3789 ( .CLK(n3906), .C(n3907) );
  CKBD0 U3790 ( .CLK(n3907), .C(n3908) );
  CKBD0 U3791 ( .CLK(n3908), .C(n3909) );
  CKBD0 U3792 ( .CLK(n3909), .C(n3910) );
  CKBD0 U3793 ( .CLK(n3910), .C(n3911) );
  BUFFD0 U3794 ( .I(n3911), .Z(n3912) );
  CKBD0 U3795 ( .CLK(n3912), .C(n3913) );
  CKBD0 U3796 ( .CLK(n3913), .C(n3914) );
  CKBD0 U3797 ( .CLK(n3914), .C(n3915) );
  CKBD0 U3798 ( .CLK(n3915), .C(n3916) );
  CKBD0 U3799 ( .CLK(n3916), .C(n3917) );
  CKBD0 U3800 ( .CLK(n3917), .C(n3918) );
  CKBD0 U3801 ( .CLK(n3918), .C(n3919) );
  CKBD0 U3802 ( .CLK(n3919), .C(n3920) );
  CKBD0 U3803 ( .CLK(n3920), .C(n3921) );
  BUFFD0 U3804 ( .I(n3921), .Z(n3922) );
  CKBD0 U3805 ( .CLK(n3922), .C(n3923) );
  CKBD0 U3806 ( .CLK(n3923), .C(n3924) );
  CKBD0 U3807 ( .CLK(n3924), .C(n3925) );
  CKBD0 U3808 ( .CLK(n3925), .C(n3926) );
  CKBD0 U3809 ( .CLK(n3926), .C(n3927) );
  CKBD0 U3810 ( .CLK(n3927), .C(n3928) );
  CKBD0 U3811 ( .CLK(n3928), .C(n3929) );
  CKBD0 U3812 ( .CLK(n3929), .C(n3930) );
  CKBD0 U3813 ( .CLK(n3930), .C(n3931) );
  BUFFD0 U3814 ( .I(n3931), .Z(n3932) );
  CKBD0 U3815 ( .CLK(n3932), .C(n3933) );
  CKBD0 U3816 ( .CLK(n3933), .C(n3934) );
  CKBD0 U3817 ( .CLK(n3934), .C(n3935) );
  CKBD0 U3818 ( .CLK(n3935), .C(n3936) );
  CKBD0 U3819 ( .CLK(n3936), .C(n3937) );
  CKBD0 U3820 ( .CLK(n3937), .C(n3938) );
  CKBD0 U3821 ( .CLK(n3938), .C(n3939) );
  CKBD0 U3822 ( .CLK(n3939), .C(n3940) );
  CKBD0 U3823 ( .CLK(n3940), .C(n3941) );
  CKBD0 U3824 ( .CLK(n3941), .C(n3942) );
  CKBD0 U3825 ( .CLK(n3942), .C(n3943) );
  BUFFD0 U3826 ( .I(n3943), .Z(n3944) );
  CKBD0 U3827 ( .CLK(n3944), .C(n3945) );
  CKBD0 U3828 ( .CLK(n3945), .C(n3946) );
  CKBD0 U3829 ( .CLK(n3946), .C(n3947) );
  CKBD0 U3830 ( .CLK(n3947), .C(n3948) );
  CKBD0 U3831 ( .CLK(n3948), .C(n3949) );
  BUFFD0 U3832 ( .I(n3949), .Z(n3950) );
  CKBD0 U3833 ( .CLK(n3950), .C(n3951) );
  BUFFD0 U3834 ( .I(n3951), .Z(n3952) );
  CKBD0 U3835 ( .CLK(n3952), .C(n3953) );
  BUFFD0 U3836 ( .I(n3953), .Z(n3954) );
  CKBD0 U3837 ( .CLK(n3954), .C(n3955) );
  BUFFD0 U3838 ( .I(n3955), .Z(n3956) );
  CKBD0 U3839 ( .CLK(n3956), .C(n3957) );
  BUFFD0 U3840 ( .I(n3957), .Z(n3958) );
  CKBD0 U3841 ( .CLK(n3958), .C(n3959) );
  BUFFD0 U3842 ( .I(n3959), .Z(n3960) );
  CKBD0 U3843 ( .CLK(n3960), .C(n3961) );
  BUFFD0 U3844 ( .I(n3961), .Z(n3962) );
  CKBD0 U3845 ( .CLK(n3962), .C(n3963) );
  BUFFD0 U3846 ( .I(n3963), .Z(n3964) );
  BUFFD0 U3847 ( .I(n3966), .Z(n3965) );
  BUFFD0 U3848 ( .I(n3967), .Z(n3966) );
  BUFFD0 U3849 ( .I(n9178), .Z(n3967) );
  CKBD0 U3850 ( .CLK(n1275), .C(n3968) );
  CKBD0 U3851 ( .CLK(n3968), .C(n3969) );
  CKBD0 U3852 ( .CLK(n3969), .C(n3970) );
  BUFFD0 U3853 ( .I(n3970), .Z(n3971) );
  CKBD0 U3854 ( .CLK(n3971), .C(n3972) );
  CKBD0 U3855 ( .CLK(n3972), .C(n3973) );
  CKBD0 U3856 ( .CLK(n3973), .C(n3974) );
  CKBD0 U3857 ( .CLK(n3974), .C(n3975) );
  CKBD0 U3858 ( .CLK(n3975), .C(n3976) );
  CKBD0 U3859 ( .CLK(n3976), .C(n3977) );
  CKBD0 U3860 ( .CLK(n3977), .C(n3978) );
  CKBD0 U3861 ( .CLK(n3978), .C(n3979) );
  CKBD0 U3862 ( .CLK(n3979), .C(n3980) );
  CKBD0 U3863 ( .CLK(n3980), .C(n3981) );
  CKBD0 U3864 ( .CLK(n3981), .C(n3982) );
  BUFFD0 U3865 ( .I(n3982), .Z(n3983) );
  CKBD0 U3866 ( .CLK(n3983), .C(n3984) );
  CKBD0 U3867 ( .CLK(n3984), .C(n3985) );
  CKBD0 U3868 ( .CLK(n3985), .C(n3986) );
  CKBD0 U3869 ( .CLK(n3986), .C(n3987) );
  CKBD0 U3870 ( .CLK(n3987), .C(n3988) );
  CKBD0 U3871 ( .CLK(n3988), .C(n3989) );
  CKBD0 U3872 ( .CLK(n3989), .C(n3990) );
  CKBD0 U3873 ( .CLK(n3990), .C(n3991) );
  CKBD0 U3874 ( .CLK(n3991), .C(n3992) );
  BUFFD0 U3875 ( .I(n3992), .Z(n3993) );
  CKBD0 U3876 ( .CLK(n3993), .C(n3994) );
  CKBD0 U3877 ( .CLK(n3994), .C(n3995) );
  CKBD0 U3878 ( .CLK(n3995), .C(n3996) );
  CKBD0 U3879 ( .CLK(n3996), .C(n3997) );
  CKBD0 U3880 ( .CLK(n3997), .C(n3998) );
  CKBD0 U3881 ( .CLK(n3998), .C(n3999) );
  CKBD0 U3882 ( .CLK(n3999), .C(n4000) );
  CKBD0 U3883 ( .CLK(n4000), .C(n4001) );
  CKBD0 U3884 ( .CLK(n4001), .C(n4002) );
  BUFFD0 U3885 ( .I(n4002), .Z(n4003) );
  CKBD0 U3886 ( .CLK(n4003), .C(n4004) );
  CKBD0 U3887 ( .CLK(n4004), .C(n4005) );
  CKBD0 U3888 ( .CLK(n4005), .C(n4006) );
  CKBD0 U3889 ( .CLK(n4006), .C(n4007) );
  CKBD0 U3890 ( .CLK(n4007), .C(n4008) );
  CKBD0 U3891 ( .CLK(n4008), .C(n4009) );
  CKBD0 U3892 ( .CLK(n4009), .C(n4010) );
  CKBD0 U3893 ( .CLK(n4010), .C(n4011) );
  CKBD0 U3894 ( .CLK(n4011), .C(n4012) );
  CKBD0 U3895 ( .CLK(n4012), .C(n4013) );
  CKBD0 U3896 ( .CLK(n4013), .C(n4014) );
  BUFFD0 U3897 ( .I(n4014), .Z(n4015) );
  CKBD0 U3898 ( .CLK(n4015), .C(n4016) );
  CKBD0 U3899 ( .CLK(n4016), .C(n4017) );
  CKBD0 U3900 ( .CLK(n4017), .C(n4018) );
  CKBD0 U3901 ( .CLK(n4018), .C(n4019) );
  CKBD0 U3902 ( .CLK(n4019), .C(n4020) );
  CKBD0 U3903 ( .CLK(n4020), .C(n4021) );
  CKBD0 U3904 ( .CLK(n4021), .C(n4022) );
  CKBD0 U3905 ( .CLK(n4022), .C(n4023) );
  CKBD0 U3906 ( .CLK(n4023), .C(n4024) );
  BUFFD0 U3907 ( .I(n4024), .Z(n4025) );
  CKBD0 U3908 ( .CLK(n4025), .C(n4026) );
  CKBD0 U3909 ( .CLK(n4026), .C(n4027) );
  CKBD0 U3910 ( .CLK(n4027), .C(n4028) );
  CKBD0 U3911 ( .CLK(n4028), .C(n4029) );
  CKBD0 U3912 ( .CLK(n4029), .C(n4030) );
  CKBD0 U3913 ( .CLK(n4030), .C(n4031) );
  CKBD0 U3914 ( .CLK(n4031), .C(n4032) );
  CKBD0 U3915 ( .CLK(n4032), .C(n4033) );
  CKBD0 U3916 ( .CLK(n4033), .C(n4034) );
  CKBD0 U3917 ( .CLK(n4034), .C(n4035) );
  BUFFD0 U3918 ( .I(n4035), .Z(n4036) );
  CKBD0 U3919 ( .CLK(n4036), .C(n4037) );
  CKBD0 U3920 ( .CLK(n4037), .C(n4038) );
  CKBD0 U3921 ( .CLK(n4038), .C(n4039) );
  CKBD0 U3922 ( .CLK(n4039), .C(n4040) );
  CKBD0 U3923 ( .CLK(n4040), .C(n4041) );
  CKBD0 U3924 ( .CLK(n4041), .C(n4042) );
  CKBD0 U3925 ( .CLK(n4042), .C(n4043) );
  CKBD0 U3926 ( .CLK(n4043), .C(n4044) );
  CKBD0 U3927 ( .CLK(n4044), .C(n4045) );
  CKBD0 U3928 ( .CLK(n4045), .C(n4046) );
  CKBD0 U3929 ( .CLK(n4046), .C(n4047) );
  BUFFD0 U3930 ( .I(n4047), .Z(n4048) );
  CKBD0 U3931 ( .CLK(n4048), .C(n4049) );
  CKBD0 U3932 ( .CLK(n4049), .C(n4050) );
  CKBD0 U3933 ( .CLK(n4050), .C(n4051) );
  CKBD0 U3934 ( .CLK(n4051), .C(n4052) );
  CKBD0 U3935 ( .CLK(n4052), .C(n4053) );
  CKBD0 U3936 ( .CLK(n4053), .C(n4054) );
  CKBD0 U3937 ( .CLK(n4054), .C(n4055) );
  CKBD0 U3938 ( .CLK(n4055), .C(n4056) );
  CKBD0 U3939 ( .CLK(n4056), .C(n4057) );
  BUFFD0 U3940 ( .I(n4057), .Z(n4058) );
  CKBD0 U3941 ( .CLK(n4058), .C(n4059) );
  CKBD0 U3942 ( .CLK(n4059), .C(n4060) );
  CKBD0 U3943 ( .CLK(n4060), .C(n4061) );
  CKBD0 U3944 ( .CLK(n4061), .C(n4062) );
  CKBD0 U3945 ( .CLK(n4062), .C(n4063) );
  CKBD0 U3946 ( .CLK(n4063), .C(n4064) );
  CKBD0 U3947 ( .CLK(n4064), .C(n4065) );
  CKBD0 U3948 ( .CLK(n4065), .C(n4066) );
  CKBD0 U3949 ( .CLK(n4066), .C(n4067) );
  BUFFD0 U3950 ( .I(n4067), .Z(n4068) );
  CKBD0 U3951 ( .CLK(n4068), .C(n4069) );
  CKBD0 U3952 ( .CLK(n4069), .C(n4070) );
  CKBD0 U3953 ( .CLK(n4070), .C(n4071) );
  CKBD0 U3954 ( .CLK(n4071), .C(n4072) );
  CKBD0 U3955 ( .CLK(n4072), .C(n4073) );
  CKBD0 U3956 ( .CLK(n4073), .C(n4074) );
  CKBD0 U3957 ( .CLK(n4074), .C(n4075) );
  CKBD0 U3958 ( .CLK(n4075), .C(n4076) );
  CKBD0 U3959 ( .CLK(n4076), .C(n4077) );
  CKBD0 U3960 ( .CLK(n4077), .C(n4078) );
  CKBD0 U3961 ( .CLK(n4078), .C(n4079) );
  BUFFD0 U3962 ( .I(n4079), .Z(n4080) );
  CKBD0 U3963 ( .CLK(n4080), .C(n4081) );
  CKBD0 U3964 ( .CLK(n4081), .C(n4082) );
  CKBD0 U3965 ( .CLK(n4082), .C(n4083) );
  CKBD0 U3966 ( .CLK(n4083), .C(n4084) );
  CKBD0 U3967 ( .CLK(n4084), .C(n4085) );
  BUFFD0 U3968 ( .I(n4085), .Z(n4086) );
  CKBD0 U3969 ( .CLK(n4086), .C(n4087) );
  BUFFD0 U3970 ( .I(n4087), .Z(n4088) );
  CKBD0 U3971 ( .CLK(n4088), .C(n4089) );
  BUFFD0 U3972 ( .I(n4089), .Z(n4090) );
  CKBD0 U3973 ( .CLK(n4090), .C(n4091) );
  BUFFD0 U3974 ( .I(n4091), .Z(n4092) );
  CKBD0 U3975 ( .CLK(n4092), .C(n4093) );
  BUFFD0 U3976 ( .I(n4093), .Z(n4094) );
  CKBD0 U3977 ( .CLK(n4094), .C(n4095) );
  BUFFD0 U3978 ( .I(n4095), .Z(n4096) );
  CKBD0 U3979 ( .CLK(n4096), .C(n4097) );
  BUFFD0 U3980 ( .I(n4097), .Z(n4098) );
  CKBD0 U3981 ( .CLK(n4098), .C(n4099) );
  BUFFD0 U3982 ( .I(n4099), .Z(n4100) );
  BUFFD0 U3983 ( .I(n4102), .Z(n4101) );
  BUFFD0 U3984 ( .I(n4103), .Z(n4102) );
  BUFFD0 U3985 ( .I(n9179), .Z(n4103) );
  CKBD0 U3986 ( .CLK(n1273), .C(n4104) );
  CKBD0 U3987 ( .CLK(n4104), .C(n4105) );
  CKBD0 U3988 ( .CLK(n4105), .C(n4106) );
  BUFFD0 U3989 ( .I(n4106), .Z(n4107) );
  CKBD0 U3990 ( .CLK(n4107), .C(n4108) );
  CKBD0 U3991 ( .CLK(n4108), .C(n4109) );
  CKBD0 U3992 ( .CLK(n4109), .C(n4110) );
  CKBD0 U3993 ( .CLK(n4110), .C(n4111) );
  CKBD0 U3994 ( .CLK(n4111), .C(n4112) );
  CKBD0 U3995 ( .CLK(n4112), .C(n4113) );
  CKBD0 U3996 ( .CLK(n4113), .C(n4114) );
  CKBD0 U3997 ( .CLK(n4114), .C(n4115) );
  CKBD0 U3998 ( .CLK(n4115), .C(n4116) );
  CKBD0 U3999 ( .CLK(n4116), .C(n4117) );
  BUFFD0 U4000 ( .I(n4117), .Z(n4118) );
  CKBD0 U4001 ( .CLK(n4118), .C(n4119) );
  CKBD0 U4002 ( .CLK(n4119), .C(n4120) );
  CKBD0 U4003 ( .CLK(n4120), .C(n4121) );
  CKBD0 U4004 ( .CLK(n4121), .C(n4122) );
  CKBD0 U4005 ( .CLK(n4122), .C(n4123) );
  CKBD0 U4006 ( .CLK(n4123), .C(n4124) );
  CKBD0 U4007 ( .CLK(n4124), .C(n4125) );
  CKBD0 U4008 ( .CLK(n4125), .C(n4126) );
  CKBD0 U4009 ( .CLK(n4126), .C(n4127) );
  CKBD0 U4010 ( .CLK(n4127), .C(n4128) );
  BUFFD0 U4011 ( .I(n4128), .Z(n4129) );
  CKBD0 U4012 ( .CLK(n4129), .C(n4130) );
  CKBD0 U4013 ( .CLK(n4130), .C(n4131) );
  CKBD0 U4014 ( .CLK(n4131), .C(n4132) );
  CKBD0 U4015 ( .CLK(n4132), .C(n4133) );
  CKBD0 U4016 ( .CLK(n4133), .C(n4134) );
  CKBD0 U4017 ( .CLK(n4134), .C(n4135) );
  CKBD0 U4018 ( .CLK(n4135), .C(n4136) );
  CKBD0 U4019 ( .CLK(n4136), .C(n4137) );
  CKBD0 U4020 ( .CLK(n4137), .C(n4138) );
  BUFFD0 U4021 ( .I(n4138), .Z(n4139) );
  CKBD0 U4022 ( .CLK(n4139), .C(n4140) );
  CKBD0 U4023 ( .CLK(n4140), .C(n4141) );
  CKBD0 U4024 ( .CLK(n4141), .C(n4142) );
  CKBD0 U4025 ( .CLK(n4142), .C(n4143) );
  CKBD0 U4026 ( .CLK(n4143), .C(n4144) );
  CKBD0 U4027 ( .CLK(n4144), .C(n4145) );
  CKBD0 U4028 ( .CLK(n4145), .C(n4146) );
  CKBD0 U4029 ( .CLK(n4146), .C(n4147) );
  CKBD0 U4030 ( .CLK(n4147), .C(n4148) );
  CKBD0 U4031 ( .CLK(n4148), .C(n4149) );
  CKBD0 U4032 ( .CLK(n4149), .C(n4150) );
  BUFFD0 U4033 ( .I(n4150), .Z(n4151) );
  CKBD0 U4034 ( .CLK(n4151), .C(n4152) );
  CKBD0 U4035 ( .CLK(n4152), .C(n4153) );
  CKBD0 U4036 ( .CLK(n4153), .C(n4154) );
  CKBD0 U4037 ( .CLK(n4154), .C(n4155) );
  CKBD0 U4038 ( .CLK(n4155), .C(n4156) );
  CKBD0 U4039 ( .CLK(n4156), .C(n4157) );
  CKBD0 U4040 ( .CLK(n4157), .C(n4158) );
  CKBD0 U4041 ( .CLK(n4158), .C(n4159) );
  CKBD0 U4042 ( .CLK(n4159), .C(n4160) );
  BUFFD0 U4043 ( .I(n4160), .Z(n4161) );
  CKBD0 U4044 ( .CLK(n4161), .C(n4162) );
  CKBD0 U4045 ( .CLK(n4162), .C(n4163) );
  CKBD0 U4046 ( .CLK(n4163), .C(n4164) );
  CKBD0 U4047 ( .CLK(n4164), .C(n4165) );
  CKBD0 U4048 ( .CLK(n4165), .C(n4166) );
  CKBD0 U4049 ( .CLK(n4166), .C(n4167) );
  CKBD0 U4050 ( .CLK(n4167), .C(n4168) );
  CKBD0 U4051 ( .CLK(n4168), .C(n4169) );
  CKBD0 U4052 ( .CLK(n4169), .C(n4170) );
  CKBD0 U4053 ( .CLK(n4170), .C(n4171) );
  CKBD0 U4054 ( .CLK(n4171), .C(n4172) );
  BUFFD0 U4055 ( .I(n4172), .Z(n4173) );
  CKBD0 U4056 ( .CLK(n4173), .C(n4174) );
  CKBD0 U4057 ( .CLK(n4174), .C(n4175) );
  CKBD0 U4058 ( .CLK(n4175), .C(n4176) );
  CKBD0 U4059 ( .CLK(n4176), .C(n4177) );
  CKBD0 U4060 ( .CLK(n4177), .C(n4178) );
  CKBD0 U4061 ( .CLK(n4178), .C(n4179) );
  CKBD0 U4062 ( .CLK(n4179), .C(n4180) );
  CKBD0 U4063 ( .CLK(n4180), .C(n4181) );
  CKBD0 U4064 ( .CLK(n4181), .C(n4182) );
  BUFFD0 U4065 ( .I(n4182), .Z(n4183) );
  CKBD0 U4066 ( .CLK(n4183), .C(n4184) );
  CKBD0 U4067 ( .CLK(n4184), .C(n4185) );
  CKBD0 U4068 ( .CLK(n4185), .C(n4186) );
  CKBD0 U4069 ( .CLK(n4186), .C(n4187) );
  CKBD0 U4070 ( .CLK(n4187), .C(n4188) );
  CKBD0 U4071 ( .CLK(n4188), .C(n4189) );
  CKBD0 U4072 ( .CLK(n4189), .C(n4190) );
  CKBD0 U4073 ( .CLK(n4190), .C(n4191) );
  CKBD0 U4074 ( .CLK(n4191), .C(n4192) );
  CKBD0 U4075 ( .CLK(n4192), .C(n4193) );
  BUFFD0 U4076 ( .I(n4193), .Z(n4194) );
  CKBD0 U4077 ( .CLK(n4194), .C(n4195) );
  CKBD0 U4078 ( .CLK(n4195), .C(n4196) );
  CKBD0 U4079 ( .CLK(n4196), .C(n4197) );
  CKBD0 U4080 ( .CLK(n4197), .C(n4198) );
  CKBD0 U4081 ( .CLK(n4198), .C(n4199) );
  CKBD0 U4082 ( .CLK(n4199), .C(n4200) );
  CKBD0 U4083 ( .CLK(n4200), .C(n4201) );
  CKBD0 U4084 ( .CLK(n4201), .C(n4202) );
  CKBD0 U4085 ( .CLK(n4202), .C(n4203) );
  CKBD0 U4086 ( .CLK(n4203), .C(n4204) );
  BUFFD0 U4087 ( .I(n4204), .Z(n4205) );
  CKBD0 U4088 ( .CLK(n4205), .C(n4206) );
  CKBD0 U4089 ( .CLK(n4206), .C(n4207) );
  CKBD0 U4090 ( .CLK(n4207), .C(n4208) );
  CKBD0 U4091 ( .CLK(n4208), .C(n4209) );
  CKBD0 U4092 ( .CLK(n4209), .C(n4210) );
  CKBD0 U4093 ( .CLK(n4210), .C(n4211) );
  CKBD0 U4094 ( .CLK(n4211), .C(n4212) );
  CKBD0 U4095 ( .CLK(n4212), .C(n4213) );
  CKBD0 U4096 ( .CLK(n4213), .C(n4214) );
  CKBD0 U4097 ( .CLK(n4214), .C(n4215) );
  BUFFD0 U4098 ( .I(n4215), .Z(n4216) );
  CKBD0 U4099 ( .CLK(n4216), .C(n4217) );
  CKBD0 U4100 ( .CLK(n4217), .C(n4218) );
  CKBD0 U4101 ( .CLK(n4218), .C(n4219) );
  CKBD0 U4102 ( .CLK(n4219), .C(n4220) );
  CKBD0 U4103 ( .CLK(n4220), .C(n4221) );
  BUFFD0 U4104 ( .I(n4221), .Z(n4222) );
  CKBD0 U4105 ( .CLK(n4222), .C(n4223) );
  BUFFD0 U4106 ( .I(n4223), .Z(n4224) );
  CKBD0 U4107 ( .CLK(n4224), .C(n4225) );
  BUFFD0 U4108 ( .I(n4225), .Z(n4226) );
  CKBD0 U4109 ( .CLK(n4226), .C(n4227) );
  BUFFD0 U4110 ( .I(n4227), .Z(n4228) );
  CKBD0 U4111 ( .CLK(n4228), .C(n4229) );
  BUFFD0 U4112 ( .I(n4229), .Z(n4230) );
  CKBD0 U4113 ( .CLK(n4230), .C(n4231) );
  BUFFD0 U4114 ( .I(n4231), .Z(n4232) );
  CKBD0 U4115 ( .CLK(n4232), .C(n4233) );
  BUFFD0 U4116 ( .I(n4233), .Z(n4234) );
  CKBD0 U4117 ( .CLK(n4234), .C(n4235) );
  BUFFD0 U4118 ( .I(n4235), .Z(n4236) );
  BUFFD0 U4119 ( .I(n4238), .Z(n4237) );
  BUFFD0 U4120 ( .I(n4239), .Z(n4238) );
  BUFFD0 U4121 ( .I(n4240), .Z(n4239) );
  BUFFD0 U4122 ( .I(n9180), .Z(n4240) );
  CKBD0 U4123 ( .CLK(n1271), .C(n4241) );
  CKBD0 U4124 ( .CLK(n4241), .C(n4242) );
  CKBD0 U4125 ( .CLK(n4242), .C(n4243) );
  BUFFD0 U4126 ( .I(n4243), .Z(n4244) );
  CKBD0 U4127 ( .CLK(n4244), .C(n4245) );
  CKBD0 U4128 ( .CLK(n4245), .C(n4246) );
  CKBD0 U4129 ( .CLK(n4246), .C(n4247) );
  CKBD0 U4130 ( .CLK(n4247), .C(n4248) );
  CKBD0 U4131 ( .CLK(n4248), .C(n4249) );
  CKBD0 U4132 ( .CLK(n4249), .C(n4250) );
  CKBD0 U4133 ( .CLK(n4250), .C(n4251) );
  CKBD0 U4134 ( .CLK(n4251), .C(n4252) );
  CKBD0 U4135 ( .CLK(n4252), .C(n4253) );
  CKBD0 U4136 ( .CLK(n4253), .C(n4254) );
  BUFFD0 U4137 ( .I(n4254), .Z(n4255) );
  CKBD0 U4138 ( .CLK(n4255), .C(n4256) );
  CKBD0 U4139 ( .CLK(n4256), .C(n4257) );
  CKBD0 U4140 ( .CLK(n4257), .C(n4258) );
  CKBD0 U4141 ( .CLK(n4258), .C(n4259) );
  CKBD0 U4142 ( .CLK(n4259), .C(n4260) );
  CKBD0 U4143 ( .CLK(n4260), .C(n4261) );
  CKBD0 U4144 ( .CLK(n4261), .C(n4262) );
  CKBD0 U4145 ( .CLK(n4262), .C(n4263) );
  CKBD0 U4146 ( .CLK(n4263), .C(n4264) );
  CKBD0 U4147 ( .CLK(n4264), .C(n4265) );
  BUFFD0 U4148 ( .I(n4265), .Z(n4266) );
  CKBD0 U4149 ( .CLK(n4266), .C(n4267) );
  CKBD0 U4150 ( .CLK(n4267), .C(n4268) );
  CKBD0 U4151 ( .CLK(n4268), .C(n4269) );
  CKBD0 U4152 ( .CLK(n4269), .C(n4270) );
  CKBD0 U4153 ( .CLK(n4270), .C(n4271) );
  CKBD0 U4154 ( .CLK(n4271), .C(n4272) );
  CKBD0 U4155 ( .CLK(n4272), .C(n4273) );
  CKBD0 U4156 ( .CLK(n4273), .C(n4274) );
  CKBD0 U4157 ( .CLK(n4274), .C(n4275) );
  CKBD0 U4158 ( .CLK(n4275), .C(n4276) );
  BUFFD0 U4159 ( .I(n4276), .Z(n4277) );
  CKBD0 U4160 ( .CLK(n4277), .C(n4278) );
  CKBD0 U4161 ( .CLK(n4278), .C(n4279) );
  CKBD0 U4162 ( .CLK(n4279), .C(n4280) );
  CKBD0 U4163 ( .CLK(n4280), .C(n4281) );
  CKBD0 U4164 ( .CLK(n4281), .C(n4282) );
  CKBD0 U4165 ( .CLK(n4282), .C(n4283) );
  CKBD0 U4166 ( .CLK(n4283), .C(n4284) );
  CKBD0 U4167 ( .CLK(n4284), .C(n4285) );
  CKBD0 U4168 ( .CLK(n4285), .C(n4286) );
  BUFFD0 U4169 ( .I(n4286), .Z(n4287) );
  CKBD0 U4170 ( .CLK(n4287), .C(n4288) );
  CKBD0 U4171 ( .CLK(n4288), .C(n4289) );
  CKBD0 U4172 ( .CLK(n4289), .C(n4290) );
  CKBD0 U4173 ( .CLK(n4290), .C(n4291) );
  CKBD0 U4174 ( .CLK(n4291), .C(n4292) );
  CKBD0 U4175 ( .CLK(n4292), .C(n4293) );
  CKBD0 U4176 ( .CLK(n4293), .C(n4294) );
  CKBD0 U4177 ( .CLK(n4294), .C(n4295) );
  CKBD0 U4178 ( .CLK(n4295), .C(n4296) );
  CKBD0 U4179 ( .CLK(n4296), .C(n4297) );
  CKBD0 U4180 ( .CLK(n4297), .C(n4298) );
  BUFFD0 U4181 ( .I(n4298), .Z(n4299) );
  CKBD0 U4182 ( .CLK(n4299), .C(n4300) );
  CKBD0 U4183 ( .CLK(n4300), .C(n4301) );
  CKBD0 U4184 ( .CLK(n4301), .C(n4302) );
  CKBD0 U4185 ( .CLK(n4302), .C(n4303) );
  CKBD0 U4186 ( .CLK(n4303), .C(n4304) );
  CKBD0 U4187 ( .CLK(n4304), .C(n4305) );
  CKBD0 U4188 ( .CLK(n4305), .C(n4306) );
  CKBD0 U4189 ( .CLK(n4306), .C(n4307) );
  CKBD0 U4190 ( .CLK(n4307), .C(n4308) );
  BUFFD0 U4191 ( .I(n4308), .Z(n4309) );
  CKBD0 U4192 ( .CLK(n4309), .C(n4310) );
  CKBD0 U4193 ( .CLK(n4310), .C(n4311) );
  CKBD0 U4194 ( .CLK(n4311), .C(n4312) );
  CKBD0 U4195 ( .CLK(n4312), .C(n4313) );
  CKBD0 U4196 ( .CLK(n4313), .C(n4314) );
  CKBD0 U4197 ( .CLK(n4314), .C(n4315) );
  CKBD0 U4198 ( .CLK(n4315), .C(n4316) );
  CKBD0 U4199 ( .CLK(n4316), .C(n4317) );
  CKBD0 U4200 ( .CLK(n4317), .C(n4318) );
  CKBD0 U4201 ( .CLK(n4318), .C(n4319) );
  CKBD0 U4202 ( .CLK(n4319), .C(n4320) );
  BUFFD0 U4203 ( .I(n4320), .Z(n4321) );
  CKBD0 U4204 ( .CLK(n4321), .C(n4322) );
  CKBD0 U4205 ( .CLK(n4322), .C(n4323) );
  CKBD0 U4206 ( .CLK(n4323), .C(n4324) );
  CKBD0 U4207 ( .CLK(n4324), .C(n4325) );
  CKBD0 U4208 ( .CLK(n4325), .C(n4326) );
  CKBD0 U4209 ( .CLK(n4326), .C(n4327) );
  CKBD0 U4210 ( .CLK(n4327), .C(n4328) );
  CKBD0 U4211 ( .CLK(n4328), .C(n4329) );
  CKBD0 U4212 ( .CLK(n4329), .C(n4330) );
  BUFFD0 U4213 ( .I(n4330), .Z(n4331) );
  CKBD0 U4214 ( .CLK(n4331), .C(n4332) );
  CKBD0 U4215 ( .CLK(n4332), .C(n4333) );
  CKBD0 U4216 ( .CLK(n4333), .C(n4334) );
  CKBD0 U4217 ( .CLK(n4334), .C(n4335) );
  CKBD0 U4218 ( .CLK(n4335), .C(n4336) );
  CKBD0 U4219 ( .CLK(n4336), .C(n4337) );
  CKBD0 U4220 ( .CLK(n4337), .C(n4338) );
  CKBD0 U4221 ( .CLK(n4338), .C(n4339) );
  CKBD0 U4222 ( .CLK(n4339), .C(n4340) );
  CKBD0 U4223 ( .CLK(n4340), .C(n4341) );
  BUFFD0 U4224 ( .I(n4341), .Z(n4342) );
  CKBD0 U4225 ( .CLK(n4342), .C(n4343) );
  CKBD0 U4226 ( .CLK(n4343), .C(n4344) );
  CKBD0 U4227 ( .CLK(n4344), .C(n4345) );
  CKBD0 U4228 ( .CLK(n4345), .C(n4346) );
  CKBD0 U4229 ( .CLK(n4346), .C(n4347) );
  CKBD0 U4230 ( .CLK(n4347), .C(n4348) );
  CKBD0 U4231 ( .CLK(n4348), .C(n4349) );
  CKBD0 U4232 ( .CLK(n4349), .C(n4350) );
  CKBD0 U4233 ( .CLK(n4350), .C(n4351) );
  CKBD0 U4234 ( .CLK(n4351), .C(n4352) );
  BUFFD0 U4235 ( .I(n4352), .Z(n4353) );
  CKBD0 U4236 ( .CLK(n4353), .C(n4354) );
  CKBD0 U4237 ( .CLK(n4354), .C(n4355) );
  CKBD0 U4238 ( .CLK(n4355), .C(n4356) );
  CKBD0 U4239 ( .CLK(n4356), .C(n4357) );
  CKBD0 U4240 ( .CLK(n4357), .C(n4358) );
  BUFFD0 U4241 ( .I(n4358), .Z(n4359) );
  CKBD0 U4242 ( .CLK(n4359), .C(n4360) );
  BUFFD0 U4243 ( .I(n4360), .Z(n4361) );
  CKBD0 U4244 ( .CLK(n4361), .C(n4362) );
  BUFFD0 U4245 ( .I(n4362), .Z(n4363) );
  CKBD0 U4246 ( .CLK(n4363), .C(n4364) );
  BUFFD0 U4247 ( .I(n4364), .Z(n4365) );
  CKBD0 U4248 ( .CLK(n4365), .C(n4366) );
  BUFFD0 U4249 ( .I(n4366), .Z(n4367) );
  CKBD0 U4250 ( .CLK(n4367), .C(n4368) );
  BUFFD0 U4251 ( .I(n4368), .Z(n4369) );
  CKBD0 U4252 ( .CLK(n4369), .C(n4370) );
  BUFFD0 U4253 ( .I(n4370), .Z(n4371) );
  CKBD0 U4254 ( .CLK(n4371), .C(n4372) );
  BUFFD0 U4255 ( .I(n4372), .Z(n4373) );
  BUFFD0 U4256 ( .I(n4375), .Z(n4374) );
  BUFFD0 U4257 ( .I(n4376), .Z(n4375) );
  BUFFD0 U4258 ( .I(n9181), .Z(n4376) );
  CKBD0 U4259 ( .CLK(n1269), .C(n4377) );
  CKBD0 U4260 ( .CLK(n4377), .C(n4378) );
  CKBD0 U4261 ( .CLK(n4378), .C(n4379) );
  BUFFD0 U4262 ( .I(n4379), .Z(n4380) );
  CKBD0 U4263 ( .CLK(n4380), .C(n4381) );
  CKBD0 U4264 ( .CLK(n4381), .C(n4382) );
  CKBD0 U4265 ( .CLK(n4382), .C(n4383) );
  CKBD0 U4266 ( .CLK(n4383), .C(n4384) );
  CKBD0 U4267 ( .CLK(n4384), .C(n4385) );
  CKBD0 U4268 ( .CLK(n4385), .C(n4386) );
  CKBD0 U4269 ( .CLK(n4386), .C(n4387) );
  CKBD0 U4270 ( .CLK(n4387), .C(n4388) );
  CKBD0 U4271 ( .CLK(n4388), .C(n4389) );
  CKBD0 U4272 ( .CLK(n4389), .C(n4390) );
  CKBD0 U4273 ( .CLK(n4390), .C(n4391) );
  BUFFD0 U4274 ( .I(n4391), .Z(n4392) );
  CKBD0 U4275 ( .CLK(n4392), .C(n4393) );
  CKBD0 U4276 ( .CLK(n4393), .C(n4394) );
  CKBD0 U4277 ( .CLK(n4394), .C(n4395) );
  CKBD0 U4278 ( .CLK(n4395), .C(n4396) );
  CKBD0 U4279 ( .CLK(n4396), .C(n4397) );
  CKBD0 U4280 ( .CLK(n4397), .C(n4398) );
  CKBD0 U4281 ( .CLK(n4398), .C(n4399) );
  CKBD0 U4282 ( .CLK(n4399), .C(n4400) );
  CKBD0 U4283 ( .CLK(n4400), .C(n4401) );
  BUFFD0 U4284 ( .I(n4401), .Z(n4402) );
  CKBD0 U4285 ( .CLK(n4402), .C(n4403) );
  CKBD0 U4286 ( .CLK(n4403), .C(n4404) );
  CKBD0 U4287 ( .CLK(n4404), .C(n4405) );
  CKBD0 U4288 ( .CLK(n4405), .C(n4406) );
  CKBD0 U4289 ( .CLK(n4406), .C(n4407) );
  CKBD0 U4290 ( .CLK(n4407), .C(n4408) );
  CKBD0 U4291 ( .CLK(n4408), .C(n4409) );
  CKBD0 U4292 ( .CLK(n4409), .C(n4410) );
  CKBD0 U4293 ( .CLK(n4410), .C(n4411) );
  BUFFD0 U4294 ( .I(n4411), .Z(n4412) );
  CKBD0 U4295 ( .CLK(n4412), .C(n4413) );
  CKBD0 U4296 ( .CLK(n4413), .C(n4414) );
  CKBD0 U4297 ( .CLK(n4414), .C(n4415) );
  CKBD0 U4298 ( .CLK(n4415), .C(n4416) );
  CKBD0 U4299 ( .CLK(n4416), .C(n4417) );
  CKBD0 U4300 ( .CLK(n4417), .C(n4418) );
  CKBD0 U4301 ( .CLK(n4418), .C(n4419) );
  CKBD0 U4302 ( .CLK(n4419), .C(n4420) );
  CKBD0 U4303 ( .CLK(n4420), .C(n4421) );
  CKBD0 U4304 ( .CLK(n4421), .C(n4422) );
  CKBD0 U4305 ( .CLK(n4422), .C(n4423) );
  BUFFD0 U4306 ( .I(n4423), .Z(n4424) );
  CKBD0 U4307 ( .CLK(n4424), .C(n4425) );
  CKBD0 U4308 ( .CLK(n4425), .C(n4426) );
  CKBD0 U4309 ( .CLK(n4426), .C(n4427) );
  CKBD0 U4310 ( .CLK(n4427), .C(n4428) );
  CKBD0 U4311 ( .CLK(n4428), .C(n4429) );
  CKBD0 U4312 ( .CLK(n4429), .C(n4430) );
  CKBD0 U4313 ( .CLK(n4430), .C(n4431) );
  CKBD0 U4314 ( .CLK(n4431), .C(n4432) );
  CKBD0 U4315 ( .CLK(n4432), .C(n4433) );
  BUFFD0 U4316 ( .I(n4433), .Z(n4434) );
  CKBD0 U4317 ( .CLK(n4434), .C(n4435) );
  CKBD0 U4318 ( .CLK(n4435), .C(n4436) );
  CKBD0 U4319 ( .CLK(n4436), .C(n4437) );
  CKBD0 U4320 ( .CLK(n4437), .C(n4438) );
  CKBD0 U4321 ( .CLK(n4438), .C(n4439) );
  CKBD0 U4322 ( .CLK(n4439), .C(n4440) );
  CKBD0 U4323 ( .CLK(n4440), .C(n4441) );
  CKBD0 U4324 ( .CLK(n4441), .C(n4442) );
  CKBD0 U4325 ( .CLK(n4442), .C(n4443) );
  CKBD0 U4326 ( .CLK(n4443), .C(n4444) );
  BUFFD0 U4327 ( .I(n4444), .Z(n4445) );
  CKBD0 U4328 ( .CLK(n4445), .C(n4446) );
  CKBD0 U4329 ( .CLK(n4446), .C(n4447) );
  CKBD0 U4330 ( .CLK(n4447), .C(n4448) );
  CKBD0 U4331 ( .CLK(n4448), .C(n4449) );
  CKBD0 U4332 ( .CLK(n4449), .C(n4450) );
  CKBD0 U4333 ( .CLK(n4450), .C(n4451) );
  CKBD0 U4334 ( .CLK(n4451), .C(n4452) );
  CKBD0 U4335 ( .CLK(n4452), .C(n4453) );
  CKBD0 U4336 ( .CLK(n4453), .C(n4454) );
  CKBD0 U4337 ( .CLK(n4454), .C(n4455) );
  CKBD0 U4338 ( .CLK(n4455), .C(n4456) );
  BUFFD0 U4339 ( .I(n4456), .Z(n4457) );
  CKBD0 U4340 ( .CLK(n4457), .C(n4458) );
  CKBD0 U4341 ( .CLK(n4458), .C(n4459) );
  CKBD0 U4342 ( .CLK(n4459), .C(n4460) );
  CKBD0 U4343 ( .CLK(n4460), .C(n4461) );
  CKBD0 U4344 ( .CLK(n4461), .C(n4462) );
  CKBD0 U4345 ( .CLK(n4462), .C(n4463) );
  CKBD0 U4346 ( .CLK(n4463), .C(n4464) );
  CKBD0 U4347 ( .CLK(n4464), .C(n4465) );
  CKBD0 U4348 ( .CLK(n4465), .C(n4466) );
  BUFFD0 U4349 ( .I(n4466), .Z(n4467) );
  CKBD0 U4350 ( .CLK(n4467), .C(n4468) );
  CKBD0 U4351 ( .CLK(n4468), .C(n4469) );
  CKBD0 U4352 ( .CLK(n4469), .C(n4470) );
  CKBD0 U4353 ( .CLK(n4470), .C(n4471) );
  CKBD0 U4354 ( .CLK(n4471), .C(n4472) );
  CKBD0 U4355 ( .CLK(n4472), .C(n4473) );
  CKBD0 U4356 ( .CLK(n4473), .C(n4474) );
  CKBD0 U4357 ( .CLK(n4474), .C(n4475) );
  CKBD0 U4358 ( .CLK(n4475), .C(n4476) );
  BUFFD0 U4359 ( .I(n4476), .Z(n4477) );
  CKBD0 U4360 ( .CLK(n4477), .C(n4478) );
  CKBD0 U4361 ( .CLK(n4478), .C(n4479) );
  CKBD0 U4362 ( .CLK(n4479), .C(n4480) );
  CKBD0 U4363 ( .CLK(n4480), .C(n4481) );
  CKBD0 U4364 ( .CLK(n4481), .C(n4482) );
  CKBD0 U4365 ( .CLK(n4482), .C(n4483) );
  CKBD0 U4366 ( .CLK(n4483), .C(n4484) );
  CKBD0 U4367 ( .CLK(n4484), .C(n4485) );
  CKBD0 U4368 ( .CLK(n4485), .C(n4486) );
  CKBD0 U4369 ( .CLK(n4486), .C(n4487) );
  CKBD0 U4370 ( .CLK(n4487), .C(n4488) );
  BUFFD0 U4371 ( .I(n4488), .Z(n4489) );
  CKBD0 U4372 ( .CLK(n4489), .C(n4490) );
  CKBD0 U4373 ( .CLK(n4490), .C(n4491) );
  CKBD0 U4374 ( .CLK(n4491), .C(n4492) );
  CKBD0 U4375 ( .CLK(n4492), .C(n4493) );
  CKBD0 U4376 ( .CLK(n4493), .C(n4494) );
  BUFFD0 U4377 ( .I(n4494), .Z(n4495) );
  CKBD0 U4378 ( .CLK(n4495), .C(n4496) );
  BUFFD0 U4379 ( .I(n4496), .Z(n4497) );
  CKBD0 U4380 ( .CLK(n4497), .C(n4498) );
  BUFFD0 U4381 ( .I(n4498), .Z(n4499) );
  CKBD0 U4382 ( .CLK(n4499), .C(n4500) );
  BUFFD0 U4383 ( .I(n4500), .Z(n4501) );
  CKBD0 U4384 ( .CLK(n4501), .C(n4502) );
  BUFFD0 U4385 ( .I(n4502), .Z(n4503) );
  CKBD0 U4386 ( .CLK(n4503), .C(n4504) );
  BUFFD0 U4387 ( .I(n4504), .Z(n4505) );
  CKBD0 U4388 ( .CLK(n4505), .C(n4506) );
  BUFFD0 U4389 ( .I(n4506), .Z(n4507) );
  CKBD0 U4390 ( .CLK(n4507), .C(n4508) );
  BUFFD0 U4391 ( .I(n4508), .Z(n4509) );
  BUFFD0 U4392 ( .I(n4511), .Z(n4510) );
  BUFFD0 U4393 ( .I(n4512), .Z(n4511) );
  BUFFD0 U4394 ( .I(n9182), .Z(n4512) );
  CKBD0 U4395 ( .CLK(n1267), .C(n4513) );
  CKBD0 U4396 ( .CLK(n4513), .C(n4514) );
  CKBD0 U4397 ( .CLK(n4514), .C(n4515) );
  BUFFD0 U4398 ( .I(n4515), .Z(n4516) );
  CKBD0 U4399 ( .CLK(n4516), .C(n4517) );
  CKBD0 U4400 ( .CLK(n4517), .C(n4518) );
  CKBD0 U4401 ( .CLK(n4518), .C(n4519) );
  CKBD0 U4402 ( .CLK(n4519), .C(n4520) );
  CKBD0 U4403 ( .CLK(n4520), .C(n4521) );
  CKBD0 U4404 ( .CLK(n4521), .C(n4522) );
  CKBD0 U4405 ( .CLK(n4522), .C(n4523) );
  CKBD0 U4406 ( .CLK(n4523), .C(n4524) );
  CKBD0 U4407 ( .CLK(n4524), .C(n4525) );
  CKBD0 U4408 ( .CLK(n4525), .C(n4526) );
  BUFFD0 U4409 ( .I(n4526), .Z(n4527) );
  CKBD0 U4410 ( .CLK(n4527), .C(n4528) );
  CKBD0 U4411 ( .CLK(n4528), .C(n4529) );
  CKBD0 U4412 ( .CLK(n4529), .C(n4530) );
  CKBD0 U4413 ( .CLK(n4530), .C(n4531) );
  CKBD0 U4414 ( .CLK(n4531), .C(n4532) );
  CKBD0 U4415 ( .CLK(n4532), .C(n4533) );
  CKBD0 U4416 ( .CLK(n4533), .C(n4534) );
  CKBD0 U4417 ( .CLK(n4534), .C(n4535) );
  CKBD0 U4418 ( .CLK(n4535), .C(n4536) );
  CKBD0 U4419 ( .CLK(n4536), .C(n4537) );
  BUFFD0 U4420 ( .I(n4537), .Z(n4538) );
  CKBD0 U4421 ( .CLK(n4538), .C(n4539) );
  CKBD0 U4422 ( .CLK(n4539), .C(n4540) );
  CKBD0 U4423 ( .CLK(n4540), .C(n4541) );
  CKBD0 U4424 ( .CLK(n4541), .C(n4542) );
  CKBD0 U4425 ( .CLK(n4542), .C(n4543) );
  CKBD0 U4426 ( .CLK(n4543), .C(n4544) );
  CKBD0 U4427 ( .CLK(n4544), .C(n4545) );
  CKBD0 U4428 ( .CLK(n4545), .C(n4546) );
  CKBD0 U4429 ( .CLK(n4546), .C(n4547) );
  BUFFD0 U4430 ( .I(n4547), .Z(n4548) );
  CKBD0 U4431 ( .CLK(n4548), .C(n4549) );
  CKBD0 U4432 ( .CLK(n4549), .C(n4550) );
  CKBD0 U4433 ( .CLK(n4550), .C(n4551) );
  CKBD0 U4434 ( .CLK(n4551), .C(n4552) );
  CKBD0 U4435 ( .CLK(n4552), .C(n4553) );
  CKBD0 U4436 ( .CLK(n4553), .C(n4554) );
  CKBD0 U4437 ( .CLK(n4554), .C(n4555) );
  CKBD0 U4438 ( .CLK(n4555), .C(n4556) );
  CKBD0 U4439 ( .CLK(n4556), .C(n4557) );
  CKBD0 U4440 ( .CLK(n4557), .C(n4558) );
  CKBD0 U4441 ( .CLK(n4558), .C(n4559) );
  BUFFD0 U4442 ( .I(n4559), .Z(n4560) );
  CKBD0 U4443 ( .CLK(n4560), .C(n4561) );
  CKBD0 U4444 ( .CLK(n4561), .C(n4562) );
  CKBD0 U4445 ( .CLK(n4562), .C(n4563) );
  CKBD0 U4446 ( .CLK(n4563), .C(n4564) );
  CKBD0 U4447 ( .CLK(n4564), .C(n4565) );
  CKBD0 U4448 ( .CLK(n4565), .C(n4566) );
  CKBD0 U4449 ( .CLK(n4566), .C(n4567) );
  CKBD0 U4450 ( .CLK(n4567), .C(n4568) );
  CKBD0 U4451 ( .CLK(n4568), .C(n4569) );
  BUFFD0 U4452 ( .I(n4569), .Z(n4570) );
  CKBD0 U4453 ( .CLK(n4570), .C(n4571) );
  CKBD0 U4454 ( .CLK(n4571), .C(n4572) );
  CKBD0 U4455 ( .CLK(n4572), .C(n4573) );
  CKBD0 U4456 ( .CLK(n4573), .C(n4574) );
  CKBD0 U4457 ( .CLK(n4574), .C(n4575) );
  CKBD0 U4458 ( .CLK(n4575), .C(n4576) );
  CKBD0 U4459 ( .CLK(n4576), .C(n4577) );
  CKBD0 U4460 ( .CLK(n4577), .C(n4578) );
  CKBD0 U4461 ( .CLK(n4578), .C(n4579) );
  CKBD0 U4462 ( .CLK(n4579), .C(n4580) );
  BUFFD0 U4463 ( .I(n4580), .Z(n4581) );
  CKBD0 U4464 ( .CLK(n4581), .C(n4582) );
  CKBD0 U4465 ( .CLK(n4582), .C(n4583) );
  CKBD0 U4466 ( .CLK(n4583), .C(n4584) );
  CKBD0 U4467 ( .CLK(n4584), .C(n4585) );
  CKBD0 U4468 ( .CLK(n4585), .C(n4586) );
  CKBD0 U4469 ( .CLK(n4586), .C(n4587) );
  CKBD0 U4470 ( .CLK(n4587), .C(n4588) );
  CKBD0 U4471 ( .CLK(n4588), .C(n4589) );
  CKBD0 U4472 ( .CLK(n4589), .C(n4590) );
  CKBD0 U4473 ( .CLK(n4590), .C(n4591) );
  BUFFD0 U4474 ( .I(n4591), .Z(n4592) );
  CKBD0 U4475 ( .CLK(n4592), .C(n4593) );
  CKBD0 U4476 ( .CLK(n4593), .C(n4594) );
  CKBD0 U4477 ( .CLK(n4594), .C(n4595) );
  CKBD0 U4478 ( .CLK(n4595), .C(n4596) );
  CKBD0 U4479 ( .CLK(n4596), .C(n4597) );
  CKBD0 U4480 ( .CLK(n4597), .C(n4598) );
  CKBD0 U4481 ( .CLK(n4598), .C(n4599) );
  CKBD0 U4482 ( .CLK(n4599), .C(n4600) );
  CKBD0 U4483 ( .CLK(n4600), .C(n4601) );
  CKBD0 U4484 ( .CLK(n4601), .C(n4602) );
  BUFFD0 U4485 ( .I(n4602), .Z(n4603) );
  CKBD0 U4486 ( .CLK(n4603), .C(n4604) );
  CKBD0 U4487 ( .CLK(n4604), .C(n4605) );
  CKBD0 U4488 ( .CLK(n4605), .C(n4606) );
  CKBD0 U4489 ( .CLK(n4606), .C(n4607) );
  CKBD0 U4490 ( .CLK(n4607), .C(n4608) );
  CKBD0 U4491 ( .CLK(n4608), .C(n4609) );
  CKBD0 U4492 ( .CLK(n4609), .C(n4610) );
  CKBD0 U4493 ( .CLK(n4610), .C(n4611) );
  CKBD0 U4494 ( .CLK(n4611), .C(n4612) );
  CKBD0 U4495 ( .CLK(n4612), .C(n4613) );
  BUFFD0 U4496 ( .I(n4613), .Z(n4614) );
  CKBD0 U4497 ( .CLK(n4614), .C(n4615) );
  CKBD0 U4498 ( .CLK(n4615), .C(n4616) );
  CKBD0 U4499 ( .CLK(n4616), .C(n4617) );
  CKBD0 U4500 ( .CLK(n4617), .C(n4618) );
  CKBD0 U4501 ( .CLK(n4618), .C(n4619) );
  CKBD0 U4502 ( .CLK(n4619), .C(n4620) );
  CKBD0 U4503 ( .CLK(n4620), .C(n4621) );
  CKBD0 U4504 ( .CLK(n4621), .C(n4622) );
  CKBD0 U4505 ( .CLK(n4622), .C(n4623) );
  CKBD0 U4506 ( .CLK(n4623), .C(n4624) );
  BUFFD0 U4507 ( .I(n4624), .Z(n4625) );
  CKBD0 U4508 ( .CLK(n4625), .C(n4626) );
  CKBD0 U4509 ( .CLK(n4626), .C(n4627) );
  CKBD0 U4510 ( .CLK(n4627), .C(n4628) );
  CKBD0 U4511 ( .CLK(n4628), .C(n4629) );
  CKBD0 U4512 ( .CLK(n4629), .C(n4630) );
  BUFFD0 U4513 ( .I(n4630), .Z(n4631) );
  CKBD0 U4514 ( .CLK(n4631), .C(n4632) );
  BUFFD0 U4515 ( .I(n4632), .Z(n4633) );
  CKBD0 U4516 ( .CLK(n4633), .C(n4634) );
  BUFFD0 U4517 ( .I(n4634), .Z(n4635) );
  CKBD0 U4518 ( .CLK(n4635), .C(n4636) );
  BUFFD0 U4519 ( .I(n4636), .Z(n4637) );
  CKBD0 U4520 ( .CLK(n4637), .C(n4638) );
  BUFFD0 U4521 ( .I(n4638), .Z(n4639) );
  CKBD0 U4522 ( .CLK(n4639), .C(n4640) );
  BUFFD0 U4523 ( .I(n4640), .Z(n4641) );
  CKBD0 U4524 ( .CLK(n4641), .C(n4642) );
  BUFFD0 U4525 ( .I(n4642), .Z(n4643) );
  CKBD0 U4526 ( .CLK(n4643), .C(n4644) );
  BUFFD0 U4527 ( .I(n4644), .Z(n4645) );
  BUFFD0 U4528 ( .I(n4647), .Z(n4646) );
  BUFFD0 U4529 ( .I(n4648), .Z(n4647) );
  BUFFD0 U4530 ( .I(n9183), .Z(n4648) );
  CKBD0 U4531 ( .CLK(n1265), .C(n4649) );
  CKBD0 U4532 ( .CLK(n4649), .C(n4650) );
  CKBD0 U4533 ( .CLK(n4650), .C(n4651) );
  CKBD0 U4534 ( .CLK(n4651), .C(n4652) );
  BUFFD0 U4535 ( .I(n4652), .Z(n4653) );
  CKBD0 U4536 ( .CLK(n4653), .C(n4654) );
  CKBD0 U4537 ( .CLK(n4654), .C(n4655) );
  CKBD0 U4538 ( .CLK(n4655), .C(n4656) );
  CKBD0 U4539 ( .CLK(n4656), .C(n4657) );
  CKBD0 U4540 ( .CLK(n4657), .C(n4658) );
  CKBD0 U4541 ( .CLK(n4658), .C(n4659) );
  CKBD0 U4542 ( .CLK(n4659), .C(n4660) );
  CKBD0 U4543 ( .CLK(n4660), .C(n4661) );
  CKBD0 U4544 ( .CLK(n4661), .C(n4662) );
  BUFFD0 U4545 ( .I(n4662), .Z(n4663) );
  CKBD0 U4546 ( .CLK(n4663), .C(n4664) );
  CKBD0 U4547 ( .CLK(n4664), .C(n4665) );
  CKBD0 U4548 ( .CLK(n4665), .C(n4666) );
  CKBD0 U4549 ( .CLK(n4666), .C(n4667) );
  CKBD0 U4550 ( .CLK(n4667), .C(n4668) );
  CKBD0 U4551 ( .CLK(n4668), .C(n4669) );
  CKBD0 U4552 ( .CLK(n4669), .C(n4670) );
  CKBD0 U4553 ( .CLK(n4670), .C(n4671) );
  CKBD0 U4554 ( .CLK(n4671), .C(n4672) );
  CKBD0 U4555 ( .CLK(n4672), .C(n4673) );
  BUFFD0 U4556 ( .I(n4673), .Z(n4674) );
  CKBD0 U4557 ( .CLK(n4674), .C(n4675) );
  CKBD0 U4558 ( .CLK(n4675), .C(n4676) );
  CKBD0 U4559 ( .CLK(n4676), .C(n4677) );
  CKBD0 U4560 ( .CLK(n4677), .C(n4678) );
  CKBD0 U4561 ( .CLK(n4678), .C(n4679) );
  CKBD0 U4562 ( .CLK(n4679), .C(n4680) );
  CKBD0 U4563 ( .CLK(n4680), .C(n4681) );
  CKBD0 U4564 ( .CLK(n4681), .C(n4682) );
  CKBD0 U4565 ( .CLK(n4682), .C(n4683) );
  CKBD0 U4566 ( .CLK(n4683), .C(n4684) );
  BUFFD0 U4567 ( .I(n4684), .Z(n4685) );
  CKBD0 U4568 ( .CLK(n4685), .C(n4686) );
  CKBD0 U4569 ( .CLK(n4686), .C(n4687) );
  CKBD0 U4570 ( .CLK(n4687), .C(n4688) );
  CKBD0 U4571 ( .CLK(n4688), .C(n4689) );
  CKBD0 U4572 ( .CLK(n4689), .C(n4690) );
  CKBD0 U4573 ( .CLK(n4690), .C(n4691) );
  CKBD0 U4574 ( .CLK(n4691), .C(n4692) );
  CKBD0 U4575 ( .CLK(n4692), .C(n4693) );
  CKBD0 U4576 ( .CLK(n4693), .C(n4694) );
  CKBD0 U4577 ( .CLK(n4694), .C(n4695) );
  BUFFD0 U4578 ( .I(n4695), .Z(n4696) );
  CKBD0 U4579 ( .CLK(n4696), .C(n4697) );
  CKBD0 U4580 ( .CLK(n4697), .C(n4698) );
  CKBD0 U4581 ( .CLK(n4698), .C(n4699) );
  CKBD0 U4582 ( .CLK(n4699), .C(n4700) );
  CKBD0 U4583 ( .CLK(n4700), .C(n4701) );
  CKBD0 U4584 ( .CLK(n4701), .C(n4702) );
  CKBD0 U4585 ( .CLK(n4702), .C(n4703) );
  CKBD0 U4586 ( .CLK(n4703), .C(n4704) );
  CKBD0 U4587 ( .CLK(n4704), .C(n4705) );
  BUFFD0 U4588 ( .I(n4705), .Z(n4706) );
  CKBD0 U4589 ( .CLK(n4706), .C(n4707) );
  CKBD0 U4590 ( .CLK(n4707), .C(n4708) );
  CKBD0 U4591 ( .CLK(n4708), .C(n4709) );
  CKBD0 U4592 ( .CLK(n4709), .C(n4710) );
  CKBD0 U4593 ( .CLK(n4710), .C(n4711) );
  CKBD0 U4594 ( .CLK(n4711), .C(n4712) );
  CKBD0 U4595 ( .CLK(n4712), .C(n4713) );
  CKBD0 U4596 ( .CLK(n4713), .C(n4714) );
  CKBD0 U4597 ( .CLK(n4714), .C(n4715) );
  CKBD0 U4598 ( .CLK(n4715), .C(n4716) );
  CKBD0 U4599 ( .CLK(n4716), .C(n4717) );
  BUFFD0 U4600 ( .I(n4717), .Z(n4718) );
  CKBD0 U4601 ( .CLK(n4718), .C(n4719) );
  CKBD0 U4602 ( .CLK(n4719), .C(n4720) );
  CKBD0 U4603 ( .CLK(n4720), .C(n4721) );
  CKBD0 U4604 ( .CLK(n4721), .C(n4722) );
  CKBD0 U4605 ( .CLK(n4722), .C(n4723) );
  CKBD0 U4606 ( .CLK(n4723), .C(n4724) );
  CKBD0 U4607 ( .CLK(n4724), .C(n4725) );
  CKBD0 U4608 ( .CLK(n4725), .C(n4726) );
  CKBD0 U4609 ( .CLK(n4726), .C(n4727) );
  BUFFD0 U4610 ( .I(n4727), .Z(n4728) );
  CKBD0 U4611 ( .CLK(n4728), .C(n4729) );
  CKBD0 U4612 ( .CLK(n4729), .C(n4730) );
  CKBD0 U4613 ( .CLK(n4730), .C(n4731) );
  CKBD0 U4614 ( .CLK(n4731), .C(n4732) );
  CKBD0 U4615 ( .CLK(n4732), .C(n4733) );
  CKBD0 U4616 ( .CLK(n4733), .C(n4734) );
  CKBD0 U4617 ( .CLK(n4734), .C(n4735) );
  CKBD0 U4618 ( .CLK(n4735), .C(n4736) );
  CKBD0 U4619 ( .CLK(n4736), .C(n4737) );
  CKBD0 U4620 ( .CLK(n4737), .C(n4738) );
  BUFFD0 U4621 ( .I(n4738), .Z(n4739) );
  CKBD0 U4622 ( .CLK(n4739), .C(n4740) );
  CKBD0 U4623 ( .CLK(n4740), .C(n4741) );
  CKBD0 U4624 ( .CLK(n4741), .C(n4742) );
  CKBD0 U4625 ( .CLK(n4742), .C(n4743) );
  CKBD0 U4626 ( .CLK(n4743), .C(n4744) );
  CKBD0 U4627 ( .CLK(n4744), .C(n4745) );
  CKBD0 U4628 ( .CLK(n4745), .C(n4746) );
  CKBD0 U4629 ( .CLK(n4746), .C(n4747) );
  CKBD0 U4630 ( .CLK(n4747), .C(n4748) );
  CKBD0 U4631 ( .CLK(n4748), .C(n4749) );
  BUFFD0 U4632 ( .I(n4749), .Z(n4750) );
  CKBD0 U4633 ( .CLK(n4750), .C(n4751) );
  CKBD0 U4634 ( .CLK(n4751), .C(n4752) );
  CKBD0 U4635 ( .CLK(n4752), .C(n4753) );
  CKBD0 U4636 ( .CLK(n4753), .C(n4754) );
  CKBD0 U4637 ( .CLK(n4754), .C(n4755) );
  CKBD0 U4638 ( .CLK(n4755), .C(n4756) );
  CKBD0 U4639 ( .CLK(n4756), .C(n4757) );
  CKBD0 U4640 ( .CLK(n4757), .C(n4758) );
  CKBD0 U4641 ( .CLK(n4758), .C(n4759) );
  CKBD0 U4642 ( .CLK(n4759), .C(n4760) );
  BUFFD0 U4643 ( .I(n4760), .Z(n4761) );
  CKBD0 U4644 ( .CLK(n4761), .C(n4762) );
  CKBD0 U4645 ( .CLK(n4762), .C(n4763) );
  CKBD0 U4646 ( .CLK(n4763), .C(n4764) );
  CKBD0 U4647 ( .CLK(n4764), .C(n4765) );
  CKBD0 U4648 ( .CLK(n4765), .C(n4766) );
  BUFFD0 U4649 ( .I(n4766), .Z(n4767) );
  CKBD0 U4650 ( .CLK(n4767), .C(n4768) );
  BUFFD0 U4651 ( .I(n4768), .Z(n4769) );
  CKBD0 U4652 ( .CLK(n4769), .C(n4770) );
  BUFFD0 U4653 ( .I(n4770), .Z(n4771) );
  CKBD0 U4654 ( .CLK(n4771), .C(n4772) );
  BUFFD0 U4655 ( .I(n4772), .Z(n4773) );
  CKBD0 U4656 ( .CLK(n4773), .C(n4774) );
  BUFFD0 U4657 ( .I(n4774), .Z(n4775) );
  CKBD0 U4658 ( .CLK(n4775), .C(n4776) );
  BUFFD0 U4659 ( .I(n4776), .Z(n4777) );
  CKBD0 U4660 ( .CLK(n4777), .C(n4778) );
  BUFFD0 U4661 ( .I(n4778), .Z(n4779) );
  CKBD0 U4662 ( .CLK(n4779), .C(n4780) );
  BUFFD0 U4663 ( .I(n4780), .Z(n4781) );
  BUFFD0 U4664 ( .I(n4783), .Z(n4782) );
  BUFFD0 U4665 ( .I(n4784), .Z(n4783) );
  BUFFD0 U4666 ( .I(n9184), .Z(n4784) );
  CKBD0 U4667 ( .CLK(n732), .C(n4785) );
  CKBD0 U4668 ( .CLK(n4785), .C(n4786) );
  CKBD0 U4669 ( .CLK(n4786), .C(n4787) );
  CKBD0 U4670 ( .CLK(n4787), .C(n4788) );
  BUFFD0 U4671 ( .I(n4788), .Z(n4789) );
  CKBD0 U4672 ( .CLK(n4789), .C(n4790) );
  CKBD0 U4673 ( .CLK(n4790), .C(n4791) );
  CKBD0 U4674 ( .CLK(n4791), .C(n4792) );
  CKBD0 U4675 ( .CLK(n4792), .C(n4793) );
  CKBD0 U4676 ( .CLK(n4793), .C(n4794) );
  CKBD0 U4677 ( .CLK(n4794), .C(n4795) );
  CKBD0 U4678 ( .CLK(n4795), .C(n4796) );
  CKBD0 U4679 ( .CLK(n4796), .C(n4797) );
  CKBD0 U4680 ( .CLK(n4797), .C(n4798) );
  BUFFD0 U4681 ( .I(n4798), .Z(n4799) );
  CKBD0 U4682 ( .CLK(n4799), .C(n4800) );
  CKBD0 U4683 ( .CLK(n4800), .C(n4801) );
  CKBD0 U4684 ( .CLK(n4801), .C(n4802) );
  CKBD0 U4685 ( .CLK(n4802), .C(n4803) );
  CKBD0 U4686 ( .CLK(n4803), .C(n4804) );
  CKBD0 U4687 ( .CLK(n4804), .C(n4805) );
  CKBD0 U4688 ( .CLK(n4805), .C(n4806) );
  CKBD0 U4689 ( .CLK(n4806), .C(n4807) );
  CKBD0 U4690 ( .CLK(n4807), .C(n4808) );
  BUFFD0 U4691 ( .I(n4808), .Z(n4809) );
  CKBD0 U4692 ( .CLK(n4809), .C(n4810) );
  CKBD0 U4693 ( .CLK(n4810), .C(n4811) );
  CKBD0 U4694 ( .CLK(n4811), .C(n4812) );
  CKBD0 U4695 ( .CLK(n4812), .C(n4813) );
  CKBD0 U4696 ( .CLK(n4813), .C(n4814) );
  CKBD0 U4697 ( .CLK(n4814), .C(n4815) );
  CKBD0 U4698 ( .CLK(n4815), .C(n4816) );
  CKBD0 U4699 ( .CLK(n4816), .C(n4817) );
  CKBD0 U4700 ( .CLK(n4817), .C(n4818) );
  CKBD0 U4701 ( .CLK(n4818), .C(n4819) );
  CKBD0 U4702 ( .CLK(n4819), .C(n4820) );
  BUFFD0 U4703 ( .I(n4820), .Z(n4821) );
  CKBD0 U4704 ( .CLK(n4821), .C(n4822) );
  CKBD0 U4705 ( .CLK(n4822), .C(n4823) );
  CKBD0 U4706 ( .CLK(n4823), .C(n4824) );
  CKBD0 U4707 ( .CLK(n4824), .C(n4825) );
  CKBD0 U4708 ( .CLK(n4825), .C(n4826) );
  CKBD0 U4709 ( .CLK(n4826), .C(n4827) );
  CKBD0 U4710 ( .CLK(n4827), .C(n4828) );
  CKBD0 U4711 ( .CLK(n4828), .C(n4829) );
  CKBD0 U4712 ( .CLK(n4829), .C(n4830) );
  BUFFD0 U4713 ( .I(n4830), .Z(n4831) );
  CKBD0 U4714 ( .CLK(n4831), .C(n4832) );
  CKBD0 U4715 ( .CLK(n4832), .C(n4833) );
  CKBD0 U4716 ( .CLK(n4833), .C(n4834) );
  CKBD0 U4717 ( .CLK(n4834), .C(n4835) );
  CKBD0 U4718 ( .CLK(n4835), .C(n4836) );
  CKBD0 U4719 ( .CLK(n4836), .C(n4837) );
  CKBD0 U4720 ( .CLK(n4837), .C(n4838) );
  CKBD0 U4721 ( .CLK(n4838), .C(n4839) );
  CKBD0 U4722 ( .CLK(n4839), .C(n4840) );
  CKBD0 U4723 ( .CLK(n4840), .C(n4841) );
  BUFFD0 U4724 ( .I(n4841), .Z(n4842) );
  CKBD0 U4725 ( .CLK(n4842), .C(n4843) );
  CKBD0 U4726 ( .CLK(n4843), .C(n4844) );
  CKBD0 U4727 ( .CLK(n4844), .C(n4845) );
  CKBD0 U4728 ( .CLK(n4845), .C(n4846) );
  CKBD0 U4729 ( .CLK(n4846), .C(n4847) );
  CKBD0 U4730 ( .CLK(n4847), .C(n4848) );
  CKBD0 U4731 ( .CLK(n4848), .C(n4849) );
  CKBD0 U4732 ( .CLK(n4849), .C(n4850) );
  CKBD0 U4733 ( .CLK(n4850), .C(n4851) );
  CKBD0 U4734 ( .CLK(n4851), .C(n4852) );
  CKBD0 U4735 ( .CLK(n4852), .C(n4853) );
  BUFFD0 U4736 ( .I(n4853), .Z(n4854) );
  CKBD0 U4737 ( .CLK(n4854), .C(n4855) );
  CKBD0 U4738 ( .CLK(n4855), .C(n4856) );
  CKBD0 U4739 ( .CLK(n4856), .C(n4857) );
  CKBD0 U4740 ( .CLK(n4857), .C(n4858) );
  CKBD0 U4741 ( .CLK(n4858), .C(n4859) );
  CKBD0 U4742 ( .CLK(n4859), .C(n4860) );
  CKBD0 U4743 ( .CLK(n4860), .C(n4861) );
  CKBD0 U4744 ( .CLK(n4861), .C(n4862) );
  CKBD0 U4745 ( .CLK(n4862), .C(n4863) );
  BUFFD0 U4746 ( .I(n4863), .Z(n4864) );
  CKBD0 U4747 ( .CLK(n4864), .C(n4865) );
  CKBD0 U4748 ( .CLK(n4865), .C(n4866) );
  CKBD0 U4749 ( .CLK(n4866), .C(n4867) );
  CKBD0 U4750 ( .CLK(n4867), .C(n4868) );
  CKBD0 U4751 ( .CLK(n4868), .C(n4869) );
  CKBD0 U4752 ( .CLK(n4869), .C(n4870) );
  CKBD0 U4753 ( .CLK(n4870), .C(n4871) );
  CKBD0 U4754 ( .CLK(n4871), .C(n4872) );
  CKBD0 U4755 ( .CLK(n4872), .C(n4873) );
  CKBD0 U4756 ( .CLK(n4873), .C(n4874) );
  BUFFD0 U4757 ( .I(n4874), .Z(n4875) );
  CKBD0 U4758 ( .CLK(n4875), .C(n4876) );
  CKBD0 U4759 ( .CLK(n4876), .C(n4877) );
  CKBD0 U4760 ( .CLK(n4877), .C(n4878) );
  CKBD0 U4761 ( .CLK(n4878), .C(n4879) );
  CKBD0 U4762 ( .CLK(n4879), .C(n4880) );
  CKBD0 U4763 ( .CLK(n4880), .C(n4881) );
  CKBD0 U4764 ( .CLK(n4881), .C(n4882) );
  CKBD0 U4765 ( .CLK(n4882), .C(n4883) );
  CKBD0 U4766 ( .CLK(n4883), .C(n4884) );
  CKBD0 U4767 ( .CLK(n4884), .C(n4885) );
  BUFFD0 U4768 ( .I(n4885), .Z(n4886) );
  CKBD0 U4769 ( .CLK(n4886), .C(n4887) );
  CKBD0 U4770 ( .CLK(n4887), .C(n4888) );
  CKBD0 U4771 ( .CLK(n4888), .C(n4889) );
  CKBD0 U4772 ( .CLK(n4889), .C(n4890) );
  CKBD0 U4773 ( .CLK(n4890), .C(n4891) );
  CKBD0 U4774 ( .CLK(n4891), .C(n4892) );
  CKBD0 U4775 ( .CLK(n4892), .C(n4893) );
  CKBD0 U4776 ( .CLK(n4893), .C(n4894) );
  CKBD0 U4777 ( .CLK(n4894), .C(n4895) );
  BUFFD0 U4778 ( .I(n4895), .Z(n4896) );
  CKBD0 U4779 ( .CLK(n4896), .C(n4897) );
  CKBD0 U4780 ( .CLK(n4897), .C(n4898) );
  CKBD0 U4781 ( .CLK(n4898), .C(n4899) );
  CKBD0 U4782 ( .CLK(n4899), .C(n4900) );
  CKBD0 U4783 ( .CLK(n4900), .C(n4901) );
  CKBD0 U4784 ( .CLK(n4901), .C(n4902) );
  BUFFD0 U4785 ( .I(n4902), .Z(n4903) );
  CKBD0 U4786 ( .CLK(n4903), .C(n4904) );
  BUFFD0 U4787 ( .I(n4904), .Z(n4905) );
  CKBD0 U4788 ( .CLK(n4905), .C(n4906) );
  BUFFD0 U4789 ( .I(n4906), .Z(n4907) );
  CKBD0 U4790 ( .CLK(n4907), .C(n4908) );
  BUFFD0 U4791 ( .I(n4908), .Z(n4909) );
  CKBD0 U4792 ( .CLK(n4909), .C(n4910) );
  BUFFD0 U4793 ( .I(n4910), .Z(n4911) );
  CKBD0 U4794 ( .CLK(n4911), .C(n4912) );
  BUFFD0 U4795 ( .I(n4912), .Z(n4913) );
  CKBD0 U4796 ( .CLK(n4913), .C(n4914) );
  BUFFD0 U4797 ( .I(n4914), .Z(n4915) );
  CKBD0 U4798 ( .CLK(n4915), .C(n4916) );
  BUFFD0 U4799 ( .I(n4916), .Z(n4917) );
  BUFFD0 U4800 ( .I(n4919), .Z(n4918) );
  BUFFD0 U4801 ( .I(n4920), .Z(n4919) );
  BUFFD0 U4802 ( .I(n9185), .Z(n4920) );
  CKBD0 U4803 ( .CLK(n1163), .C(n4921) );
  CKBD0 U4804 ( .CLK(n4921), .C(n4922) );
  CKBD0 U4805 ( .CLK(n4922), .C(n4923) );
  BUFFD0 U4806 ( .I(n4923), .Z(n4924) );
  CKBD0 U4807 ( .CLK(n4924), .C(n4925) );
  CKBD0 U4808 ( .CLK(n4925), .C(n4926) );
  CKBD0 U4809 ( .CLK(n4926), .C(n4927) );
  CKBD0 U4810 ( .CLK(n4927), .C(n4928) );
  CKBD0 U4811 ( .CLK(n4928), .C(n4929) );
  CKBD0 U4812 ( .CLK(n4929), .C(n4930) );
  CKBD0 U4813 ( .CLK(n4930), .C(n4931) );
  CKBD0 U4814 ( .CLK(n4931), .C(n4932) );
  CKBD0 U4815 ( .CLK(n4932), .C(n4933) );
  CKBD0 U4816 ( .CLK(n4933), .C(n4934) );
  BUFFD0 U4817 ( .I(n4934), .Z(n4935) );
  CKBD0 U4818 ( .CLK(n4935), .C(n4936) );
  CKBD0 U4819 ( .CLK(n4936), .C(n4937) );
  CKBD0 U4820 ( .CLK(n4937), .C(n4938) );
  CKBD0 U4821 ( .CLK(n4938), .C(n4939) );
  CKBD0 U4822 ( .CLK(n4939), .C(n4940) );
  CKBD0 U4823 ( .CLK(n4940), .C(n4941) );
  CKBD0 U4824 ( .CLK(n4941), .C(n4942) );
  CKBD0 U4825 ( .CLK(n4942), .C(n4943) );
  CKBD0 U4826 ( .CLK(n4943), .C(n4944) );
  CKBD0 U4827 ( .CLK(n4944), .C(n4945) );
  BUFFD0 U4828 ( .I(n4945), .Z(n4946) );
  CKBD0 U4829 ( .CLK(n4946), .C(n4947) );
  CKBD0 U4830 ( .CLK(n4947), .C(n4948) );
  CKBD0 U4831 ( .CLK(n4948), .C(n4949) );
  CKBD0 U4832 ( .CLK(n4949), .C(n4950) );
  CKBD0 U4833 ( .CLK(n4950), .C(n4951) );
  CKBD0 U4834 ( .CLK(n4951), .C(n4952) );
  CKBD0 U4835 ( .CLK(n4952), .C(n4953) );
  CKBD0 U4836 ( .CLK(n4953), .C(n4954) );
  CKBD0 U4837 ( .CLK(n4954), .C(n4955) );
  CKBD0 U4838 ( .CLK(n4955), .C(n4956) );
  BUFFD0 U4839 ( .I(n4956), .Z(n4957) );
  CKBD0 U4840 ( .CLK(n4957), .C(n4958) );
  CKBD0 U4841 ( .CLK(n4958), .C(n4959) );
  CKBD0 U4842 ( .CLK(n4959), .C(n4960) );
  CKBD0 U4843 ( .CLK(n4960), .C(n4961) );
  CKBD0 U4844 ( .CLK(n4961), .C(n4962) );
  CKBD0 U4845 ( .CLK(n4962), .C(n4963) );
  CKBD0 U4846 ( .CLK(n4963), .C(n4964) );
  CKBD0 U4847 ( .CLK(n4964), .C(n4965) );
  CKBD0 U4848 ( .CLK(n4965), .C(n4966) );
  BUFFD0 U4849 ( .I(n4966), .Z(n4967) );
  CKBD0 U4850 ( .CLK(n4967), .C(n4968) );
  CKBD0 U4851 ( .CLK(n4968), .C(n4969) );
  CKBD0 U4852 ( .CLK(n4969), .C(n4970) );
  CKBD0 U4853 ( .CLK(n4970), .C(n4971) );
  CKBD0 U4854 ( .CLK(n4971), .C(n4972) );
  CKBD0 U4855 ( .CLK(n4972), .C(n4973) );
  CKBD0 U4856 ( .CLK(n4973), .C(n4974) );
  CKBD0 U4857 ( .CLK(n4974), .C(n4975) );
  CKBD0 U4858 ( .CLK(n4975), .C(n4976) );
  CKBD0 U4859 ( .CLK(n4976), .C(n4977) );
  CKBD0 U4860 ( .CLK(n4977), .C(n4978) );
  BUFFD0 U4861 ( .I(n4978), .Z(n4979) );
  CKBD0 U4862 ( .CLK(n4979), .C(n4980) );
  CKBD0 U4863 ( .CLK(n4980), .C(n4981) );
  CKBD0 U4864 ( .CLK(n4981), .C(n4982) );
  CKBD0 U4865 ( .CLK(n4982), .C(n4983) );
  CKBD0 U4866 ( .CLK(n4983), .C(n4984) );
  CKBD0 U4867 ( .CLK(n4984), .C(n4985) );
  CKBD0 U4868 ( .CLK(n4985), .C(n4986) );
  CKBD0 U4869 ( .CLK(n4986), .C(n4987) );
  CKBD0 U4870 ( .CLK(n4987), .C(n4988) );
  BUFFD0 U4871 ( .I(n4988), .Z(n4989) );
  CKBD0 U4872 ( .CLK(n4989), .C(n4990) );
  CKBD0 U4873 ( .CLK(n4990), .C(n4991) );
  CKBD0 U4874 ( .CLK(n4991), .C(n4992) );
  CKBD0 U4875 ( .CLK(n4992), .C(n4993) );
  CKBD0 U4876 ( .CLK(n4993), .C(n4994) );
  CKBD0 U4877 ( .CLK(n4994), .C(n4995) );
  CKBD0 U4878 ( .CLK(n4995), .C(n4996) );
  CKBD0 U4879 ( .CLK(n4996), .C(n4997) );
  CKBD0 U4880 ( .CLK(n4997), .C(n4998) );
  CKBD0 U4881 ( .CLK(n4998), .C(n4999) );
  BUFFD0 U4882 ( .I(n4999), .Z(n5000) );
  CKBD0 U4883 ( .CLK(n5000), .C(n5001) );
  CKBD0 U4884 ( .CLK(n5001), .C(n5002) );
  CKBD0 U4885 ( .CLK(n5002), .C(n5003) );
  CKBD0 U4886 ( .CLK(n5003), .C(n5004) );
  CKBD0 U4887 ( .CLK(n5004), .C(n5005) );
  CKBD0 U4888 ( .CLK(n5005), .C(n5006) );
  CKBD0 U4889 ( .CLK(n5006), .C(n5007) );
  CKBD0 U4890 ( .CLK(n5007), .C(n5008) );
  CKBD0 U4891 ( .CLK(n5008), .C(n5009) );
  CKBD0 U4892 ( .CLK(n5009), .C(n5010) );
  BUFFD0 U4893 ( .I(n5010), .Z(n5011) );
  CKBD0 U4894 ( .CLK(n5011), .C(n5012) );
  CKBD0 U4895 ( .CLK(n5012), .C(n5013) );
  CKBD0 U4896 ( .CLK(n5013), .C(n5014) );
  CKBD0 U4897 ( .CLK(n5014), .C(n5015) );
  CKBD0 U4898 ( .CLK(n5015), .C(n5016) );
  CKBD0 U4899 ( .CLK(n5016), .C(n5017) );
  CKBD0 U4900 ( .CLK(n5017), .C(n5018) );
  CKBD0 U4901 ( .CLK(n5018), .C(n5019) );
  CKBD0 U4902 ( .CLK(n5019), .C(n5020) );
  CKBD0 U4903 ( .CLK(n5020), .C(n5021) );
  BUFFD0 U4904 ( .I(n5021), .Z(n5022) );
  CKBD0 U4905 ( .CLK(n5022), .C(n5023) );
  CKBD0 U4906 ( .CLK(n5023), .C(n5024) );
  CKBD0 U4907 ( .CLK(n5024), .C(n5025) );
  CKBD0 U4908 ( .CLK(n5025), .C(n5026) );
  CKBD0 U4909 ( .CLK(n5026), .C(n5027) );
  CKBD0 U4910 ( .CLK(n5027), .C(n5028) );
  CKBD0 U4911 ( .CLK(n5028), .C(n5029) );
  CKBD0 U4912 ( .CLK(n5029), .C(n5030) );
  CKBD0 U4913 ( .CLK(n5030), .C(n5031) );
  BUFFD0 U4914 ( .I(n5031), .Z(n5032) );
  CKBD0 U4915 ( .CLK(n5032), .C(n5033) );
  CKBD0 U4916 ( .CLK(n5033), .C(n5034) );
  CKBD0 U4917 ( .CLK(n5034), .C(n5035) );
  CKBD0 U4918 ( .CLK(n5035), .C(n5036) );
  CKBD0 U4919 ( .CLK(n5036), .C(n5037) );
  CKBD0 U4920 ( .CLK(n5037), .C(n5038) );
  BUFFD0 U4921 ( .I(n5038), .Z(n5039) );
  CKBD0 U4922 ( .CLK(n5039), .C(n5040) );
  BUFFD0 U4923 ( .I(n5040), .Z(n5041) );
  CKBD0 U4924 ( .CLK(n5041), .C(n5042) );
  BUFFD0 U4925 ( .I(n5042), .Z(n5043) );
  CKBD0 U4926 ( .CLK(n5043), .C(n5044) );
  BUFFD0 U4927 ( .I(n5044), .Z(n5045) );
  CKBD0 U4928 ( .CLK(n5045), .C(n5046) );
  BUFFD0 U4929 ( .I(n5046), .Z(n5047) );
  CKBD0 U4930 ( .CLK(n5047), .C(n5048) );
  BUFFD0 U4931 ( .I(n5048), .Z(n5049) );
  CKBD0 U4932 ( .CLK(n5049), .C(n5050) );
  BUFFD0 U4933 ( .I(n5050), .Z(n5051) );
  CKBD0 U4934 ( .CLK(n5051), .C(n5052) );
  BUFFD0 U4935 ( .I(n5052), .Z(n5053) );
  BUFFD0 U4936 ( .I(n5055), .Z(n5054) );
  BUFFD0 U4937 ( .I(n5056), .Z(n5055) );
  BUFFD0 U4938 ( .I(n9186), .Z(n5056) );
  CKBD0 U4939 ( .CLK(n1161), .C(n5057) );
  CKBD0 U4940 ( .CLK(n5057), .C(n5058) );
  CKBD0 U4941 ( .CLK(n5058), .C(n5059) );
  BUFFD0 U4942 ( .I(n5059), .Z(n5060) );
  CKBD0 U4943 ( .CLK(n5060), .C(n5061) );
  CKBD0 U4944 ( .CLK(n5061), .C(n5062) );
  CKBD0 U4945 ( .CLK(n5062), .C(n5063) );
  CKBD0 U4946 ( .CLK(n5063), .C(n5064) );
  CKBD0 U4947 ( .CLK(n5064), .C(n5065) );
  CKBD0 U4948 ( .CLK(n5065), .C(n5066) );
  CKBD0 U4949 ( .CLK(n5066), .C(n5067) );
  CKBD0 U4950 ( .CLK(n5067), .C(n5068) );
  CKBD0 U4951 ( .CLK(n5068), .C(n5069) );
  CKBD0 U4952 ( .CLK(n5069), .C(n5070) );
  BUFFD0 U4953 ( .I(n5070), .Z(n5071) );
  CKBD0 U4954 ( .CLK(n5071), .C(n5072) );
  CKBD0 U4955 ( .CLK(n5072), .C(n5073) );
  CKBD0 U4956 ( .CLK(n5073), .C(n5074) );
  CKBD0 U4957 ( .CLK(n5074), .C(n5075) );
  CKBD0 U4958 ( .CLK(n5075), .C(n5076) );
  CKBD0 U4959 ( .CLK(n5076), .C(n5077) );
  CKBD0 U4960 ( .CLK(n5077), .C(n5078) );
  CKBD0 U4961 ( .CLK(n5078), .C(n5079) );
  CKBD0 U4962 ( .CLK(n5079), .C(n5080) );
  CKBD0 U4963 ( .CLK(n5080), .C(n5081) );
  BUFFD0 U4964 ( .I(n5081), .Z(n5082) );
  CKBD0 U4965 ( .CLK(n5082), .C(n5083) );
  CKBD0 U4966 ( .CLK(n5083), .C(n5084) );
  CKBD0 U4967 ( .CLK(n5084), .C(n5085) );
  CKBD0 U4968 ( .CLK(n5085), .C(n5086) );
  CKBD0 U4969 ( .CLK(n5086), .C(n5087) );
  CKBD0 U4970 ( .CLK(n5087), .C(n5088) );
  CKBD0 U4971 ( .CLK(n5088), .C(n5089) );
  CKBD0 U4972 ( .CLK(n5089), .C(n5090) );
  CKBD0 U4973 ( .CLK(n5090), .C(n5091) );
  CKBD0 U4974 ( .CLK(n5091), .C(n5092) );
  BUFFD0 U4975 ( .I(n5092), .Z(n5093) );
  CKBD0 U4976 ( .CLK(n5093), .C(n5094) );
  CKBD0 U4977 ( .CLK(n5094), .C(n5095) );
  CKBD0 U4978 ( .CLK(n5095), .C(n5096) );
  CKBD0 U4979 ( .CLK(n5096), .C(n5097) );
  CKBD0 U4980 ( .CLK(n5097), .C(n5098) );
  CKBD0 U4981 ( .CLK(n5098), .C(n5099) );
  CKBD0 U4982 ( .CLK(n5099), .C(n5100) );
  CKBD0 U4983 ( .CLK(n5100), .C(n5101) );
  CKBD0 U4984 ( .CLK(n5101), .C(n5102) );
  BUFFD0 U4985 ( .I(n5102), .Z(n5103) );
  CKBD0 U4986 ( .CLK(n5103), .C(n5104) );
  CKBD0 U4987 ( .CLK(n5104), .C(n5105) );
  CKBD0 U4988 ( .CLK(n5105), .C(n5106) );
  CKBD0 U4989 ( .CLK(n5106), .C(n5107) );
  CKBD0 U4990 ( .CLK(n5107), .C(n5108) );
  CKBD0 U4991 ( .CLK(n5108), .C(n5109) );
  CKBD0 U4992 ( .CLK(n5109), .C(n5110) );
  CKBD0 U4993 ( .CLK(n5110), .C(n5111) );
  CKBD0 U4994 ( .CLK(n5111), .C(n5112) );
  CKBD0 U4995 ( .CLK(n5112), .C(n5113) );
  CKBD0 U4996 ( .CLK(n5113), .C(n5114) );
  BUFFD0 U4997 ( .I(n5114), .Z(n5115) );
  CKBD0 U4998 ( .CLK(n5115), .C(n5116) );
  CKBD0 U4999 ( .CLK(n5116), .C(n5117) );
  CKBD0 U5000 ( .CLK(n5117), .C(n5118) );
  CKBD0 U5001 ( .CLK(n5118), .C(n5119) );
  CKBD0 U5002 ( .CLK(n5119), .C(n5120) );
  CKBD0 U5003 ( .CLK(n5120), .C(n5121) );
  CKBD0 U5004 ( .CLK(n5121), .C(n5122) );
  CKBD0 U5005 ( .CLK(n5122), .C(n5123) );
  CKBD0 U5006 ( .CLK(n5123), .C(n5124) );
  BUFFD0 U5007 ( .I(n5124), .Z(n5125) );
  CKBD0 U5008 ( .CLK(n5125), .C(n5126) );
  CKBD0 U5009 ( .CLK(n5126), .C(n5127) );
  CKBD0 U5010 ( .CLK(n5127), .C(n5128) );
  CKBD0 U5011 ( .CLK(n5128), .C(n5129) );
  CKBD0 U5012 ( .CLK(n5129), .C(n5130) );
  CKBD0 U5013 ( .CLK(n5130), .C(n5131) );
  CKBD0 U5014 ( .CLK(n5131), .C(n5132) );
  CKBD0 U5015 ( .CLK(n5132), .C(n5133) );
  CKBD0 U5016 ( .CLK(n5133), .C(n5134) );
  CKBD0 U5017 ( .CLK(n5134), .C(n5135) );
  BUFFD0 U5018 ( .I(n5135), .Z(n5136) );
  CKBD0 U5019 ( .CLK(n5136), .C(n5137) );
  CKBD0 U5020 ( .CLK(n5137), .C(n5138) );
  CKBD0 U5021 ( .CLK(n5138), .C(n5139) );
  CKBD0 U5022 ( .CLK(n5139), .C(n5140) );
  CKBD0 U5023 ( .CLK(n5140), .C(n5141) );
  CKBD0 U5024 ( .CLK(n5141), .C(n5142) );
  CKBD0 U5025 ( .CLK(n5142), .C(n5143) );
  CKBD0 U5026 ( .CLK(n5143), .C(n5144) );
  CKBD0 U5027 ( .CLK(n5144), .C(n5145) );
  CKBD0 U5028 ( .CLK(n5145), .C(n5146) );
  BUFFD0 U5029 ( .I(n5146), .Z(n5147) );
  CKBD0 U5030 ( .CLK(n5147), .C(n5148) );
  CKBD0 U5031 ( .CLK(n5148), .C(n5149) );
  CKBD0 U5032 ( .CLK(n5149), .C(n5150) );
  CKBD0 U5033 ( .CLK(n5150), .C(n5151) );
  CKBD0 U5034 ( .CLK(n5151), .C(n5152) );
  CKBD0 U5035 ( .CLK(n5152), .C(n5153) );
  CKBD0 U5036 ( .CLK(n5153), .C(n5154) );
  CKBD0 U5037 ( .CLK(n5154), .C(n5155) );
  CKBD0 U5038 ( .CLK(n5155), .C(n5156) );
  CKBD0 U5039 ( .CLK(n5156), .C(n5157) );
  BUFFD0 U5040 ( .I(n5157), .Z(n5158) );
  CKBD0 U5041 ( .CLK(n5158), .C(n5159) );
  CKBD0 U5042 ( .CLK(n5159), .C(n5160) );
  CKBD0 U5043 ( .CLK(n5160), .C(n5161) );
  CKBD0 U5044 ( .CLK(n5161), .C(n5162) );
  CKBD0 U5045 ( .CLK(n5162), .C(n5163) );
  CKBD0 U5046 ( .CLK(n5163), .C(n5164) );
  CKBD0 U5047 ( .CLK(n5164), .C(n5165) );
  CKBD0 U5048 ( .CLK(n5165), .C(n5166) );
  CKBD0 U5049 ( .CLK(n5166), .C(n5167) );
  CKBD0 U5050 ( .CLK(n5167), .C(n5168) );
  BUFFD0 U5051 ( .I(n5168), .Z(n5169) );
  CKBD0 U5052 ( .CLK(n5169), .C(n5170) );
  CKBD0 U5053 ( .CLK(n5170), .C(n5171) );
  CKBD0 U5054 ( .CLK(n5171), .C(n5172) );
  CKBD0 U5055 ( .CLK(n5172), .C(n5173) );
  CKBD0 U5056 ( .CLK(n5173), .C(n5174) );
  BUFFD0 U5057 ( .I(n5174), .Z(n5175) );
  CKBD0 U5058 ( .CLK(n5175), .C(n5176) );
  BUFFD0 U5059 ( .I(n5176), .Z(n5177) );
  CKBD0 U5060 ( .CLK(n5177), .C(n5178) );
  BUFFD0 U5061 ( .I(n5178), .Z(n5179) );
  CKBD0 U5062 ( .CLK(n5179), .C(n5180) );
  BUFFD0 U5063 ( .I(n5180), .Z(n5181) );
  CKBD0 U5064 ( .CLK(n5181), .C(n5182) );
  BUFFD0 U5065 ( .I(n5182), .Z(n5183) );
  CKBD0 U5066 ( .CLK(n5183), .C(n5184) );
  BUFFD0 U5067 ( .I(n5184), .Z(n5185) );
  CKBD0 U5068 ( .CLK(n5185), .C(n5186) );
  BUFFD0 U5069 ( .I(n5186), .Z(n5187) );
  CKBD0 U5070 ( .CLK(n5187), .C(n5188) );
  BUFFD0 U5071 ( .I(n5188), .Z(n5189) );
  BUFFD0 U5072 ( .I(Decoder[12]), .Z(n5190) );
  BUFFD0 U5073 ( .I(n5192), .Z(n5191) );
  BUFFD0 U5074 ( .I(n5193), .Z(n5192) );
  BUFFD0 U5075 ( .I(n9187), .Z(n5193) );
  CKBD0 U5076 ( .CLK(n1159), .C(n5194) );
  CKBD0 U5077 ( .CLK(n5194), .C(n5195) );
  CKBD0 U5078 ( .CLK(n5195), .C(n5196) );
  CKBD0 U5079 ( .CLK(n5196), .C(n5197) );
  BUFFD0 U5080 ( .I(n5197), .Z(n5198) );
  CKBD0 U5081 ( .CLK(n5198), .C(n5199) );
  CKBD0 U5082 ( .CLK(n5199), .C(n5200) );
  CKBD0 U5083 ( .CLK(n5200), .C(n5201) );
  CKBD0 U5084 ( .CLK(n5201), .C(n5202) );
  CKBD0 U5085 ( .CLK(n5202), .C(n5203) );
  CKBD0 U5086 ( .CLK(n5203), .C(n5204) );
  CKBD0 U5087 ( .CLK(n5204), .C(n5205) );
  CKBD0 U5088 ( .CLK(n5205), .C(n5206) );
  CKBD0 U5089 ( .CLK(n5206), .C(n5207) );
  BUFFD0 U5090 ( .I(n5207), .Z(n5208) );
  CKBD0 U5091 ( .CLK(n5208), .C(n5209) );
  CKBD0 U5092 ( .CLK(n5209), .C(n5210) );
  CKBD0 U5093 ( .CLK(n5210), .C(n5211) );
  CKBD0 U5094 ( .CLK(n5211), .C(n5212) );
  CKBD0 U5095 ( .CLK(n5212), .C(n5213) );
  CKBD0 U5096 ( .CLK(n5213), .C(n5214) );
  CKBD0 U5097 ( .CLK(n5214), .C(n5215) );
  CKBD0 U5098 ( .CLK(n5215), .C(n5216) );
  CKBD0 U5099 ( .CLK(n5216), .C(n5217) );
  BUFFD0 U5100 ( .I(n5217), .Z(n5218) );
  CKBD0 U5101 ( .CLK(n5218), .C(n5219) );
  CKBD0 U5102 ( .CLK(n5219), .C(n5220) );
  CKBD0 U5103 ( .CLK(n5220), .C(n5221) );
  CKBD0 U5104 ( .CLK(n5221), .C(n5222) );
  CKBD0 U5105 ( .CLK(n5222), .C(n5223) );
  CKBD0 U5106 ( .CLK(n5223), .C(n5224) );
  CKBD0 U5107 ( .CLK(n5224), .C(n5225) );
  CKBD0 U5108 ( .CLK(n5225), .C(n5226) );
  CKBD0 U5109 ( .CLK(n5226), .C(n5227) );
  CKBD0 U5110 ( .CLK(n5227), .C(n5228) );
  CKBD0 U5111 ( .CLK(n5228), .C(n5229) );
  BUFFD0 U5112 ( .I(n5229), .Z(n5230) );
  CKBD0 U5113 ( .CLK(n5230), .C(n5231) );
  CKBD0 U5114 ( .CLK(n5231), .C(n5232) );
  CKBD0 U5115 ( .CLK(n5232), .C(n5233) );
  CKBD0 U5116 ( .CLK(n5233), .C(n5234) );
  CKBD0 U5117 ( .CLK(n5234), .C(n5235) );
  CKBD0 U5118 ( .CLK(n5235), .C(n5236) );
  CKBD0 U5119 ( .CLK(n5236), .C(n5237) );
  CKBD0 U5120 ( .CLK(n5237), .C(n5238) );
  CKBD0 U5121 ( .CLK(n5238), .C(n5239) );
  CKBD0 U5122 ( .CLK(n5239), .C(n5240) );
  BUFFD0 U5123 ( .I(n5240), .Z(n5241) );
  CKBD0 U5124 ( .CLK(n5241), .C(n5242) );
  CKBD0 U5125 ( .CLK(n5242), .C(n5243) );
  CKBD0 U5126 ( .CLK(n5243), .C(n5244) );
  CKBD0 U5127 ( .CLK(n5244), .C(n5245) );
  CKBD0 U5128 ( .CLK(n5245), .C(n5246) );
  CKBD0 U5129 ( .CLK(n5246), .C(n5247) );
  CKBD0 U5130 ( .CLK(n5247), .C(n5248) );
  CKBD0 U5131 ( .CLK(n5248), .C(n5249) );
  CKBD0 U5132 ( .CLK(n5249), .C(n5250) );
  BUFFD0 U5133 ( .I(n5250), .Z(n5251) );
  CKBD0 U5134 ( .CLK(n5251), .C(n5252) );
  CKBD0 U5135 ( .CLK(n5252), .C(n5253) );
  CKBD0 U5136 ( .CLK(n5253), .C(n5254) );
  CKBD0 U5137 ( .CLK(n5254), .C(n5255) );
  CKBD0 U5138 ( .CLK(n5255), .C(n5256) );
  CKBD0 U5139 ( .CLK(n5256), .C(n5257) );
  CKBD0 U5140 ( .CLK(n5257), .C(n5258) );
  CKBD0 U5141 ( .CLK(n5258), .C(n5259) );
  CKBD0 U5142 ( .CLK(n5259), .C(n5260) );
  CKBD0 U5143 ( .CLK(n5260), .C(n5261) );
  CKBD0 U5144 ( .CLK(n5261), .C(n5262) );
  BUFFD0 U5145 ( .I(n5262), .Z(n5263) );
  CKBD0 U5146 ( .CLK(n5263), .C(n5264) );
  CKBD0 U5147 ( .CLK(n5264), .C(n5265) );
  CKBD0 U5148 ( .CLK(n5265), .C(n5266) );
  CKBD0 U5149 ( .CLK(n5266), .C(n5267) );
  CKBD0 U5150 ( .CLK(n5267), .C(n5268) );
  CKBD0 U5151 ( .CLK(n5268), .C(n5269) );
  CKBD0 U5152 ( .CLK(n5269), .C(n5270) );
  CKBD0 U5153 ( .CLK(n5270), .C(n5271) );
  CKBD0 U5154 ( .CLK(n5271), .C(n5272) );
  BUFFD0 U5155 ( .I(n5272), .Z(n5273) );
  CKBD0 U5156 ( .CLK(n5273), .C(n5274) );
  CKBD0 U5157 ( .CLK(n5274), .C(n5275) );
  CKBD0 U5158 ( .CLK(n5275), .C(n5276) );
  CKBD0 U5159 ( .CLK(n5276), .C(n5277) );
  CKBD0 U5160 ( .CLK(n5277), .C(n5278) );
  CKBD0 U5161 ( .CLK(n5278), .C(n5279) );
  CKBD0 U5162 ( .CLK(n5279), .C(n5280) );
  CKBD0 U5163 ( .CLK(n5280), .C(n5281) );
  CKBD0 U5164 ( .CLK(n5281), .C(n5282) );
  CKBD0 U5165 ( .CLK(n5282), .C(n5283) );
  BUFFD0 U5166 ( .I(n5283), .Z(n5284) );
  CKBD0 U5167 ( .CLK(n5284), .C(n5285) );
  CKBD0 U5168 ( .CLK(n5285), .C(n5286) );
  CKBD0 U5169 ( .CLK(n5286), .C(n5287) );
  CKBD0 U5170 ( .CLK(n5287), .C(n5288) );
  CKBD0 U5171 ( .CLK(n5288), .C(n5289) );
  CKBD0 U5172 ( .CLK(n5289), .C(n5290) );
  CKBD0 U5173 ( .CLK(n5290), .C(n5291) );
  CKBD0 U5174 ( .CLK(n5291), .C(n5292) );
  CKBD0 U5175 ( .CLK(n5292), .C(n5293) );
  CKBD0 U5176 ( .CLK(n5293), .C(n5294) );
  BUFFD0 U5177 ( .I(n5294), .Z(n5295) );
  CKBD0 U5178 ( .CLK(n5295), .C(n5296) );
  CKBD0 U5179 ( .CLK(n5296), .C(n5297) );
  CKBD0 U5180 ( .CLK(n5297), .C(n5298) );
  CKBD0 U5181 ( .CLK(n5298), .C(n5299) );
  CKBD0 U5182 ( .CLK(n5299), .C(n5300) );
  CKBD0 U5183 ( .CLK(n5300), .C(n5301) );
  CKBD0 U5184 ( .CLK(n5301), .C(n5302) );
  CKBD0 U5185 ( .CLK(n5302), .C(n5303) );
  CKBD0 U5186 ( .CLK(n5303), .C(n5304) );
  BUFFD0 U5187 ( .I(n5304), .Z(n5305) );
  CKBD0 U5188 ( .CLK(n5305), .C(n5306) );
  CKBD0 U5189 ( .CLK(n5306), .C(n5307) );
  CKBD0 U5190 ( .CLK(n5307), .C(n5308) );
  CKBD0 U5191 ( .CLK(n5308), .C(n5309) );
  CKBD0 U5192 ( .CLK(n5309), .C(n5310) );
  CKBD0 U5193 ( .CLK(n5310), .C(n5311) );
  BUFFD0 U5194 ( .I(n5311), .Z(n5312) );
  CKBD0 U5195 ( .CLK(n5312), .C(n5313) );
  BUFFD0 U5196 ( .I(n5313), .Z(n5314) );
  CKBD0 U5197 ( .CLK(n5314), .C(n5315) );
  BUFFD0 U5198 ( .I(n5315), .Z(n5316) );
  CKBD0 U5199 ( .CLK(n5316), .C(n5317) );
  BUFFD0 U5200 ( .I(n5317), .Z(n5318) );
  CKBD0 U5201 ( .CLK(n5318), .C(n5319) );
  BUFFD0 U5202 ( .I(n5319), .Z(n5320) );
  CKBD0 U5203 ( .CLK(n5320), .C(n5321) );
  BUFFD0 U5204 ( .I(n5321), .Z(n5322) );
  CKBD0 U5205 ( .CLK(n5322), .C(n5323) );
  BUFFD0 U5206 ( .I(n5323), .Z(n5324) );
  CKBD0 U5207 ( .CLK(n5324), .C(n5325) );
  BUFFD0 U5208 ( .I(n5325), .Z(n5326) );
  BUFFD0 U5209 ( .I(n5328), .Z(n5327) );
  BUFFD0 U5210 ( .I(n5329), .Z(n5328) );
  BUFFD0 U5211 ( .I(n9188), .Z(n5329) );
  CKBD0 U5212 ( .CLK(n1157), .C(n5330) );
  CKBD0 U5213 ( .CLK(n5330), .C(n5331) );
  CKBD0 U5214 ( .CLK(n5331), .C(n5332) );
  BUFFD0 U5215 ( .I(n5332), .Z(n5333) );
  CKBD0 U5216 ( .CLK(n5333), .C(n5334) );
  CKBD0 U5217 ( .CLK(n5334), .C(n5335) );
  CKBD0 U5218 ( .CLK(n5335), .C(n5336) );
  CKBD0 U5219 ( .CLK(n5336), .C(n5337) );
  CKBD0 U5220 ( .CLK(n5337), .C(n5338) );
  CKBD0 U5221 ( .CLK(n5338), .C(n5339) );
  CKBD0 U5222 ( .CLK(n5339), .C(n5340) );
  CKBD0 U5223 ( .CLK(n5340), .C(n5341) );
  CKBD0 U5224 ( .CLK(n5341), .C(n5342) );
  CKBD0 U5225 ( .CLK(n5342), .C(n5343) );
  BUFFD0 U5226 ( .I(n5343), .Z(n5344) );
  CKBD0 U5227 ( .CLK(n5344), .C(n5345) );
  CKBD0 U5228 ( .CLK(n5345), .C(n5346) );
  CKBD0 U5229 ( .CLK(n5346), .C(n5347) );
  CKBD0 U5230 ( .CLK(n5347), .C(n5348) );
  CKBD0 U5231 ( .CLK(n5348), .C(n5349) );
  CKBD0 U5232 ( .CLK(n5349), .C(n5350) );
  CKBD0 U5233 ( .CLK(n5350), .C(n5351) );
  CKBD0 U5234 ( .CLK(n5351), .C(n5352) );
  CKBD0 U5235 ( .CLK(n5352), .C(n5353) );
  CKBD0 U5236 ( .CLK(n5353), .C(n5354) );
  BUFFD0 U5237 ( .I(n5354), .Z(n5355) );
  CKBD0 U5238 ( .CLK(n5355), .C(n5356) );
  CKBD0 U5239 ( .CLK(n5356), .C(n5357) );
  CKBD0 U5240 ( .CLK(n5357), .C(n5358) );
  CKBD0 U5241 ( .CLK(n5358), .C(n5359) );
  CKBD0 U5242 ( .CLK(n5359), .C(n5360) );
  CKBD0 U5243 ( .CLK(n5360), .C(n5361) );
  CKBD0 U5244 ( .CLK(n5361), .C(n5362) );
  CKBD0 U5245 ( .CLK(n5362), .C(n5363) );
  CKBD0 U5246 ( .CLK(n5363), .C(n5364) );
  CKBD0 U5247 ( .CLK(n5364), .C(n5365) );
  BUFFD0 U5248 ( .I(n5365), .Z(n5366) );
  CKBD0 U5249 ( .CLK(n5366), .C(n5367) );
  CKBD0 U5250 ( .CLK(n5367), .C(n5368) );
  CKBD0 U5251 ( .CLK(n5368), .C(n5369) );
  CKBD0 U5252 ( .CLK(n5369), .C(n5370) );
  CKBD0 U5253 ( .CLK(n5370), .C(n5371) );
  CKBD0 U5254 ( .CLK(n5371), .C(n5372) );
  CKBD0 U5255 ( .CLK(n5372), .C(n5373) );
  CKBD0 U5256 ( .CLK(n5373), .C(n5374) );
  CKBD0 U5257 ( .CLK(n5374), .C(n5375) );
  BUFFD0 U5258 ( .I(n5375), .Z(n5376) );
  CKBD0 U5259 ( .CLK(n5376), .C(n5377) );
  CKBD0 U5260 ( .CLK(n5377), .C(n5378) );
  CKBD0 U5261 ( .CLK(n5378), .C(n5379) );
  CKBD0 U5262 ( .CLK(n5379), .C(n5380) );
  CKBD0 U5263 ( .CLK(n5380), .C(n5381) );
  CKBD0 U5264 ( .CLK(n5381), .C(n5382) );
  CKBD0 U5265 ( .CLK(n5382), .C(n5383) );
  CKBD0 U5266 ( .CLK(n5383), .C(n5384) );
  CKBD0 U5267 ( .CLK(n5384), .C(n5385) );
  CKBD0 U5268 ( .CLK(n5385), .C(n5386) );
  CKBD0 U5269 ( .CLK(n5386), .C(n5387) );
  BUFFD0 U5270 ( .I(n5387), .Z(n5388) );
  CKBD0 U5271 ( .CLK(n5388), .C(n5389) );
  CKBD0 U5272 ( .CLK(n5389), .C(n5390) );
  CKBD0 U5273 ( .CLK(n5390), .C(n5391) );
  CKBD0 U5274 ( .CLK(n5391), .C(n5392) );
  CKBD0 U5275 ( .CLK(n5392), .C(n5393) );
  CKBD0 U5276 ( .CLK(n5393), .C(n5394) );
  CKBD0 U5277 ( .CLK(n5394), .C(n5395) );
  CKBD0 U5278 ( .CLK(n5395), .C(n5396) );
  CKBD0 U5279 ( .CLK(n5396), .C(n5397) );
  BUFFD0 U5280 ( .I(n5397), .Z(n5398) );
  CKBD0 U5281 ( .CLK(n5398), .C(n5399) );
  CKBD0 U5282 ( .CLK(n5399), .C(n5400) );
  CKBD0 U5283 ( .CLK(n5400), .C(n5401) );
  CKBD0 U5284 ( .CLK(n5401), .C(n5402) );
  CKBD0 U5285 ( .CLK(n5402), .C(n5403) );
  CKBD0 U5286 ( .CLK(n5403), .C(n5404) );
  CKBD0 U5287 ( .CLK(n5404), .C(n5405) );
  CKBD0 U5288 ( .CLK(n5405), .C(n5406) );
  CKBD0 U5289 ( .CLK(n5406), .C(n5407) );
  CKBD0 U5290 ( .CLK(n5407), .C(n5408) );
  BUFFD0 U5291 ( .I(n5408), .Z(n5409) );
  CKBD0 U5292 ( .CLK(n5409), .C(n5410) );
  CKBD0 U5293 ( .CLK(n5410), .C(n5411) );
  CKBD0 U5294 ( .CLK(n5411), .C(n5412) );
  CKBD0 U5295 ( .CLK(n5412), .C(n5413) );
  CKBD0 U5296 ( .CLK(n5413), .C(n5414) );
  CKBD0 U5297 ( .CLK(n5414), .C(n5415) );
  CKBD0 U5298 ( .CLK(n5415), .C(n5416) );
  CKBD0 U5299 ( .CLK(n5416), .C(n5417) );
  CKBD0 U5300 ( .CLK(n5417), .C(n5418) );
  CKBD0 U5301 ( .CLK(n5418), .C(n5419) );
  BUFFD0 U5302 ( .I(n5419), .Z(n5420) );
  CKBD0 U5303 ( .CLK(n5420), .C(n5421) );
  CKBD0 U5304 ( .CLK(n5421), .C(n5422) );
  CKBD0 U5305 ( .CLK(n5422), .C(n5423) );
  CKBD0 U5306 ( .CLK(n5423), .C(n5424) );
  CKBD0 U5307 ( .CLK(n5424), .C(n5425) );
  CKBD0 U5308 ( .CLK(n5425), .C(n5426) );
  CKBD0 U5309 ( .CLK(n5426), .C(n5427) );
  CKBD0 U5310 ( .CLK(n5427), .C(n5428) );
  CKBD0 U5311 ( .CLK(n5428), .C(n5429) );
  CKBD0 U5312 ( .CLK(n5429), .C(n5430) );
  BUFFD0 U5313 ( .I(n5430), .Z(n5431) );
  CKBD0 U5314 ( .CLK(n5431), .C(n5432) );
  CKBD0 U5315 ( .CLK(n5432), .C(n5433) );
  CKBD0 U5316 ( .CLK(n5433), .C(n5434) );
  CKBD0 U5317 ( .CLK(n5434), .C(n5435) );
  CKBD0 U5318 ( .CLK(n5435), .C(n5436) );
  CKBD0 U5319 ( .CLK(n5436), .C(n5437) );
  CKBD0 U5320 ( .CLK(n5437), .C(n5438) );
  CKBD0 U5321 ( .CLK(n5438), .C(n5439) );
  CKBD0 U5322 ( .CLK(n5439), .C(n5440) );
  BUFFD0 U5323 ( .I(n5440), .Z(n5441) );
  CKBD0 U5324 ( .CLK(n5441), .C(n5442) );
  CKBD0 U5325 ( .CLK(n5442), .C(n5443) );
  CKBD0 U5326 ( .CLK(n5443), .C(n5444) );
  CKBD0 U5327 ( .CLK(n5444), .C(n5445) );
  CKBD0 U5328 ( .CLK(n5445), .C(n5446) );
  CKBD0 U5329 ( .CLK(n5446), .C(n5447) );
  BUFFD0 U5330 ( .I(n5447), .Z(n5448) );
  CKBD0 U5331 ( .CLK(n5448), .C(n5449) );
  BUFFD0 U5332 ( .I(n5449), .Z(n5450) );
  CKBD0 U5333 ( .CLK(n5450), .C(n5451) );
  BUFFD0 U5334 ( .I(n5451), .Z(n5452) );
  CKBD0 U5335 ( .CLK(n5452), .C(n5453) );
  BUFFD0 U5336 ( .I(n5453), .Z(n5454) );
  CKBD0 U5337 ( .CLK(n5454), .C(n5455) );
  BUFFD0 U5338 ( .I(n5455), .Z(n5456) );
  CKBD0 U5339 ( .CLK(n5456), .C(n5457) );
  BUFFD0 U5340 ( .I(n5457), .Z(n5458) );
  CKBD0 U5341 ( .CLK(n5458), .C(n5459) );
  BUFFD0 U5342 ( .I(n5459), .Z(n5460) );
  CKBD0 U5343 ( .CLK(n5460), .C(n5461) );
  BUFFD0 U5344 ( .I(n5461), .Z(n5462) );
  BUFFD0 U5345 ( .I(n5464), .Z(n5463) );
  BUFFD0 U5346 ( .I(n5465), .Z(n5464) );
  BUFFD0 U5347 ( .I(n9189), .Z(n5465) );
  CKBD0 U5348 ( .CLK(n1155), .C(n5466) );
  CKBD0 U5349 ( .CLK(n5466), .C(n5467) );
  CKBD0 U5350 ( .CLK(n5467), .C(n5468) );
  BUFFD0 U5351 ( .I(n5468), .Z(n5469) );
  CKBD0 U5352 ( .CLK(n5469), .C(n5470) );
  CKBD0 U5353 ( .CLK(n5470), .C(n5471) );
  CKBD0 U5354 ( .CLK(n5471), .C(n5472) );
  CKBD0 U5355 ( .CLK(n5472), .C(n5473) );
  CKBD0 U5356 ( .CLK(n5473), .C(n5474) );
  CKBD0 U5357 ( .CLK(n5474), .C(n5475) );
  CKBD0 U5358 ( .CLK(n5475), .C(n5476) );
  CKBD0 U5359 ( .CLK(n5476), .C(n5477) );
  CKBD0 U5360 ( .CLK(n5477), .C(n5478) );
  CKBD0 U5361 ( .CLK(n5478), .C(n5479) );
  BUFFD0 U5362 ( .I(n5479), .Z(n5480) );
  CKBD0 U5363 ( .CLK(n5480), .C(n5481) );
  CKBD0 U5364 ( .CLK(n5481), .C(n5482) );
  CKBD0 U5365 ( .CLK(n5482), .C(n5483) );
  CKBD0 U5366 ( .CLK(n5483), .C(n5484) );
  CKBD0 U5367 ( .CLK(n5484), .C(n5485) );
  CKBD0 U5368 ( .CLK(n5485), .C(n5486) );
  CKBD0 U5369 ( .CLK(n5486), .C(n5487) );
  CKBD0 U5370 ( .CLK(n5487), .C(n5488) );
  CKBD0 U5371 ( .CLK(n5488), .C(n5489) );
  CKBD0 U5372 ( .CLK(n5489), .C(n5490) );
  BUFFD0 U5373 ( .I(n5490), .Z(n5491) );
  CKBD0 U5374 ( .CLK(n5491), .C(n5492) );
  CKBD0 U5375 ( .CLK(n5492), .C(n5493) );
  CKBD0 U5376 ( .CLK(n5493), .C(n5494) );
  CKBD0 U5377 ( .CLK(n5494), .C(n5495) );
  CKBD0 U5378 ( .CLK(n5495), .C(n5496) );
  CKBD0 U5379 ( .CLK(n5496), .C(n5497) );
  CKBD0 U5380 ( .CLK(n5497), .C(n5498) );
  CKBD0 U5381 ( .CLK(n5498), .C(n5499) );
  CKBD0 U5382 ( .CLK(n5499), .C(n5500) );
  CKBD0 U5383 ( .CLK(n5500), .C(n5501) );
  BUFFD0 U5384 ( .I(n5501), .Z(n5502) );
  CKBD0 U5385 ( .CLK(n5502), .C(n5503) );
  CKBD0 U5386 ( .CLK(n5503), .C(n5504) );
  CKBD0 U5387 ( .CLK(n5504), .C(n5505) );
  CKBD0 U5388 ( .CLK(n5505), .C(n5506) );
  CKBD0 U5389 ( .CLK(n5506), .C(n5507) );
  CKBD0 U5390 ( .CLK(n5507), .C(n5508) );
  CKBD0 U5391 ( .CLK(n5508), .C(n5509) );
  CKBD0 U5392 ( .CLK(n5509), .C(n5510) );
  CKBD0 U5393 ( .CLK(n5510), .C(n5511) );
  BUFFD0 U5394 ( .I(n5511), .Z(n5512) );
  CKBD0 U5395 ( .CLK(n5512), .C(n5513) );
  CKBD0 U5396 ( .CLK(n5513), .C(n5514) );
  CKBD0 U5397 ( .CLK(n5514), .C(n5515) );
  CKBD0 U5398 ( .CLK(n5515), .C(n5516) );
  CKBD0 U5399 ( .CLK(n5516), .C(n5517) );
  CKBD0 U5400 ( .CLK(n5517), .C(n5518) );
  CKBD0 U5401 ( .CLK(n5518), .C(n5519) );
  CKBD0 U5402 ( .CLK(n5519), .C(n5520) );
  CKBD0 U5403 ( .CLK(n5520), .C(n5521) );
  CKBD0 U5404 ( .CLK(n5521), .C(n5522) );
  CKBD0 U5405 ( .CLK(n5522), .C(n5523) );
  BUFFD0 U5406 ( .I(n5523), .Z(n5524) );
  CKBD0 U5407 ( .CLK(n5524), .C(n5525) );
  CKBD0 U5408 ( .CLK(n5525), .C(n5526) );
  CKBD0 U5409 ( .CLK(n5526), .C(n5527) );
  CKBD0 U5410 ( .CLK(n5527), .C(n5528) );
  CKBD0 U5411 ( .CLK(n5528), .C(n5529) );
  CKBD0 U5412 ( .CLK(n5529), .C(n5530) );
  CKBD0 U5413 ( .CLK(n5530), .C(n5531) );
  CKBD0 U5414 ( .CLK(n5531), .C(n5532) );
  CKBD0 U5415 ( .CLK(n5532), .C(n5533) );
  BUFFD0 U5416 ( .I(n5533), .Z(n5534) );
  CKBD0 U5417 ( .CLK(n5534), .C(n5535) );
  CKBD0 U5418 ( .CLK(n5535), .C(n5536) );
  CKBD0 U5419 ( .CLK(n5536), .C(n5537) );
  CKBD0 U5420 ( .CLK(n5537), .C(n5538) );
  CKBD0 U5421 ( .CLK(n5538), .C(n5539) );
  CKBD0 U5422 ( .CLK(n5539), .C(n5540) );
  CKBD0 U5423 ( .CLK(n5540), .C(n5541) );
  CKBD0 U5424 ( .CLK(n5541), .C(n5542) );
  CKBD0 U5425 ( .CLK(n5542), .C(n5543) );
  CKBD0 U5426 ( .CLK(n5543), .C(n5544) );
  BUFFD0 U5427 ( .I(n5544), .Z(n5545) );
  CKBD0 U5428 ( .CLK(n5545), .C(n5546) );
  CKBD0 U5429 ( .CLK(n5546), .C(n5547) );
  CKBD0 U5430 ( .CLK(n5547), .C(n5548) );
  CKBD0 U5431 ( .CLK(n5548), .C(n5549) );
  CKBD0 U5432 ( .CLK(n5549), .C(n5550) );
  CKBD0 U5433 ( .CLK(n5550), .C(n5551) );
  CKBD0 U5434 ( .CLK(n5551), .C(n5552) );
  CKBD0 U5435 ( .CLK(n5552), .C(n5553) );
  CKBD0 U5436 ( .CLK(n5553), .C(n5554) );
  CKBD0 U5437 ( .CLK(n5554), .C(n5555) );
  BUFFD0 U5438 ( .I(n5555), .Z(n5556) );
  CKBD0 U5439 ( .CLK(n5556), .C(n5557) );
  CKBD0 U5440 ( .CLK(n5557), .C(n5558) );
  CKBD0 U5441 ( .CLK(n5558), .C(n5559) );
  CKBD0 U5442 ( .CLK(n5559), .C(n5560) );
  CKBD0 U5443 ( .CLK(n5560), .C(n5561) );
  CKBD0 U5444 ( .CLK(n5561), .C(n5562) );
  CKBD0 U5445 ( .CLK(n5562), .C(n5563) );
  CKBD0 U5446 ( .CLK(n5563), .C(n5564) );
  CKBD0 U5447 ( .CLK(n5564), .C(n5565) );
  CKBD0 U5448 ( .CLK(n5565), .C(n5566) );
  BUFFD0 U5449 ( .I(n5566), .Z(n5567) );
  CKBD0 U5450 ( .CLK(n5567), .C(n5568) );
  CKBD0 U5451 ( .CLK(n5568), .C(n5569) );
  CKBD0 U5452 ( .CLK(n5569), .C(n5570) );
  CKBD0 U5453 ( .CLK(n5570), .C(n5571) );
  CKBD0 U5454 ( .CLK(n5571), .C(n5572) );
  CKBD0 U5455 ( .CLK(n5572), .C(n5573) );
  CKBD0 U5456 ( .CLK(n5573), .C(n5574) );
  CKBD0 U5457 ( .CLK(n5574), .C(n5575) );
  CKBD0 U5458 ( .CLK(n5575), .C(n5576) );
  CKBD0 U5459 ( .CLK(n5576), .C(n5577) );
  BUFFD0 U5460 ( .I(n5577), .Z(n5578) );
  CKBD0 U5461 ( .CLK(n5578), .C(n5579) );
  CKBD0 U5462 ( .CLK(n5579), .C(n5580) );
  CKBD0 U5463 ( .CLK(n5580), .C(n5581) );
  CKBD0 U5464 ( .CLK(n5581), .C(n5582) );
  CKBD0 U5465 ( .CLK(n5582), .C(n5583) );
  BUFFD0 U5466 ( .I(n5583), .Z(n5584) );
  CKBD0 U5467 ( .CLK(n5584), .C(n5585) );
  BUFFD0 U5468 ( .I(n5585), .Z(n5586) );
  CKBD0 U5469 ( .CLK(n5586), .C(n5587) );
  BUFFD0 U5470 ( .I(n5587), .Z(n5588) );
  CKBD0 U5471 ( .CLK(n5588), .C(n5589) );
  BUFFD0 U5472 ( .I(n5589), .Z(n5590) );
  CKBD0 U5473 ( .CLK(n5590), .C(n5591) );
  BUFFD0 U5474 ( .I(n5591), .Z(n5592) );
  CKBD0 U5475 ( .CLK(n5592), .C(n5593) );
  BUFFD0 U5476 ( .I(n5593), .Z(n5594) );
  CKBD0 U5477 ( .CLK(n5594), .C(n5595) );
  BUFFD0 U5478 ( .I(n5595), .Z(n5596) );
  CKBD0 U5479 ( .CLK(n5596), .C(n5597) );
  BUFFD0 U5480 ( .I(n5597), .Z(n5598) );
  BUFFD0 U5481 ( .I(n5600), .Z(n5599) );
  BUFFD0 U5482 ( .I(n5601), .Z(n5600) );
  BUFFD0 U5483 ( .I(n9190), .Z(n5601) );
  CKBD0 U5484 ( .CLK(n1153), .C(n5602) );
  CKBD0 U5485 ( .CLK(n5602), .C(n5603) );
  CKBD0 U5486 ( .CLK(n5603), .C(n5604) );
  BUFFD0 U5487 ( .I(n5604), .Z(n5605) );
  CKBD0 U5488 ( .CLK(n5605), .C(n5606) );
  CKBD0 U5489 ( .CLK(n5606), .C(n5607) );
  CKBD0 U5490 ( .CLK(n5607), .C(n5608) );
  CKBD0 U5491 ( .CLK(n5608), .C(n5609) );
  CKBD0 U5492 ( .CLK(n5609), .C(n5610) );
  CKBD0 U5493 ( .CLK(n5610), .C(n5611) );
  CKBD0 U5494 ( .CLK(n5611), .C(n5612) );
  CKBD0 U5495 ( .CLK(n5612), .C(n5613) );
  CKBD0 U5496 ( .CLK(n5613), .C(n5614) );
  CKBD0 U5497 ( .CLK(n5614), .C(n5615) );
  BUFFD0 U5498 ( .I(n5615), .Z(n5616) );
  CKBD0 U5499 ( .CLK(n5616), .C(n5617) );
  CKBD0 U5500 ( .CLK(n5617), .C(n5618) );
  CKBD0 U5501 ( .CLK(n5618), .C(n5619) );
  CKBD0 U5502 ( .CLK(n5619), .C(n5620) );
  CKBD0 U5503 ( .CLK(n5620), .C(n5621) );
  CKBD0 U5504 ( .CLK(n5621), .C(n5622) );
  CKBD0 U5505 ( .CLK(n5622), .C(n5623) );
  CKBD0 U5506 ( .CLK(n5623), .C(n5624) );
  CKBD0 U5507 ( .CLK(n5624), .C(n5625) );
  CKBD0 U5508 ( .CLK(n5625), .C(n5626) );
  BUFFD0 U5509 ( .I(n5626), .Z(n5627) );
  CKBD0 U5510 ( .CLK(n5627), .C(n5628) );
  CKBD0 U5511 ( .CLK(n5628), .C(n5629) );
  CKBD0 U5512 ( .CLK(n5629), .C(n5630) );
  CKBD0 U5513 ( .CLK(n5630), .C(n5631) );
  CKBD0 U5514 ( .CLK(n5631), .C(n5632) );
  CKBD0 U5515 ( .CLK(n5632), .C(n5633) );
  CKBD0 U5516 ( .CLK(n5633), .C(n5634) );
  CKBD0 U5517 ( .CLK(n5634), .C(n5635) );
  CKBD0 U5518 ( .CLK(n5635), .C(n5636) );
  CKBD0 U5519 ( .CLK(n5636), .C(n5637) );
  BUFFD0 U5520 ( .I(n5637), .Z(n5638) );
  CKBD0 U5521 ( .CLK(n5638), .C(n5639) );
  CKBD0 U5522 ( .CLK(n5639), .C(n5640) );
  CKBD0 U5523 ( .CLK(n5640), .C(n5641) );
  CKBD0 U5524 ( .CLK(n5641), .C(n5642) );
  CKBD0 U5525 ( .CLK(n5642), .C(n5643) );
  CKBD0 U5526 ( .CLK(n5643), .C(n5644) );
  CKBD0 U5527 ( .CLK(n5644), .C(n5645) );
  CKBD0 U5528 ( .CLK(n5645), .C(n5646) );
  CKBD0 U5529 ( .CLK(n5646), .C(n5647) );
  CKBD0 U5530 ( .CLK(n5647), .C(n5648) );
  BUFFD0 U5531 ( .I(n5648), .Z(n5649) );
  CKBD0 U5532 ( .CLK(n5649), .C(n5650) );
  CKBD0 U5533 ( .CLK(n5650), .C(n5651) );
  CKBD0 U5534 ( .CLK(n5651), .C(n5652) );
  CKBD0 U5535 ( .CLK(n5652), .C(n5653) );
  CKBD0 U5536 ( .CLK(n5653), .C(n5654) );
  CKBD0 U5537 ( .CLK(n5654), .C(n5655) );
  CKBD0 U5538 ( .CLK(n5655), .C(n5656) );
  CKBD0 U5539 ( .CLK(n5656), .C(n5657) );
  CKBD0 U5540 ( .CLK(n5657), .C(n5658) );
  CKBD0 U5541 ( .CLK(n5658), .C(n5659) );
  BUFFD0 U5542 ( .I(n5659), .Z(n5660) );
  CKBD0 U5543 ( .CLK(n5660), .C(n5661) );
  CKBD0 U5544 ( .CLK(n5661), .C(n5662) );
  CKBD0 U5545 ( .CLK(n5662), .C(n5663) );
  CKBD0 U5546 ( .CLK(n5663), .C(n5664) );
  CKBD0 U5547 ( .CLK(n5664), .C(n5665) );
  CKBD0 U5548 ( .CLK(n5665), .C(n5666) );
  CKBD0 U5549 ( .CLK(n5666), .C(n5667) );
  CKBD0 U5550 ( .CLK(n5667), .C(n5668) );
  CKBD0 U5551 ( .CLK(n5668), .C(n5669) );
  BUFFD0 U5552 ( .I(n5669), .Z(n5670) );
  CKBD0 U5553 ( .CLK(n5670), .C(n5671) );
  CKBD0 U5554 ( .CLK(n5671), .C(n5672) );
  CKBD0 U5555 ( .CLK(n5672), .C(n5673) );
  CKBD0 U5556 ( .CLK(n5673), .C(n5674) );
  CKBD0 U5557 ( .CLK(n5674), .C(n5675) );
  CKBD0 U5558 ( .CLK(n5675), .C(n5676) );
  CKBD0 U5559 ( .CLK(n5676), .C(n5677) );
  CKBD0 U5560 ( .CLK(n5677), .C(n5678) );
  CKBD0 U5561 ( .CLK(n5678), .C(n5679) );
  CKBD0 U5562 ( .CLK(n5679), .C(n5680) );
  CKBD0 U5563 ( .CLK(n5680), .C(n5681) );
  BUFFD0 U5564 ( .I(n5681), .Z(n5682) );
  CKBD0 U5565 ( .CLK(n5682), .C(n5683) );
  CKBD0 U5566 ( .CLK(n5683), .C(n5684) );
  CKBD0 U5567 ( .CLK(n5684), .C(n5685) );
  CKBD0 U5568 ( .CLK(n5685), .C(n5686) );
  CKBD0 U5569 ( .CLK(n5686), .C(n5687) );
  CKBD0 U5570 ( .CLK(n5687), .C(n5688) );
  CKBD0 U5571 ( .CLK(n5688), .C(n5689) );
  CKBD0 U5572 ( .CLK(n5689), .C(n5690) );
  CKBD0 U5573 ( .CLK(n5690), .C(n5691) );
  BUFFD0 U5574 ( .I(n5691), .Z(n5692) );
  CKBD0 U5575 ( .CLK(n5692), .C(n5693) );
  CKBD0 U5576 ( .CLK(n5693), .C(n5694) );
  CKBD0 U5577 ( .CLK(n5694), .C(n5695) );
  CKBD0 U5578 ( .CLK(n5695), .C(n5696) );
  CKBD0 U5579 ( .CLK(n5696), .C(n5697) );
  CKBD0 U5580 ( .CLK(n5697), .C(n5698) );
  CKBD0 U5581 ( .CLK(n5698), .C(n5699) );
  CKBD0 U5582 ( .CLK(n5699), .C(n5700) );
  CKBD0 U5583 ( .CLK(n5700), .C(n5701) );
  BUFFD0 U5584 ( .I(n5701), .Z(n5702) );
  CKBD0 U5585 ( .CLK(n5702), .C(n5703) );
  CKBD0 U5586 ( .CLK(n5703), .C(n5704) );
  CKBD0 U5587 ( .CLK(n5704), .C(n5705) );
  CKBD0 U5588 ( .CLK(n5705), .C(n5706) );
  CKBD0 U5589 ( .CLK(n5706), .C(n5707) );
  CKBD0 U5590 ( .CLK(n5707), .C(n5708) );
  CKBD0 U5591 ( .CLK(n5708), .C(n5709) );
  CKBD0 U5592 ( .CLK(n5709), .C(n5710) );
  CKBD0 U5593 ( .CLK(n5710), .C(n5711) );
  CKBD0 U5594 ( .CLK(n5711), .C(n5712) );
  CKBD0 U5595 ( .CLK(n5712), .C(n5713) );
  BUFFD0 U5596 ( .I(n5713), .Z(n5714) );
  CKBD0 U5597 ( .CLK(n5714), .C(n5715) );
  CKBD0 U5598 ( .CLK(n5715), .C(n5716) );
  CKBD0 U5599 ( .CLK(n5716), .C(n5717) );
  CKBD0 U5600 ( .CLK(n5717), .C(n5718) );
  CKBD0 U5601 ( .CLK(n5718), .C(n5719) );
  BUFFD0 U5602 ( .I(n5719), .Z(n5720) );
  CKBD0 U5603 ( .CLK(n5720), .C(n5721) );
  BUFFD0 U5604 ( .I(n5721), .Z(n5722) );
  CKBD0 U5605 ( .CLK(n5722), .C(n5723) );
  BUFFD0 U5606 ( .I(n5723), .Z(n5724) );
  CKBD0 U5607 ( .CLK(n5724), .C(n5725) );
  BUFFD0 U5608 ( .I(n5725), .Z(n5726) );
  CKBD0 U5609 ( .CLK(n5726), .C(n5727) );
  BUFFD0 U5610 ( .I(n5727), .Z(n5728) );
  CKBD0 U5611 ( .CLK(n5728), .C(n5729) );
  BUFFD0 U5612 ( .I(n5729), .Z(n5730) );
  CKBD0 U5613 ( .CLK(n5730), .C(n5731) );
  BUFFD0 U5614 ( .I(n5731), .Z(n5732) );
  CKBD0 U5615 ( .CLK(n5732), .C(n5733) );
  BUFFD0 U5616 ( .I(n5733), .Z(n5734) );
  BUFFD0 U5617 ( .I(n5736), .Z(n5735) );
  BUFFD0 U5618 ( .I(n5737), .Z(n5736) );
  BUFFD0 U5619 ( .I(n9191), .Z(n5737) );
  CKBD0 U5620 ( .CLK(n1151), .C(n5738) );
  CKBD0 U5621 ( .CLK(n5738), .C(n5739) );
  CKBD0 U5622 ( .CLK(n5739), .C(n5740) );
  BUFFD0 U5623 ( .I(n5740), .Z(n5741) );
  CKBD0 U5624 ( .CLK(n5741), .C(n5742) );
  CKBD0 U5625 ( .CLK(n5742), .C(n5743) );
  CKBD0 U5626 ( .CLK(n5743), .C(n5744) );
  CKBD0 U5627 ( .CLK(n5744), .C(n5745) );
  CKBD0 U5628 ( .CLK(n5745), .C(n5746) );
  CKBD0 U5629 ( .CLK(n5746), .C(n5747) );
  CKBD0 U5630 ( .CLK(n5747), .C(n5748) );
  CKBD0 U5631 ( .CLK(n5748), .C(n5749) );
  CKBD0 U5632 ( .CLK(n5749), .C(n5750) );
  CKBD0 U5633 ( .CLK(n5750), .C(n5751) );
  CKBD0 U5634 ( .CLK(n5751), .C(n5752) );
  BUFFD0 U5635 ( .I(n5752), .Z(n5753) );
  CKBD0 U5636 ( .CLK(n5753), .C(n5754) );
  CKBD0 U5637 ( .CLK(n5754), .C(n5755) );
  CKBD0 U5638 ( .CLK(n5755), .C(n5756) );
  CKBD0 U5639 ( .CLK(n5756), .C(n5757) );
  CKBD0 U5640 ( .CLK(n5757), .C(n5758) );
  CKBD0 U5641 ( .CLK(n5758), .C(n5759) );
  CKBD0 U5642 ( .CLK(n5759), .C(n5760) );
  CKBD0 U5643 ( .CLK(n5760), .C(n5761) );
  CKBD0 U5644 ( .CLK(n5761), .C(n5762) );
  BUFFD0 U5645 ( .I(n5762), .Z(n5763) );
  CKBD0 U5646 ( .CLK(n5763), .C(n5764) );
  CKBD0 U5647 ( .CLK(n5764), .C(n5765) );
  CKBD0 U5648 ( .CLK(n5765), .C(n5766) );
  CKBD0 U5649 ( .CLK(n5766), .C(n5767) );
  CKBD0 U5650 ( .CLK(n5767), .C(n5768) );
  CKBD0 U5651 ( .CLK(n5768), .C(n5769) );
  CKBD0 U5652 ( .CLK(n5769), .C(n5770) );
  CKBD0 U5653 ( .CLK(n5770), .C(n5771) );
  CKBD0 U5654 ( .CLK(n5771), .C(n5772) );
  BUFFD0 U5655 ( .I(n5772), .Z(n5773) );
  CKBD0 U5656 ( .CLK(n5773), .C(n5774) );
  CKBD0 U5657 ( .CLK(n5774), .C(n5775) );
  CKBD0 U5658 ( .CLK(n5775), .C(n5776) );
  CKBD0 U5659 ( .CLK(n5776), .C(n5777) );
  CKBD0 U5660 ( .CLK(n5777), .C(n5778) );
  CKBD0 U5661 ( .CLK(n5778), .C(n5779) );
  CKBD0 U5662 ( .CLK(n5779), .C(n5780) );
  CKBD0 U5663 ( .CLK(n5780), .C(n5781) );
  CKBD0 U5664 ( .CLK(n5781), .C(n5782) );
  CKBD0 U5665 ( .CLK(n5782), .C(n5783) );
  CKBD0 U5666 ( .CLK(n5783), .C(n5784) );
  BUFFD0 U5667 ( .I(n5784), .Z(n5785) );
  CKBD0 U5668 ( .CLK(n5785), .C(n5786) );
  CKBD0 U5669 ( .CLK(n5786), .C(n5787) );
  CKBD0 U5670 ( .CLK(n5787), .C(n5788) );
  CKBD0 U5671 ( .CLK(n5788), .C(n5789) );
  CKBD0 U5672 ( .CLK(n5789), .C(n5790) );
  CKBD0 U5673 ( .CLK(n5790), .C(n5791) );
  CKBD0 U5674 ( .CLK(n5791), .C(n5792) );
  CKBD0 U5675 ( .CLK(n5792), .C(n5793) );
  CKBD0 U5676 ( .CLK(n5793), .C(n5794) );
  BUFFD0 U5677 ( .I(n5794), .Z(n5795) );
  CKBD0 U5678 ( .CLK(n5795), .C(n5796) );
  CKBD0 U5679 ( .CLK(n5796), .C(n5797) );
  CKBD0 U5680 ( .CLK(n5797), .C(n5798) );
  CKBD0 U5681 ( .CLK(n5798), .C(n5799) );
  CKBD0 U5682 ( .CLK(n5799), .C(n5800) );
  CKBD0 U5683 ( .CLK(n5800), .C(n5801) );
  CKBD0 U5684 ( .CLK(n5801), .C(n5802) );
  CKBD0 U5685 ( .CLK(n5802), .C(n5803) );
  CKBD0 U5686 ( .CLK(n5803), .C(n5804) );
  CKBD0 U5687 ( .CLK(n5804), .C(n5805) );
  BUFFD0 U5688 ( .I(n5805), .Z(n5806) );
  CKBD0 U5689 ( .CLK(n5806), .C(n5807) );
  CKBD0 U5690 ( .CLK(n5807), .C(n5808) );
  CKBD0 U5691 ( .CLK(n5808), .C(n5809) );
  CKBD0 U5692 ( .CLK(n5809), .C(n5810) );
  CKBD0 U5693 ( .CLK(n5810), .C(n5811) );
  CKBD0 U5694 ( .CLK(n5811), .C(n5812) );
  CKBD0 U5695 ( .CLK(n5812), .C(n5813) );
  CKBD0 U5696 ( .CLK(n5813), .C(n5814) );
  CKBD0 U5697 ( .CLK(n5814), .C(n5815) );
  CKBD0 U5698 ( .CLK(n5815), .C(n5816) );
  BUFFD0 U5699 ( .I(n5816), .Z(n5817) );
  CKBD0 U5700 ( .CLK(n5817), .C(n5818) );
  CKBD0 U5701 ( .CLK(n5818), .C(n5819) );
  CKBD0 U5702 ( .CLK(n5819), .C(n5820) );
  CKBD0 U5703 ( .CLK(n5820), .C(n5821) );
  CKBD0 U5704 ( .CLK(n5821), .C(n5822) );
  CKBD0 U5705 ( .CLK(n5822), .C(n5823) );
  CKBD0 U5706 ( .CLK(n5823), .C(n5824) );
  CKBD0 U5707 ( .CLK(n5824), .C(n5825) );
  CKBD0 U5708 ( .CLK(n5825), .C(n5826) );
  CKBD0 U5709 ( .CLK(n5826), .C(n5827) );
  BUFFD0 U5710 ( .I(n5827), .Z(n5828) );
  CKBD0 U5711 ( .CLK(n5828), .C(n5829) );
  CKBD0 U5712 ( .CLK(n5829), .C(n5830) );
  CKBD0 U5713 ( .CLK(n5830), .C(n5831) );
  CKBD0 U5714 ( .CLK(n5831), .C(n5832) );
  CKBD0 U5715 ( .CLK(n5832), .C(n5833) );
  CKBD0 U5716 ( .CLK(n5833), .C(n5834) );
  CKBD0 U5717 ( .CLK(n5834), .C(n5835) );
  CKBD0 U5718 ( .CLK(n5835), .C(n5836) );
  CKBD0 U5719 ( .CLK(n5836), .C(n5837) );
  BUFFD0 U5720 ( .I(n5837), .Z(n5838) );
  CKBD0 U5721 ( .CLK(n5838), .C(n5839) );
  CKBD0 U5722 ( .CLK(n5839), .C(n5840) );
  CKBD0 U5723 ( .CLK(n5840), .C(n5841) );
  CKBD0 U5724 ( .CLK(n5841), .C(n5842) );
  CKBD0 U5725 ( .CLK(n5842), .C(n5843) );
  CKBD0 U5726 ( .CLK(n5843), .C(n5844) );
  CKBD0 U5727 ( .CLK(n5844), .C(n5845) );
  CKBD0 U5728 ( .CLK(n5845), .C(n5846) );
  CKBD0 U5729 ( .CLK(n5846), .C(n5847) );
  CKBD0 U5730 ( .CLK(n5847), .C(n5848) );
  CKBD0 U5731 ( .CLK(n5848), .C(n5849) );
  BUFFD0 U5732 ( .I(n5849), .Z(n5850) );
  CKBD0 U5733 ( .CLK(n5850), .C(n5851) );
  CKBD0 U5734 ( .CLK(n5851), .C(n5852) );
  CKBD0 U5735 ( .CLK(n5852), .C(n5853) );
  CKBD0 U5736 ( .CLK(n5853), .C(n5854) );
  CKBD0 U5737 ( .CLK(n5854), .C(n5855) );
  BUFFD0 U5738 ( .I(n5855), .Z(n5856) );
  CKBD0 U5739 ( .CLK(n5856), .C(n5857) );
  BUFFD0 U5740 ( .I(n5857), .Z(n5858) );
  CKBD0 U5741 ( .CLK(n5858), .C(n5859) );
  BUFFD0 U5742 ( .I(n5859), .Z(n5860) );
  CKBD0 U5743 ( .CLK(n5860), .C(n5861) );
  BUFFD0 U5744 ( .I(n5861), .Z(n5862) );
  CKBD0 U5745 ( .CLK(n5862), .C(n5863) );
  BUFFD0 U5746 ( .I(n5863), .Z(n5864) );
  CKBD0 U5747 ( .CLK(n5864), .C(n5865) );
  BUFFD0 U5748 ( .I(n5865), .Z(n5866) );
  CKBD0 U5749 ( .CLK(n5866), .C(n5867) );
  BUFFD0 U5750 ( .I(n5867), .Z(n5868) );
  CKBD0 U5751 ( .CLK(n5868), .C(n5869) );
  BUFFD0 U5752 ( .I(n5869), .Z(n5870) );
  BUFFD0 U5753 ( .I(n5872), .Z(n5871) );
  BUFFD0 U5754 ( .I(n5873), .Z(n5872) );
  BUFFD0 U5755 ( .I(n9192), .Z(n5873) );
  CKBD0 U5756 ( .CLK(n2605), .C(n5874) );
  CKBD0 U5757 ( .CLK(n5874), .C(n5875) );
  CKBD0 U5758 ( .CLK(n5875), .C(n5876) );
  BUFFD0 U5759 ( .I(n5876), .Z(n5877) );
  CKBD0 U5760 ( .CLK(n5877), .C(n5878) );
  CKBD0 U5761 ( .CLK(n5878), .C(n5879) );
  CKBD0 U5762 ( .CLK(n5879), .C(n5880) );
  CKBD0 U5763 ( .CLK(n5880), .C(n5881) );
  CKBD0 U5764 ( .CLK(n5881), .C(n5882) );
  CKBD0 U5765 ( .CLK(n5882), .C(n5883) );
  CKBD0 U5766 ( .CLK(n5883), .C(n5884) );
  CKBD0 U5767 ( .CLK(n5884), .C(n5885) );
  CKBD0 U5768 ( .CLK(n5885), .C(n5886) );
  CKBD0 U5769 ( .CLK(n5886), .C(n5887) );
  BUFFD0 U5770 ( .I(n5887), .Z(n5888) );
  CKBD0 U5771 ( .CLK(n5888), .C(n5889) );
  CKBD0 U5772 ( .CLK(n5889), .C(n5890) );
  CKBD0 U5773 ( .CLK(n5890), .C(n5891) );
  CKBD0 U5774 ( .CLK(n5891), .C(n5892) );
  CKBD0 U5775 ( .CLK(n5892), .C(n5893) );
  CKBD0 U5776 ( .CLK(n5893), .C(n5894) );
  CKBD0 U5777 ( .CLK(n5894), .C(n5895) );
  CKBD0 U5778 ( .CLK(n5895), .C(n5896) );
  CKBD0 U5779 ( .CLK(n5896), .C(n5897) );
  CKBD0 U5780 ( .CLK(n5897), .C(n5898) );
  BUFFD0 U5781 ( .I(n5898), .Z(n5899) );
  CKBD0 U5782 ( .CLK(n5899), .C(n5900) );
  CKBD0 U5783 ( .CLK(n5900), .C(n5901) );
  CKBD0 U5784 ( .CLK(n5901), .C(n5902) );
  CKBD0 U5785 ( .CLK(n5902), .C(n5903) );
  CKBD0 U5786 ( .CLK(n5903), .C(n5904) );
  CKBD0 U5787 ( .CLK(n5904), .C(n5905) );
  CKBD0 U5788 ( .CLK(n5905), .C(n5906) );
  CKBD0 U5789 ( .CLK(n5906), .C(n5907) );
  CKBD0 U5790 ( .CLK(n5907), .C(n5908) );
  BUFFD0 U5791 ( .I(n5908), .Z(n5909) );
  CKBD0 U5792 ( .CLK(n5909), .C(n5910) );
  CKBD0 U5793 ( .CLK(n5910), .C(n5911) );
  CKBD0 U5794 ( .CLK(n5911), .C(n5912) );
  CKBD0 U5795 ( .CLK(n5912), .C(n5913) );
  CKBD0 U5796 ( .CLK(n5913), .C(n5914) );
  CKBD0 U5797 ( .CLK(n5914), .C(n5915) );
  CKBD0 U5798 ( .CLK(n5915), .C(n5916) );
  CKBD0 U5799 ( .CLK(n5916), .C(n5917) );
  CKBD0 U5800 ( .CLK(n5917), .C(n5918) );
  CKBD0 U5801 ( .CLK(n5918), .C(n5919) );
  CKBD0 U5802 ( .CLK(n5919), .C(n5920) );
  BUFFD0 U5803 ( .I(n5920), .Z(n5921) );
  CKBD0 U5804 ( .CLK(n5921), .C(n5922) );
  CKBD0 U5805 ( .CLK(n5922), .C(n5923) );
  CKBD0 U5806 ( .CLK(n5923), .C(n5924) );
  CKBD0 U5807 ( .CLK(n5924), .C(n5925) );
  CKBD0 U5808 ( .CLK(n5925), .C(n5926) );
  CKBD0 U5809 ( .CLK(n5926), .C(n5927) );
  CKBD0 U5810 ( .CLK(n5927), .C(n5928) );
  CKBD0 U5811 ( .CLK(n5928), .C(n5929) );
  CKBD0 U5812 ( .CLK(n5929), .C(n5930) );
  BUFFD0 U5813 ( .I(n5930), .Z(n5931) );
  CKBD0 U5814 ( .CLK(n5931), .C(n5932) );
  CKBD0 U5815 ( .CLK(n5932), .C(n5933) );
  CKBD0 U5816 ( .CLK(n5933), .C(n5934) );
  CKBD0 U5817 ( .CLK(n5934), .C(n5935) );
  CKBD0 U5818 ( .CLK(n5935), .C(n5936) );
  CKBD0 U5819 ( .CLK(n5936), .C(n5937) );
  CKBD0 U5820 ( .CLK(n5937), .C(n5938) );
  CKBD0 U5821 ( .CLK(n5938), .C(n5939) );
  CKBD0 U5822 ( .CLK(n5939), .C(n5940) );
  CKBD0 U5823 ( .CLK(n5940), .C(n5941) );
  CKBD0 U5824 ( .CLK(n5941), .C(n5942) );
  BUFFD0 U5825 ( .I(n5942), .Z(n5943) );
  CKBD0 U5826 ( .CLK(n5943), .C(n5944) );
  CKBD0 U5827 ( .CLK(n5944), .C(n5945) );
  CKBD0 U5828 ( .CLK(n5945), .C(n5946) );
  CKBD0 U5829 ( .CLK(n5946), .C(n5947) );
  CKBD0 U5830 ( .CLK(n5947), .C(n5948) );
  CKBD0 U5831 ( .CLK(n5948), .C(n5949) );
  CKBD0 U5832 ( .CLK(n5949), .C(n5950) );
  CKBD0 U5833 ( .CLK(n5950), .C(n5951) );
  CKBD0 U5834 ( .CLK(n5951), .C(n5952) );
  BUFFD0 U5835 ( .I(n5952), .Z(n5953) );
  CKBD0 U5836 ( .CLK(n5953), .C(n5954) );
  CKBD0 U5837 ( .CLK(n5954), .C(n5955) );
  CKBD0 U5838 ( .CLK(n5955), .C(n5956) );
  CKBD0 U5839 ( .CLK(n5956), .C(n5957) );
  CKBD0 U5840 ( .CLK(n5957), .C(n5958) );
  CKBD0 U5841 ( .CLK(n5958), .C(n5959) );
  CKBD0 U5842 ( .CLK(n5959), .C(n5960) );
  CKBD0 U5843 ( .CLK(n5960), .C(n5961) );
  CKBD0 U5844 ( .CLK(n5961), .C(n5962) );
  CKBD0 U5845 ( .CLK(n5962), .C(n5963) );
  BUFFD0 U5846 ( .I(n5963), .Z(n5964) );
  CKBD0 U5847 ( .CLK(n5964), .C(n5965) );
  CKBD0 U5848 ( .CLK(n5965), .C(n5966) );
  CKBD0 U5849 ( .CLK(n5966), .C(n5967) );
  CKBD0 U5850 ( .CLK(n5967), .C(n5968) );
  CKBD0 U5851 ( .CLK(n5968), .C(n5969) );
  CKBD0 U5852 ( .CLK(n5969), .C(n5970) );
  CKBD0 U5853 ( .CLK(n5970), .C(n5971) );
  CKBD0 U5854 ( .CLK(n5971), .C(n5972) );
  CKBD0 U5855 ( .CLK(n5972), .C(n5973) );
  CKBD0 U5856 ( .CLK(n5973), .C(n5974) );
  BUFFD0 U5857 ( .I(n5974), .Z(n5975) );
  CKBD0 U5858 ( .CLK(n5975), .C(n5976) );
  CKBD0 U5859 ( .CLK(n5976), .C(n5977) );
  CKBD0 U5860 ( .CLK(n5977), .C(n5978) );
  CKBD0 U5861 ( .CLK(n5978), .C(n5979) );
  CKBD0 U5862 ( .CLK(n5979), .C(n5980) );
  CKBD0 U5863 ( .CLK(n5980), .C(n5981) );
  CKBD0 U5864 ( .CLK(n5981), .C(n5982) );
  CKBD0 U5865 ( .CLK(n5982), .C(n5983) );
  CKBD0 U5866 ( .CLK(n5983), .C(n5984) );
  CKBD0 U5867 ( .CLK(n5984), .C(n5985) );
  BUFFD0 U5868 ( .I(n5985), .Z(n5986) );
  CKBD0 U5869 ( .CLK(n5986), .C(n5987) );
  CKBD0 U5870 ( .CLK(n5987), .C(n5988) );
  CKBD0 U5871 ( .CLK(n5988), .C(n5989) );
  CKBD0 U5872 ( .CLK(n5989), .C(n5990) );
  CKBD0 U5873 ( .CLK(n5990), .C(n5991) );
  BUFFD0 U5874 ( .I(n5991), .Z(n5992) );
  CKBD0 U5875 ( .CLK(n5992), .C(n5993) );
  BUFFD0 U5876 ( .I(n5993), .Z(n5994) );
  CKBD0 U5877 ( .CLK(n5994), .C(n5995) );
  BUFFD0 U5878 ( .I(n5995), .Z(n5996) );
  CKBD0 U5879 ( .CLK(n5996), .C(n5997) );
  BUFFD0 U5880 ( .I(n5997), .Z(n5998) );
  CKBD0 U5881 ( .CLK(n5998), .C(n5999) );
  BUFFD0 U5882 ( .I(n5999), .Z(n6000) );
  CKBD0 U5883 ( .CLK(n6000), .C(n6001) );
  BUFFD0 U5884 ( .I(n6001), .Z(n6002) );
  CKBD0 U5885 ( .CLK(n6002), .C(n6003) );
  BUFFD0 U5886 ( .I(n6003), .Z(n6004) );
  CKBD0 U5887 ( .CLK(n6004), .C(n6005) );
  BUFFD0 U5888 ( .I(n6005), .Z(n6006) );
  BUFFD0 U5889 ( .I(n6008), .Z(n6007) );
  BUFFD0 U5890 ( .I(n6009), .Z(n6008) );
  BUFFD0 U5891 ( .I(n6010), .Z(n6009) );
  BUFFD0 U5892 ( .I(n9193), .Z(n6010) );
  CKBD0 U5893 ( .CLK(n950), .C(n6011) );
  CKBD0 U5894 ( .CLK(n6011), .C(n6012) );
  CKBD0 U5895 ( .CLK(n6012), .C(n6013) );
  BUFFD0 U5896 ( .I(n6013), .Z(n6014) );
  CKBD0 U5897 ( .CLK(n6014), .C(n6015) );
  CKBD0 U5898 ( .CLK(n6015), .C(n6016) );
  CKBD0 U5899 ( .CLK(n6016), .C(n6017) );
  CKBD0 U5900 ( .CLK(n6017), .C(n6018) );
  CKBD0 U5901 ( .CLK(n6018), .C(n6019) );
  CKBD0 U5902 ( .CLK(n6019), .C(n6020) );
  CKBD0 U5903 ( .CLK(n6020), .C(n6021) );
  CKBD0 U5904 ( .CLK(n6021), .C(n6022) );
  CKBD0 U5905 ( .CLK(n6022), .C(n6023) );
  CKBD0 U5906 ( .CLK(n6023), .C(n6024) );
  BUFFD0 U5907 ( .I(n6024), .Z(n6025) );
  CKBD0 U5908 ( .CLK(n6025), .C(n6026) );
  CKBD0 U5909 ( .CLK(n6026), .C(n6027) );
  CKBD0 U5910 ( .CLK(n6027), .C(n6028) );
  CKBD0 U5911 ( .CLK(n6028), .C(n6029) );
  CKBD0 U5912 ( .CLK(n6029), .C(n6030) );
  CKBD0 U5913 ( .CLK(n6030), .C(n6031) );
  CKBD0 U5914 ( .CLK(n6031), .C(n6032) );
  CKBD0 U5915 ( .CLK(n6032), .C(n6033) );
  CKBD0 U5916 ( .CLK(n6033), .C(n6034) );
  CKBD0 U5917 ( .CLK(n6034), .C(n6035) );
  BUFFD0 U5918 ( .I(n6035), .Z(n6036) );
  CKBD0 U5919 ( .CLK(n6036), .C(n6037) );
  CKBD0 U5920 ( .CLK(n6037), .C(n6038) );
  CKBD0 U5921 ( .CLK(n6038), .C(n6039) );
  CKBD0 U5922 ( .CLK(n6039), .C(n6040) );
  CKBD0 U5923 ( .CLK(n6040), .C(n6041) );
  CKBD0 U5924 ( .CLK(n6041), .C(n6042) );
  CKBD0 U5925 ( .CLK(n6042), .C(n6043) );
  CKBD0 U5926 ( .CLK(n6043), .C(n6044) );
  CKBD0 U5927 ( .CLK(n6044), .C(n6045) );
  BUFFD0 U5928 ( .I(n6045), .Z(n6046) );
  CKBD0 U5929 ( .CLK(n6046), .C(n6047) );
  CKBD0 U5930 ( .CLK(n6047), .C(n6048) );
  CKBD0 U5931 ( .CLK(n6048), .C(n6049) );
  CKBD0 U5932 ( .CLK(n6049), .C(n6050) );
  CKBD0 U5933 ( .CLK(n6050), .C(n6051) );
  CKBD0 U5934 ( .CLK(n6051), .C(n6052) );
  CKBD0 U5935 ( .CLK(n6052), .C(n6053) );
  CKBD0 U5936 ( .CLK(n6053), .C(n6054) );
  CKBD0 U5937 ( .CLK(n6054), .C(n6055) );
  CKBD0 U5938 ( .CLK(n6055), .C(n6056) );
  CKBD0 U5939 ( .CLK(n6056), .C(n6057) );
  BUFFD0 U5940 ( .I(n6057), .Z(n6058) );
  CKBD0 U5941 ( .CLK(n6058), .C(n6059) );
  CKBD0 U5942 ( .CLK(n6059), .C(n6060) );
  CKBD0 U5943 ( .CLK(n6060), .C(n6061) );
  CKBD0 U5944 ( .CLK(n6061), .C(n6062) );
  CKBD0 U5945 ( .CLK(n6062), .C(n6063) );
  CKBD0 U5946 ( .CLK(n6063), .C(n6064) );
  CKBD0 U5947 ( .CLK(n6064), .C(n6065) );
  CKBD0 U5948 ( .CLK(n6065), .C(n6066) );
  CKBD0 U5949 ( .CLK(n6066), .C(n6067) );
  BUFFD0 U5950 ( .I(n6067), .Z(n6068) );
  CKBD0 U5951 ( .CLK(n6068), .C(n6069) );
  CKBD0 U5952 ( .CLK(n6069), .C(n6070) );
  CKBD0 U5953 ( .CLK(n6070), .C(n6071) );
  CKBD0 U5954 ( .CLK(n6071), .C(n6072) );
  CKBD0 U5955 ( .CLK(n6072), .C(n6073) );
  CKBD0 U5956 ( .CLK(n6073), .C(n6074) );
  CKBD0 U5957 ( .CLK(n6074), .C(n6075) );
  CKBD0 U5958 ( .CLK(n6075), .C(n6076) );
  CKBD0 U5959 ( .CLK(n6076), .C(n6077) );
  CKBD0 U5960 ( .CLK(n6077), .C(n6078) );
  BUFFD0 U5961 ( .I(n6078), .Z(n6079) );
  CKBD0 U5962 ( .CLK(n6079), .C(n6080) );
  CKBD0 U5963 ( .CLK(n6080), .C(n6081) );
  CKBD0 U5964 ( .CLK(n6081), .C(n6082) );
  CKBD0 U5965 ( .CLK(n6082), .C(n6083) );
  CKBD0 U5966 ( .CLK(n6083), .C(n6084) );
  CKBD0 U5967 ( .CLK(n6084), .C(n6085) );
  CKBD0 U5968 ( .CLK(n6085), .C(n6086) );
  CKBD0 U5969 ( .CLK(n6086), .C(n6087) );
  CKBD0 U5970 ( .CLK(n6087), .C(n6088) );
  CKBD0 U5971 ( .CLK(n6088), .C(n6089) );
  BUFFD0 U5972 ( .I(n6089), .Z(n6090) );
  CKBD0 U5973 ( .CLK(n6090), .C(n6091) );
  CKBD0 U5974 ( .CLK(n6091), .C(n6092) );
  CKBD0 U5975 ( .CLK(n6092), .C(n6093) );
  CKBD0 U5976 ( .CLK(n6093), .C(n6094) );
  CKBD0 U5977 ( .CLK(n6094), .C(n6095) );
  CKBD0 U5978 ( .CLK(n6095), .C(n6096) );
  CKBD0 U5979 ( .CLK(n6096), .C(n6097) );
  CKBD0 U5980 ( .CLK(n6097), .C(n6098) );
  CKBD0 U5981 ( .CLK(n6098), .C(n6099) );
  CKBD0 U5982 ( .CLK(n6099), .C(n6100) );
  BUFFD0 U5983 ( .I(n6100), .Z(n6101) );
  CKBD0 U5984 ( .CLK(n6101), .C(n6102) );
  CKBD0 U5985 ( .CLK(n6102), .C(n6103) );
  CKBD0 U5986 ( .CLK(n6103), .C(n6104) );
  CKBD0 U5987 ( .CLK(n6104), .C(n6105) );
  CKBD0 U5988 ( .CLK(n6105), .C(n6106) );
  CKBD0 U5989 ( .CLK(n6106), .C(n6107) );
  CKBD0 U5990 ( .CLK(n6107), .C(n6108) );
  CKBD0 U5991 ( .CLK(n6108), .C(n6109) );
  CKBD0 U5992 ( .CLK(n6109), .C(n6110) );
  CKBD0 U5993 ( .CLK(n6110), .C(n6111) );
  BUFFD0 U5994 ( .I(n6111), .Z(n6112) );
  CKBD0 U5995 ( .CLK(n6112), .C(n6113) );
  CKBD0 U5996 ( .CLK(n6113), .C(n6114) );
  CKBD0 U5997 ( .CLK(n6114), .C(n6115) );
  CKBD0 U5998 ( .CLK(n6115), .C(n6116) );
  CKBD0 U5999 ( .CLK(n6116), .C(n6117) );
  CKBD0 U6000 ( .CLK(n6117), .C(n6118) );
  CKBD0 U6001 ( .CLK(n6118), .C(n6119) );
  CKBD0 U6002 ( .CLK(n6119), .C(n6120) );
  CKBD0 U6003 ( .CLK(n6120), .C(n6121) );
  CKBD0 U6004 ( .CLK(n6121), .C(n6122) );
  BUFFD0 U6005 ( .I(n6122), .Z(n6123) );
  CKBD0 U6006 ( .CLK(n6123), .C(n6124) );
  CKBD0 U6007 ( .CLK(n6124), .C(n6125) );
  CKBD0 U6008 ( .CLK(n6125), .C(n6126) );
  CKBD0 U6009 ( .CLK(n6126), .C(n6127) );
  CKBD0 U6010 ( .CLK(n6127), .C(n6128) );
  BUFFD0 U6011 ( .I(n6128), .Z(n6129) );
  CKBD0 U6012 ( .CLK(n6129), .C(n6130) );
  BUFFD0 U6013 ( .I(n6130), .Z(n6131) );
  CKBD0 U6014 ( .CLK(n6131), .C(n6132) );
  BUFFD0 U6015 ( .I(n6132), .Z(n6133) );
  CKBD0 U6016 ( .CLK(n6133), .C(n6134) );
  BUFFD0 U6017 ( .I(n6134), .Z(n6135) );
  CKBD0 U6018 ( .CLK(n6135), .C(n6136) );
  BUFFD0 U6019 ( .I(n6136), .Z(n6137) );
  CKBD0 U6020 ( .CLK(n6137), .C(n6138) );
  BUFFD0 U6021 ( .I(n6138), .Z(n6139) );
  CKBD0 U6022 ( .CLK(n6139), .C(n6140) );
  BUFFD0 U6023 ( .I(n6140), .Z(n6141) );
  CKBD0 U6024 ( .CLK(n6141), .C(n6142) );
  BUFFD0 U6025 ( .I(n6142), .Z(n6143) );
  BUFFD0 U6026 ( .I(n9194), .Z(n6144) );
  BUFFD0 U6027 ( .I(n6146), .Z(n6145) );
  BUFFD0 U6028 ( .I(n6147), .Z(n6146) );
  BUFFD0 U6029 ( .I(Decoder[5]), .Z(n6147) );
  CKBD0 U6030 ( .CLK(n948), .C(n6148) );
  CKBD0 U6031 ( .CLK(n6148), .C(n6149) );
  CKBD0 U6032 ( .CLK(n6149), .C(n6150) );
  BUFFD0 U6033 ( .I(n6150), .Z(n6151) );
  CKBD0 U6034 ( .CLK(n6151), .C(n6152) );
  CKBD0 U6035 ( .CLK(n6152), .C(n6153) );
  CKBD0 U6036 ( .CLK(n6153), .C(n6154) );
  CKBD0 U6037 ( .CLK(n6154), .C(n6155) );
  CKBD0 U6038 ( .CLK(n6155), .C(n6156) );
  CKBD0 U6039 ( .CLK(n6156), .C(n6157) );
  CKBD0 U6040 ( .CLK(n6157), .C(n6158) );
  CKBD0 U6041 ( .CLK(n6158), .C(n6159) );
  CKBD0 U6042 ( .CLK(n6159), .C(n6160) );
  CKBD0 U6043 ( .CLK(n6160), .C(n6161) );
  BUFFD0 U6044 ( .I(n6161), .Z(n6162) );
  CKBD0 U6045 ( .CLK(n6162), .C(n6163) );
  CKBD0 U6046 ( .CLK(n6163), .C(n6164) );
  CKBD0 U6047 ( .CLK(n6164), .C(n6165) );
  CKBD0 U6048 ( .CLK(n6165), .C(n6166) );
  CKBD0 U6049 ( .CLK(n6166), .C(n6167) );
  CKBD0 U6050 ( .CLK(n6167), .C(n6168) );
  CKBD0 U6051 ( .CLK(n6168), .C(n6169) );
  CKBD0 U6052 ( .CLK(n6169), .C(n6170) );
  CKBD0 U6053 ( .CLK(n6170), .C(n6171) );
  CKBD0 U6054 ( .CLK(n6171), .C(n6172) );
  BUFFD0 U6055 ( .I(n6172), .Z(n6173) );
  CKBD0 U6056 ( .CLK(n6173), .C(n6174) );
  CKBD0 U6057 ( .CLK(n6174), .C(n6175) );
  CKBD0 U6058 ( .CLK(n6175), .C(n6176) );
  CKBD0 U6059 ( .CLK(n6176), .C(n6177) );
  CKBD0 U6060 ( .CLK(n6177), .C(n6178) );
  CKBD0 U6061 ( .CLK(n6178), .C(n6179) );
  CKBD0 U6062 ( .CLK(n6179), .C(n6180) );
  CKBD0 U6063 ( .CLK(n6180), .C(n6181) );
  CKBD0 U6064 ( .CLK(n6181), .C(n6182) );
  CKBD0 U6065 ( .CLK(n6182), .C(n6183) );
  BUFFD0 U6066 ( .I(n6183), .Z(n6184) );
  CKBD0 U6067 ( .CLK(n6184), .C(n6185) );
  CKBD0 U6068 ( .CLK(n6185), .C(n6186) );
  CKBD0 U6069 ( .CLK(n6186), .C(n6187) );
  CKBD0 U6070 ( .CLK(n6187), .C(n6188) );
  CKBD0 U6071 ( .CLK(n6188), .C(n6189) );
  CKBD0 U6072 ( .CLK(n6189), .C(n6190) );
  CKBD0 U6073 ( .CLK(n6190), .C(n6191) );
  CKBD0 U6074 ( .CLK(n6191), .C(n6192) );
  CKBD0 U6075 ( .CLK(n6192), .C(n6193) );
  BUFFD0 U6076 ( .I(n6193), .Z(n6194) );
  CKBD0 U6077 ( .CLK(n6194), .C(n6195) );
  CKBD0 U6078 ( .CLK(n6195), .C(n6196) );
  CKBD0 U6079 ( .CLK(n6196), .C(n6197) );
  CKBD0 U6080 ( .CLK(n6197), .C(n6198) );
  CKBD0 U6081 ( .CLK(n6198), .C(n6199) );
  CKBD0 U6082 ( .CLK(n6199), .C(n6200) );
  CKBD0 U6083 ( .CLK(n6200), .C(n6201) );
  CKBD0 U6084 ( .CLK(n6201), .C(n6202) );
  CKBD0 U6085 ( .CLK(n6202), .C(n6203) );
  CKBD0 U6086 ( .CLK(n6203), .C(n6204) );
  CKBD0 U6087 ( .CLK(n6204), .C(n6205) );
  BUFFD0 U6088 ( .I(n6205), .Z(n6206) );
  CKBD0 U6089 ( .CLK(n6206), .C(n6207) );
  CKBD0 U6090 ( .CLK(n6207), .C(n6208) );
  CKBD0 U6091 ( .CLK(n6208), .C(n6209) );
  CKBD0 U6092 ( .CLK(n6209), .C(n6210) );
  CKBD0 U6093 ( .CLK(n6210), .C(n6211) );
  CKBD0 U6094 ( .CLK(n6211), .C(n6212) );
  CKBD0 U6095 ( .CLK(n6212), .C(n6213) );
  CKBD0 U6096 ( .CLK(n6213), .C(n6214) );
  CKBD0 U6097 ( .CLK(n6214), .C(n6215) );
  BUFFD0 U6098 ( .I(n6215), .Z(n6216) );
  CKBD0 U6099 ( .CLK(n6216), .C(n6217) );
  CKBD0 U6100 ( .CLK(n6217), .C(n6218) );
  CKBD0 U6101 ( .CLK(n6218), .C(n6219) );
  CKBD0 U6102 ( .CLK(n6219), .C(n6220) );
  CKBD0 U6103 ( .CLK(n6220), .C(n6221) );
  CKBD0 U6104 ( .CLK(n6221), .C(n6222) );
  CKBD0 U6105 ( .CLK(n6222), .C(n6223) );
  CKBD0 U6106 ( .CLK(n6223), .C(n6224) );
  CKBD0 U6107 ( .CLK(n6224), .C(n6225) );
  CKBD0 U6108 ( .CLK(n6225), .C(n6226) );
  BUFFD0 U6109 ( .I(n6226), .Z(n6227) );
  CKBD0 U6110 ( .CLK(n6227), .C(n6228) );
  CKBD0 U6111 ( .CLK(n6228), .C(n6229) );
  CKBD0 U6112 ( .CLK(n6229), .C(n6230) );
  CKBD0 U6113 ( .CLK(n6230), .C(n6231) );
  CKBD0 U6114 ( .CLK(n6231), .C(n6232) );
  CKBD0 U6115 ( .CLK(n6232), .C(n6233) );
  CKBD0 U6116 ( .CLK(n6233), .C(n6234) );
  CKBD0 U6117 ( .CLK(n6234), .C(n6235) );
  CKBD0 U6118 ( .CLK(n6235), .C(n6236) );
  CKBD0 U6119 ( .CLK(n6236), .C(n6237) );
  BUFFD0 U6120 ( .I(n6237), .Z(n6238) );
  CKBD0 U6121 ( .CLK(n6238), .C(n6239) );
  CKBD0 U6122 ( .CLK(n6239), .C(n6240) );
  CKBD0 U6123 ( .CLK(n6240), .C(n6241) );
  CKBD0 U6124 ( .CLK(n6241), .C(n6242) );
  CKBD0 U6125 ( .CLK(n6242), .C(n6243) );
  CKBD0 U6126 ( .CLK(n6243), .C(n6244) );
  CKBD0 U6127 ( .CLK(n6244), .C(n6245) );
  CKBD0 U6128 ( .CLK(n6245), .C(n6246) );
  CKBD0 U6129 ( .CLK(n6246), .C(n6247) );
  CKBD0 U6130 ( .CLK(n6247), .C(n6248) );
  BUFFD0 U6131 ( .I(n6248), .Z(n6249) );
  CKBD0 U6132 ( .CLK(n6249), .C(n6250) );
  CKBD0 U6133 ( .CLK(n6250), .C(n6251) );
  CKBD0 U6134 ( .CLK(n6251), .C(n6252) );
  CKBD0 U6135 ( .CLK(n6252), .C(n6253) );
  CKBD0 U6136 ( .CLK(n6253), .C(n6254) );
  CKBD0 U6137 ( .CLK(n6254), .C(n6255) );
  CKBD0 U6138 ( .CLK(n6255), .C(n6256) );
  CKBD0 U6139 ( .CLK(n6256), .C(n6257) );
  CKBD0 U6140 ( .CLK(n6257), .C(n6258) );
  CKBD0 U6141 ( .CLK(n6258), .C(n6259) );
  BUFFD0 U6142 ( .I(n6259), .Z(n6260) );
  CKBD0 U6143 ( .CLK(n6260), .C(n6261) );
  CKBD0 U6144 ( .CLK(n6261), .C(n6262) );
  CKBD0 U6145 ( .CLK(n6262), .C(n6263) );
  CKBD0 U6146 ( .CLK(n6263), .C(n6264) );
  CKBD0 U6147 ( .CLK(n6264), .C(n6265) );
  BUFFD0 U6148 ( .I(n6265), .Z(n6266) );
  CKBD0 U6149 ( .CLK(n6266), .C(n6267) );
  BUFFD0 U6150 ( .I(n6267), .Z(n6268) );
  CKBD0 U6151 ( .CLK(n6268), .C(n6269) );
  BUFFD0 U6152 ( .I(n6269), .Z(n6270) );
  CKBD0 U6153 ( .CLK(n6270), .C(n6271) );
  BUFFD0 U6154 ( .I(n6271), .Z(n6272) );
  CKBD0 U6155 ( .CLK(n6272), .C(n6273) );
  BUFFD0 U6156 ( .I(n6273), .Z(n6274) );
  CKBD0 U6157 ( .CLK(n6274), .C(n6275) );
  BUFFD0 U6158 ( .I(n6275), .Z(n6276) );
  CKBD0 U6159 ( .CLK(n6276), .C(n6277) );
  BUFFD0 U6160 ( .I(n6277), .Z(n6278) );
  CKBD0 U6161 ( .CLK(n6278), .C(n6279) );
  BUFFD0 U6162 ( .I(n6279), .Z(n6280) );
  BUFFD0 U6163 ( .I(n9195), .Z(n6281) );
  BUFFD0 U6164 ( .I(n6283), .Z(n6282) );
  BUFFD0 U6165 ( .I(n6284), .Z(n6283) );
  BUFFD0 U6166 ( .I(Decoder[4]), .Z(n6284) );
  CKBD0 U6167 ( .CLK(n946), .C(n6285) );
  CKBD0 U6168 ( .CLK(n6285), .C(n6286) );
  CKBD0 U6169 ( .CLK(n6286), .C(n6287) );
  CKBD0 U6170 ( .CLK(n6287), .C(n6288) );
  BUFFD0 U6171 ( .I(n6288), .Z(n6289) );
  CKBD0 U6172 ( .CLK(n6289), .C(n6290) );
  CKBD0 U6173 ( .CLK(n6290), .C(n6291) );
  CKBD0 U6174 ( .CLK(n6291), .C(n6292) );
  CKBD0 U6175 ( .CLK(n6292), .C(n6293) );
  CKBD0 U6176 ( .CLK(n6293), .C(n6294) );
  CKBD0 U6177 ( .CLK(n6294), .C(n6295) );
  CKBD0 U6178 ( .CLK(n6295), .C(n6296) );
  CKBD0 U6179 ( .CLK(n6296), .C(n6297) );
  CKBD0 U6180 ( .CLK(n6297), .C(n6298) );
  BUFFD0 U6181 ( .I(n6298), .Z(n6299) );
  CKBD0 U6182 ( .CLK(n6299), .C(n6300) );
  CKBD0 U6183 ( .CLK(n6300), .C(n6301) );
  CKBD0 U6184 ( .CLK(n6301), .C(n6302) );
  CKBD0 U6185 ( .CLK(n6302), .C(n6303) );
  CKBD0 U6186 ( .CLK(n6303), .C(n6304) );
  CKBD0 U6187 ( .CLK(n6304), .C(n6305) );
  CKBD0 U6188 ( .CLK(n6305), .C(n6306) );
  CKBD0 U6189 ( .CLK(n6306), .C(n6307) );
  CKBD0 U6190 ( .CLK(n6307), .C(n6308) );
  CKBD0 U6191 ( .CLK(n6308), .C(n6309) );
  BUFFD0 U6192 ( .I(n6309), .Z(n6310) );
  CKBD0 U6193 ( .CLK(n6310), .C(n6311) );
  CKBD0 U6194 ( .CLK(n6311), .C(n6312) );
  CKBD0 U6195 ( .CLK(n6312), .C(n6313) );
  CKBD0 U6196 ( .CLK(n6313), .C(n6314) );
  CKBD0 U6197 ( .CLK(n6314), .C(n6315) );
  CKBD0 U6198 ( .CLK(n6315), .C(n6316) );
  CKBD0 U6199 ( .CLK(n6316), .C(n6317) );
  CKBD0 U6200 ( .CLK(n6317), .C(n6318) );
  CKBD0 U6201 ( .CLK(n6318), .C(n6319) );
  CKBD0 U6202 ( .CLK(n6319), .C(n6320) );
  BUFFD0 U6203 ( .I(n6320), .Z(n6321) );
  CKBD0 U6204 ( .CLK(n6321), .C(n6322) );
  CKBD0 U6205 ( .CLK(n6322), .C(n6323) );
  CKBD0 U6206 ( .CLK(n6323), .C(n6324) );
  CKBD0 U6207 ( .CLK(n6324), .C(n6325) );
  CKBD0 U6208 ( .CLK(n6325), .C(n6326) );
  CKBD0 U6209 ( .CLK(n6326), .C(n6327) );
  CKBD0 U6210 ( .CLK(n6327), .C(n6328) );
  CKBD0 U6211 ( .CLK(n6328), .C(n6329) );
  CKBD0 U6212 ( .CLK(n6329), .C(n6330) );
  CKBD0 U6213 ( .CLK(n6330), .C(n6331) );
  BUFFD0 U6214 ( .I(n6331), .Z(n6332) );
  CKBD0 U6215 ( .CLK(n6332), .C(n6333) );
  CKBD0 U6216 ( .CLK(n6333), .C(n6334) );
  CKBD0 U6217 ( .CLK(n6334), .C(n6335) );
  CKBD0 U6218 ( .CLK(n6335), .C(n6336) );
  CKBD0 U6219 ( .CLK(n6336), .C(n6337) );
  CKBD0 U6220 ( .CLK(n6337), .C(n6338) );
  CKBD0 U6221 ( .CLK(n6338), .C(n6339) );
  CKBD0 U6222 ( .CLK(n6339), .C(n6340) );
  CKBD0 U6223 ( .CLK(n6340), .C(n6341) );
  BUFFD0 U6224 ( .I(n6341), .Z(n6342) );
  CKBD0 U6225 ( .CLK(n6342), .C(n6343) );
  CKBD0 U6226 ( .CLK(n6343), .C(n6344) );
  CKBD0 U6227 ( .CLK(n6344), .C(n6345) );
  CKBD0 U6228 ( .CLK(n6345), .C(n6346) );
  CKBD0 U6229 ( .CLK(n6346), .C(n6347) );
  CKBD0 U6230 ( .CLK(n6347), .C(n6348) );
  CKBD0 U6231 ( .CLK(n6348), .C(n6349) );
  CKBD0 U6232 ( .CLK(n6349), .C(n6350) );
  CKBD0 U6233 ( .CLK(n6350), .C(n6351) );
  CKBD0 U6234 ( .CLK(n6351), .C(n6352) );
  CKBD0 U6235 ( .CLK(n6352), .C(n6353) );
  BUFFD0 U6236 ( .I(n6353), .Z(n6354) );
  CKBD0 U6237 ( .CLK(n6354), .C(n6355) );
  CKBD0 U6238 ( .CLK(n6355), .C(n6356) );
  CKBD0 U6239 ( .CLK(n6356), .C(n6357) );
  CKBD0 U6240 ( .CLK(n6357), .C(n6358) );
  CKBD0 U6241 ( .CLK(n6358), .C(n6359) );
  CKBD0 U6242 ( .CLK(n6359), .C(n6360) );
  CKBD0 U6243 ( .CLK(n6360), .C(n6361) );
  CKBD0 U6244 ( .CLK(n6361), .C(n6362) );
  CKBD0 U6245 ( .CLK(n6362), .C(n6363) );
  BUFFD0 U6246 ( .I(n6363), .Z(n6364) );
  CKBD0 U6247 ( .CLK(n6364), .C(n6365) );
  CKBD0 U6248 ( .CLK(n6365), .C(n6366) );
  CKBD0 U6249 ( .CLK(n6366), .C(n6367) );
  CKBD0 U6250 ( .CLK(n6367), .C(n6368) );
  CKBD0 U6251 ( .CLK(n6368), .C(n6369) );
  CKBD0 U6252 ( .CLK(n6369), .C(n6370) );
  CKBD0 U6253 ( .CLK(n6370), .C(n6371) );
  CKBD0 U6254 ( .CLK(n6371), .C(n6372) );
  CKBD0 U6255 ( .CLK(n6372), .C(n6373) );
  BUFFD0 U6256 ( .I(n6373), .Z(n6374) );
  CKBD0 U6257 ( .CLK(n6374), .C(n6375) );
  CKBD0 U6258 ( .CLK(n6375), .C(n6376) );
  CKBD0 U6259 ( .CLK(n6376), .C(n6377) );
  CKBD0 U6260 ( .CLK(n6377), .C(n6378) );
  CKBD0 U6261 ( .CLK(n6378), .C(n6379) );
  CKBD0 U6262 ( .CLK(n6379), .C(n6380) );
  CKBD0 U6263 ( .CLK(n6380), .C(n6381) );
  CKBD0 U6264 ( .CLK(n6381), .C(n6382) );
  CKBD0 U6265 ( .CLK(n6382), .C(n6383) );
  CKBD0 U6266 ( .CLK(n6383), .C(n6384) );
  CKBD0 U6267 ( .CLK(n6384), .C(n6385) );
  BUFFD0 U6268 ( .I(n6385), .Z(n6386) );
  CKBD0 U6269 ( .CLK(n6386), .C(n6387) );
  CKBD0 U6270 ( .CLK(n6387), .C(n6388) );
  CKBD0 U6271 ( .CLK(n6388), .C(n6389) );
  CKBD0 U6272 ( .CLK(n6389), .C(n6390) );
  CKBD0 U6273 ( .CLK(n6390), .C(n6391) );
  CKBD0 U6274 ( .CLK(n6391), .C(n6392) );
  CKBD0 U6275 ( .CLK(n6392), .C(n6393) );
  CKBD0 U6276 ( .CLK(n6393), .C(n6394) );
  CKBD0 U6277 ( .CLK(n6394), .C(n6395) );
  CKBD0 U6278 ( .CLK(n6395), .C(n6396) );
  BUFFD0 U6279 ( .I(n6396), .Z(n6397) );
  CKBD0 U6280 ( .CLK(n6397), .C(n6398) );
  CKBD0 U6281 ( .CLK(n6398), .C(n6399) );
  CKBD0 U6282 ( .CLK(n6399), .C(n6400) );
  CKBD0 U6283 ( .CLK(n6400), .C(n6401) );
  CKBD0 U6284 ( .CLK(n6401), .C(n6402) );
  BUFFD0 U6285 ( .I(n6402), .Z(n6403) );
  CKBD0 U6286 ( .CLK(n6403), .C(n6404) );
  BUFFD0 U6287 ( .I(n6404), .Z(n6405) );
  CKBD0 U6288 ( .CLK(n6405), .C(n6406) );
  BUFFD0 U6289 ( .I(n6406), .Z(n6407) );
  CKBD0 U6290 ( .CLK(n6407), .C(n6408) );
  BUFFD0 U6291 ( .I(n6408), .Z(n6409) );
  CKBD0 U6292 ( .CLK(n6409), .C(n6410) );
  BUFFD0 U6293 ( .I(n6410), .Z(n6411) );
  CKBD0 U6294 ( .CLK(n6411), .C(n6412) );
  BUFFD0 U6295 ( .I(n6412), .Z(n6413) );
  CKBD0 U6296 ( .CLK(n6413), .C(n6414) );
  BUFFD0 U6297 ( .I(n6414), .Z(n6415) );
  CKBD0 U6298 ( .CLK(n6415), .C(n6416) );
  BUFFD0 U6299 ( .I(n6416), .Z(n6417) );
  BUFFD0 U6300 ( .I(n9196), .Z(n6418) );
  BUFFD0 U6301 ( .I(n6420), .Z(n6419) );
  BUFFD0 U6302 ( .I(n6421), .Z(n6420) );
  BUFFD0 U6303 ( .I(Decoder[3]), .Z(n6421) );
  CKBD0 U6304 ( .CLK(n944), .C(n6422) );
  CKBD0 U6305 ( .CLK(n6422), .C(n6423) );
  CKBD0 U6306 ( .CLK(n6423), .C(n6424) );
  BUFFD0 U6307 ( .I(n6424), .Z(n6425) );
  CKBD0 U6308 ( .CLK(n6425), .C(n6426) );
  CKBD0 U6309 ( .CLK(n6426), .C(n6427) );
  CKBD0 U6310 ( .CLK(n6427), .C(n6428) );
  CKBD0 U6311 ( .CLK(n6428), .C(n6429) );
  CKBD0 U6312 ( .CLK(n6429), .C(n6430) );
  CKBD0 U6313 ( .CLK(n6430), .C(n6431) );
  CKBD0 U6314 ( .CLK(n6431), .C(n6432) );
  CKBD0 U6315 ( .CLK(n6432), .C(n6433) );
  CKBD0 U6316 ( .CLK(n6433), .C(n6434) );
  CKBD0 U6317 ( .CLK(n6434), .C(n6435) );
  BUFFD0 U6318 ( .I(n6435), .Z(n6436) );
  CKBD0 U6319 ( .CLK(n6436), .C(n6437) );
  CKBD0 U6320 ( .CLK(n6437), .C(n6438) );
  CKBD0 U6321 ( .CLK(n6438), .C(n6439) );
  CKBD0 U6322 ( .CLK(n6439), .C(n6440) );
  CKBD0 U6323 ( .CLK(n6440), .C(n6441) );
  CKBD0 U6324 ( .CLK(n6441), .C(n6442) );
  CKBD0 U6325 ( .CLK(n6442), .C(n6443) );
  CKBD0 U6326 ( .CLK(n6443), .C(n6444) );
  CKBD0 U6327 ( .CLK(n6444), .C(n6445) );
  CKBD0 U6328 ( .CLK(n6445), .C(n6446) );
  BUFFD0 U6329 ( .I(n6446), .Z(n6447) );
  CKBD0 U6330 ( .CLK(n6447), .C(n6448) );
  CKBD0 U6331 ( .CLK(n6448), .C(n6449) );
  CKBD0 U6332 ( .CLK(n6449), .C(n6450) );
  CKBD0 U6333 ( .CLK(n6450), .C(n6451) );
  CKBD0 U6334 ( .CLK(n6451), .C(n6452) );
  CKBD0 U6335 ( .CLK(n6452), .C(n6453) );
  CKBD0 U6336 ( .CLK(n6453), .C(n6454) );
  CKBD0 U6337 ( .CLK(n6454), .C(n6455) );
  CKBD0 U6338 ( .CLK(n6455), .C(n6456) );
  BUFFD0 U6339 ( .I(n6456), .Z(n6457) );
  CKBD0 U6340 ( .CLK(n6457), .C(n6458) );
  CKBD0 U6341 ( .CLK(n6458), .C(n6459) );
  CKBD0 U6342 ( .CLK(n6459), .C(n6460) );
  CKBD0 U6343 ( .CLK(n6460), .C(n6461) );
  CKBD0 U6344 ( .CLK(n6461), .C(n6462) );
  CKBD0 U6345 ( .CLK(n6462), .C(n6463) );
  CKBD0 U6346 ( .CLK(n6463), .C(n6464) );
  CKBD0 U6347 ( .CLK(n6464), .C(n6465) );
  CKBD0 U6348 ( .CLK(n6465), .C(n6466) );
  CKBD0 U6349 ( .CLK(n6466), .C(n6467) );
  CKBD0 U6350 ( .CLK(n6467), .C(n6468) );
  BUFFD0 U6351 ( .I(n6468), .Z(n6469) );
  CKBD0 U6352 ( .CLK(n6469), .C(n6470) );
  CKBD0 U6353 ( .CLK(n6470), .C(n6471) );
  CKBD0 U6354 ( .CLK(n6471), .C(n6472) );
  CKBD0 U6355 ( .CLK(n6472), .C(n6473) );
  CKBD0 U6356 ( .CLK(n6473), .C(n6474) );
  CKBD0 U6357 ( .CLK(n6474), .C(n6475) );
  CKBD0 U6358 ( .CLK(n6475), .C(n6476) );
  CKBD0 U6359 ( .CLK(n6476), .C(n6477) );
  CKBD0 U6360 ( .CLK(n6477), .C(n6478) );
  CKBD0 U6361 ( .CLK(n6478), .C(n6479) );
  BUFFD0 U6362 ( .I(n6479), .Z(n6480) );
  CKBD0 U6363 ( .CLK(n6480), .C(n6481) );
  CKBD0 U6364 ( .CLK(n6481), .C(n6482) );
  CKBD0 U6365 ( .CLK(n6482), .C(n6483) );
  CKBD0 U6366 ( .CLK(n6483), .C(n6484) );
  CKBD0 U6367 ( .CLK(n6484), .C(n6485) );
  CKBD0 U6368 ( .CLK(n6485), .C(n6486) );
  CKBD0 U6369 ( .CLK(n6486), .C(n6487) );
  CKBD0 U6370 ( .CLK(n6487), .C(n6488) );
  CKBD0 U6371 ( .CLK(n6488), .C(n6489) );
  BUFFD0 U6372 ( .I(n6489), .Z(n6490) );
  CKBD0 U6373 ( .CLK(n6490), .C(n6491) );
  CKBD0 U6374 ( .CLK(n6491), .C(n6492) );
  CKBD0 U6375 ( .CLK(n6492), .C(n6493) );
  CKBD0 U6376 ( .CLK(n6493), .C(n6494) );
  CKBD0 U6377 ( .CLK(n6494), .C(n6495) );
  CKBD0 U6378 ( .CLK(n6495), .C(n6496) );
  CKBD0 U6379 ( .CLK(n6496), .C(n6497) );
  CKBD0 U6380 ( .CLK(n6497), .C(n6498) );
  CKBD0 U6381 ( .CLK(n6498), .C(n6499) );
  CKBD0 U6382 ( .CLK(n6499), .C(n6500) );
  CKBD0 U6383 ( .CLK(n6500), .C(n6501) );
  BUFFD0 U6384 ( .I(n6501), .Z(n6502) );
  CKBD0 U6385 ( .CLK(n6502), .C(n6503) );
  CKBD0 U6386 ( .CLK(n6503), .C(n6504) );
  CKBD0 U6387 ( .CLK(n6504), .C(n6505) );
  CKBD0 U6388 ( .CLK(n6505), .C(n6506) );
  CKBD0 U6389 ( .CLK(n6506), .C(n6507) );
  CKBD0 U6390 ( .CLK(n6507), .C(n6508) );
  CKBD0 U6391 ( .CLK(n6508), .C(n6509) );
  CKBD0 U6392 ( .CLK(n6509), .C(n6510) );
  CKBD0 U6393 ( .CLK(n6510), .C(n6511) );
  BUFFD0 U6394 ( .I(n6511), .Z(n6512) );
  CKBD0 U6395 ( .CLK(n6512), .C(n6513) );
  CKBD0 U6396 ( .CLK(n6513), .C(n6514) );
  CKBD0 U6397 ( .CLK(n6514), .C(n6515) );
  CKBD0 U6398 ( .CLK(n6515), .C(n6516) );
  CKBD0 U6399 ( .CLK(n6516), .C(n6517) );
  CKBD0 U6400 ( .CLK(n6517), .C(n6518) );
  CKBD0 U6401 ( .CLK(n6518), .C(n6519) );
  CKBD0 U6402 ( .CLK(n6519), .C(n6520) );
  CKBD0 U6403 ( .CLK(n6520), .C(n6521) );
  BUFFD0 U6404 ( .I(n6521), .Z(n6522) );
  CKBD0 U6405 ( .CLK(n6522), .C(n6523) );
  CKBD0 U6406 ( .CLK(n6523), .C(n6524) );
  CKBD0 U6407 ( .CLK(n6524), .C(n6525) );
  CKBD0 U6408 ( .CLK(n6525), .C(n6526) );
  CKBD0 U6409 ( .CLK(n6526), .C(n6527) );
  CKBD0 U6410 ( .CLK(n6527), .C(n6528) );
  CKBD0 U6411 ( .CLK(n6528), .C(n6529) );
  CKBD0 U6412 ( .CLK(n6529), .C(n6530) );
  CKBD0 U6413 ( .CLK(n6530), .C(n6531) );
  CKBD0 U6414 ( .CLK(n6531), .C(n6532) );
  CKBD0 U6415 ( .CLK(n6532), .C(n6533) );
  BUFFD0 U6416 ( .I(n6533), .Z(n6534) );
  CKBD0 U6417 ( .CLK(n6534), .C(n6535) );
  CKBD0 U6418 ( .CLK(n6535), .C(n6536) );
  CKBD0 U6419 ( .CLK(n6536), .C(n6537) );
  CKBD0 U6420 ( .CLK(n6537), .C(n6538) );
  CKBD0 U6421 ( .CLK(n6538), .C(n6539) );
  BUFFD0 U6422 ( .I(n6539), .Z(n6540) );
  CKBD0 U6423 ( .CLK(n6540), .C(n6541) );
  BUFFD0 U6424 ( .I(n6541), .Z(n6542) );
  CKBD0 U6425 ( .CLK(n6542), .C(n6543) );
  BUFFD0 U6426 ( .I(n6543), .Z(n6544) );
  CKBD0 U6427 ( .CLK(n6544), .C(n6545) );
  BUFFD0 U6428 ( .I(n6545), .Z(n6546) );
  CKBD0 U6429 ( .CLK(n6546), .C(n6547) );
  BUFFD0 U6430 ( .I(n6547), .Z(n6548) );
  CKBD0 U6431 ( .CLK(n6548), .C(n6549) );
  BUFFD0 U6432 ( .I(n6549), .Z(n6550) );
  CKBD0 U6433 ( .CLK(n6550), .C(n6551) );
  BUFFD0 U6434 ( .I(n6551), .Z(n6552) );
  CKBD0 U6435 ( .CLK(n6552), .C(n6553) );
  BUFFD0 U6436 ( .I(n6553), .Z(n6554) );
  BUFFD0 U6437 ( .I(n9197), .Z(n6555) );
  BUFFD0 U6438 ( .I(n6557), .Z(n6556) );
  BUFFD0 U6439 ( .I(n6558), .Z(n6557) );
  BUFFD0 U6440 ( .I(Decoder[2]), .Z(n6558) );
  CKBD0 U6441 ( .CLK(n942), .C(n6559) );
  CKBD0 U6442 ( .CLK(n6559), .C(n6560) );
  CKBD0 U6443 ( .CLK(n6560), .C(n6561) );
  CKBD0 U6444 ( .CLK(n6561), .C(n6562) );
  BUFFD0 U6445 ( .I(n6562), .Z(n6563) );
  CKBD0 U6446 ( .CLK(n6563), .C(n6564) );
  CKBD0 U6447 ( .CLK(n6564), .C(n6565) );
  CKBD0 U6448 ( .CLK(n6565), .C(n6566) );
  CKBD0 U6449 ( .CLK(n6566), .C(n6567) );
  CKBD0 U6450 ( .CLK(n6567), .C(n6568) );
  CKBD0 U6451 ( .CLK(n6568), .C(n6569) );
  CKBD0 U6452 ( .CLK(n6569), .C(n6570) );
  CKBD0 U6453 ( .CLK(n6570), .C(n6571) );
  CKBD0 U6454 ( .CLK(n6571), .C(n6572) );
  BUFFD0 U6455 ( .I(n6572), .Z(n6573) );
  CKBD0 U6456 ( .CLK(n6573), .C(n6574) );
  CKBD0 U6457 ( .CLK(n6574), .C(n6575) );
  CKBD0 U6458 ( .CLK(n6575), .C(n6576) );
  CKBD0 U6459 ( .CLK(n6576), .C(n6577) );
  CKBD0 U6460 ( .CLK(n6577), .C(n6578) );
  CKBD0 U6461 ( .CLK(n6578), .C(n6579) );
  CKBD0 U6462 ( .CLK(n6579), .C(n6580) );
  CKBD0 U6463 ( .CLK(n6580), .C(n6581) );
  CKBD0 U6464 ( .CLK(n6581), .C(n6582) );
  CKBD0 U6465 ( .CLK(n6582), .C(n6583) );
  BUFFD0 U6466 ( .I(n6583), .Z(n6584) );
  CKBD0 U6467 ( .CLK(n6584), .C(n6585) );
  CKBD0 U6468 ( .CLK(n6585), .C(n6586) );
  CKBD0 U6469 ( .CLK(n6586), .C(n6587) );
  CKBD0 U6470 ( .CLK(n6587), .C(n6588) );
  CKBD0 U6471 ( .CLK(n6588), .C(n6589) );
  CKBD0 U6472 ( .CLK(n6589), .C(n6590) );
  CKBD0 U6473 ( .CLK(n6590), .C(n6591) );
  CKBD0 U6474 ( .CLK(n6591), .C(n6592) );
  CKBD0 U6475 ( .CLK(n6592), .C(n6593) );
  CKBD0 U6476 ( .CLK(n6593), .C(n6594) );
  BUFFD0 U6477 ( .I(n6594), .Z(n6595) );
  CKBD0 U6478 ( .CLK(n6595), .C(n6596) );
  CKBD0 U6479 ( .CLK(n6596), .C(n6597) );
  CKBD0 U6480 ( .CLK(n6597), .C(n6598) );
  CKBD0 U6481 ( .CLK(n6598), .C(n6599) );
  CKBD0 U6482 ( .CLK(n6599), .C(n6600) );
  CKBD0 U6483 ( .CLK(n6600), .C(n6601) );
  CKBD0 U6484 ( .CLK(n6601), .C(n6602) );
  CKBD0 U6485 ( .CLK(n6602), .C(n6603) );
  CKBD0 U6486 ( .CLK(n6603), .C(n6604) );
  BUFFD0 U6487 ( .I(n6604), .Z(n6605) );
  CKBD0 U6488 ( .CLK(n6605), .C(n6606) );
  CKBD0 U6489 ( .CLK(n6606), .C(n6607) );
  CKBD0 U6490 ( .CLK(n6607), .C(n6608) );
  CKBD0 U6491 ( .CLK(n6608), .C(n6609) );
  CKBD0 U6492 ( .CLK(n6609), .C(n6610) );
  CKBD0 U6493 ( .CLK(n6610), .C(n6611) );
  CKBD0 U6494 ( .CLK(n6611), .C(n6612) );
  CKBD0 U6495 ( .CLK(n6612), .C(n6613) );
  CKBD0 U6496 ( .CLK(n6613), .C(n6614) );
  CKBD0 U6497 ( .CLK(n6614), .C(n6615) );
  CKBD0 U6498 ( .CLK(n6615), .C(n6616) );
  BUFFD0 U6499 ( .I(n6616), .Z(n6617) );
  CKBD0 U6500 ( .CLK(n6617), .C(n6618) );
  CKBD0 U6501 ( .CLK(n6618), .C(n6619) );
  CKBD0 U6502 ( .CLK(n6619), .C(n6620) );
  CKBD0 U6503 ( .CLK(n6620), .C(n6621) );
  CKBD0 U6504 ( .CLK(n6621), .C(n6622) );
  CKBD0 U6505 ( .CLK(n6622), .C(n6623) );
  CKBD0 U6506 ( .CLK(n6623), .C(n6624) );
  CKBD0 U6507 ( .CLK(n6624), .C(n6625) );
  CKBD0 U6508 ( .CLK(n6625), .C(n6626) );
  BUFFD0 U6509 ( .I(n6626), .Z(n6627) );
  CKBD0 U6510 ( .CLK(n6627), .C(n6628) );
  CKBD0 U6511 ( .CLK(n6628), .C(n6629) );
  CKBD0 U6512 ( .CLK(n6629), .C(n6630) );
  CKBD0 U6513 ( .CLK(n6630), .C(n6631) );
  CKBD0 U6514 ( .CLK(n6631), .C(n6632) );
  CKBD0 U6515 ( .CLK(n6632), .C(n6633) );
  CKBD0 U6516 ( .CLK(n6633), .C(n6634) );
  CKBD0 U6517 ( .CLK(n6634), .C(n6635) );
  CKBD0 U6518 ( .CLK(n6635), .C(n6636) );
  CKBD0 U6519 ( .CLK(n6636), .C(n6637) );
  BUFFD0 U6520 ( .I(n6637), .Z(n6638) );
  CKBD0 U6521 ( .CLK(n6638), .C(n6639) );
  CKBD0 U6522 ( .CLK(n6639), .C(n6640) );
  CKBD0 U6523 ( .CLK(n6640), .C(n6641) );
  CKBD0 U6524 ( .CLK(n6641), .C(n6642) );
  CKBD0 U6525 ( .CLK(n6642), .C(n6643) );
  CKBD0 U6526 ( .CLK(n6643), .C(n6644) );
  CKBD0 U6527 ( .CLK(n6644), .C(n6645) );
  CKBD0 U6528 ( .CLK(n6645), .C(n6646) );
  CKBD0 U6529 ( .CLK(n6646), .C(n6647) );
  CKBD0 U6530 ( .CLK(n6647), .C(n6648) );
  CKBD0 U6531 ( .CLK(n6648), .C(n6649) );
  BUFFD0 U6532 ( .I(n6649), .Z(n6650) );
  CKBD0 U6533 ( .CLK(n6650), .C(n6651) );
  CKBD0 U6534 ( .CLK(n6651), .C(n6652) );
  CKBD0 U6535 ( .CLK(n6652), .C(n6653) );
  CKBD0 U6536 ( .CLK(n6653), .C(n6654) );
  CKBD0 U6537 ( .CLK(n6654), .C(n6655) );
  CKBD0 U6538 ( .CLK(n6655), .C(n6656) );
  CKBD0 U6539 ( .CLK(n6656), .C(n6657) );
  CKBD0 U6540 ( .CLK(n6657), .C(n6658) );
  CKBD0 U6541 ( .CLK(n6658), .C(n6659) );
  BUFFD0 U6542 ( .I(n6659), .Z(n6660) );
  CKBD0 U6543 ( .CLK(n6660), .C(n6661) );
  CKBD0 U6544 ( .CLK(n6661), .C(n6662) );
  CKBD0 U6545 ( .CLK(n6662), .C(n6663) );
  CKBD0 U6546 ( .CLK(n6663), .C(n6664) );
  CKBD0 U6547 ( .CLK(n6664), .C(n6665) );
  CKBD0 U6548 ( .CLK(n6665), .C(n6666) );
  CKBD0 U6549 ( .CLK(n6666), .C(n6667) );
  CKBD0 U6550 ( .CLK(n6667), .C(n6668) );
  CKBD0 U6551 ( .CLK(n6668), .C(n6669) );
  BUFFD0 U6552 ( .I(n6669), .Z(n6670) );
  CKBD0 U6553 ( .CLK(n6670), .C(n6671) );
  CKBD0 U6554 ( .CLK(n6671), .C(n6672) );
  CKBD0 U6555 ( .CLK(n6672), .C(n6673) );
  CKBD0 U6556 ( .CLK(n6673), .C(n6674) );
  CKBD0 U6557 ( .CLK(n6674), .C(n6675) );
  CKBD0 U6558 ( .CLK(n6675), .C(n6676) );
  BUFFD0 U6559 ( .I(n6676), .Z(n6677) );
  CKBD0 U6560 ( .CLK(n6677), .C(n6678) );
  BUFFD0 U6561 ( .I(n6678), .Z(n6679) );
  CKBD0 U6562 ( .CLK(n6679), .C(n6680) );
  BUFFD0 U6563 ( .I(n6680), .Z(n6681) );
  CKBD0 U6564 ( .CLK(n6681), .C(n6682) );
  BUFFD0 U6565 ( .I(n6682), .Z(n6683) );
  CKBD0 U6566 ( .CLK(n6683), .C(n6684) );
  BUFFD0 U6567 ( .I(n6684), .Z(n6685) );
  CKBD0 U6568 ( .CLK(n6685), .C(n6686) );
  BUFFD0 U6569 ( .I(n6686), .Z(n6687) );
  CKBD0 U6570 ( .CLK(n6687), .C(n6688) );
  BUFFD0 U6571 ( .I(n6688), .Z(n6689) );
  CKBD0 U6572 ( .CLK(n6689), .C(n6690) );
  BUFFD0 U6573 ( .I(n6690), .Z(n6691) );
  BUFFD0 U6574 ( .I(n9198), .Z(n6692) );
  BUFFD0 U6575 ( .I(n6694), .Z(n6693) );
  BUFFD0 U6576 ( .I(n6695), .Z(n6694) );
  BUFFD0 U6577 ( .I(Decoder[1]), .Z(n6695) );
  CKBD0 U6578 ( .CLK(n940), .C(n6696) );
  CKBD0 U6579 ( .CLK(n6696), .C(n6697) );
  CKBD0 U6580 ( .CLK(n6697), .C(n6698) );
  BUFFD0 U6581 ( .I(n6698), .Z(n6699) );
  CKBD0 U6582 ( .CLK(n6699), .C(n6700) );
  CKBD0 U6583 ( .CLK(n6700), .C(n6701) );
  CKBD0 U6584 ( .CLK(n6701), .C(n6702) );
  CKBD0 U6585 ( .CLK(n6702), .C(n6703) );
  CKBD0 U6586 ( .CLK(n6703), .C(n6704) );
  CKBD0 U6587 ( .CLK(n6704), .C(n6705) );
  CKBD0 U6588 ( .CLK(n6705), .C(n6706) );
  CKBD0 U6589 ( .CLK(n6706), .C(n6707) );
  CKBD0 U6590 ( .CLK(n6707), .C(n6708) );
  CKBD0 U6591 ( .CLK(n6708), .C(n6709) );
  BUFFD0 U6592 ( .I(n6709), .Z(n6710) );
  CKBD0 U6593 ( .CLK(n6710), .C(n6711) );
  CKBD0 U6594 ( .CLK(n6711), .C(n6712) );
  CKBD0 U6595 ( .CLK(n6712), .C(n6713) );
  CKBD0 U6596 ( .CLK(n6713), .C(n6714) );
  CKBD0 U6597 ( .CLK(n6714), .C(n6715) );
  CKBD0 U6598 ( .CLK(n6715), .C(n6716) );
  CKBD0 U6599 ( .CLK(n6716), .C(n6717) );
  CKBD0 U6600 ( .CLK(n6717), .C(n6718) );
  CKBD0 U6601 ( .CLK(n6718), .C(n6719) );
  CKBD0 U6602 ( .CLK(n6719), .C(n6720) );
  BUFFD0 U6603 ( .I(n6720), .Z(n6721) );
  CKBD0 U6604 ( .CLK(n6721), .C(n6722) );
  CKBD0 U6605 ( .CLK(n6722), .C(n6723) );
  CKBD0 U6606 ( .CLK(n6723), .C(n6724) );
  CKBD0 U6607 ( .CLK(n6724), .C(n6725) );
  CKBD0 U6608 ( .CLK(n6725), .C(n6726) );
  CKBD0 U6609 ( .CLK(n6726), .C(n6727) );
  CKBD0 U6610 ( .CLK(n6727), .C(n6728) );
  CKBD0 U6611 ( .CLK(n6728), .C(n6729) );
  CKBD0 U6612 ( .CLK(n6729), .C(n6730) );
  BUFFD0 U6613 ( .I(n6730), .Z(n6731) );
  CKBD0 U6614 ( .CLK(n6731), .C(n6732) );
  CKBD0 U6615 ( .CLK(n6732), .C(n6733) );
  CKBD0 U6616 ( .CLK(n6733), .C(n6734) );
  CKBD0 U6617 ( .CLK(n6734), .C(n6735) );
  CKBD0 U6618 ( .CLK(n6735), .C(n6736) );
  CKBD0 U6619 ( .CLK(n6736), .C(n6737) );
  CKBD0 U6620 ( .CLK(n6737), .C(n6738) );
  CKBD0 U6621 ( .CLK(n6738), .C(n6739) );
  CKBD0 U6622 ( .CLK(n6739), .C(n6740) );
  CKBD0 U6623 ( .CLK(n6740), .C(n6741) );
  CKBD0 U6624 ( .CLK(n6741), .C(n6742) );
  BUFFD0 U6625 ( .I(n6742), .Z(n6743) );
  CKBD0 U6626 ( .CLK(n6743), .C(n6744) );
  CKBD0 U6627 ( .CLK(n6744), .C(n6745) );
  CKBD0 U6628 ( .CLK(n6745), .C(n6746) );
  CKBD0 U6629 ( .CLK(n6746), .C(n6747) );
  CKBD0 U6630 ( .CLK(n6747), .C(n6748) );
  CKBD0 U6631 ( .CLK(n6748), .C(n6749) );
  CKBD0 U6632 ( .CLK(n6749), .C(n6750) );
  CKBD0 U6633 ( .CLK(n6750), .C(n6751) );
  CKBD0 U6634 ( .CLK(n6751), .C(n6752) );
  BUFFD0 U6635 ( .I(n6752), .Z(n6753) );
  CKBD0 U6636 ( .CLK(n6753), .C(n6754) );
  CKBD0 U6637 ( .CLK(n6754), .C(n6755) );
  CKBD0 U6638 ( .CLK(n6755), .C(n6756) );
  CKBD0 U6639 ( .CLK(n6756), .C(n6757) );
  CKBD0 U6640 ( .CLK(n6757), .C(n6758) );
  CKBD0 U6641 ( .CLK(n6758), .C(n6759) );
  CKBD0 U6642 ( .CLK(n6759), .C(n6760) );
  CKBD0 U6643 ( .CLK(n6760), .C(n6761) );
  CKBD0 U6644 ( .CLK(n6761), .C(n6762) );
  CKBD0 U6645 ( .CLK(n6762), .C(n6763) );
  BUFFD0 U6646 ( .I(n6763), .Z(n6764) );
  CKBD0 U6647 ( .CLK(n6764), .C(n6765) );
  CKBD0 U6648 ( .CLK(n6765), .C(n6766) );
  CKBD0 U6649 ( .CLK(n6766), .C(n6767) );
  CKBD0 U6650 ( .CLK(n6767), .C(n6768) );
  CKBD0 U6651 ( .CLK(n6768), .C(n6769) );
  CKBD0 U6652 ( .CLK(n6769), .C(n6770) );
  CKBD0 U6653 ( .CLK(n6770), .C(n6771) );
  CKBD0 U6654 ( .CLK(n6771), .C(n6772) );
  CKBD0 U6655 ( .CLK(n6772), .C(n6773) );
  CKBD0 U6656 ( .CLK(n6773), .C(n6774) );
  BUFFD0 U6657 ( .I(n6774), .Z(n6775) );
  CKBD0 U6658 ( .CLK(n6775), .C(n6776) );
  CKBD0 U6659 ( .CLK(n6776), .C(n6777) );
  CKBD0 U6660 ( .CLK(n6777), .C(n6778) );
  CKBD0 U6661 ( .CLK(n6778), .C(n6779) );
  CKBD0 U6662 ( .CLK(n6779), .C(n6780) );
  CKBD0 U6663 ( .CLK(n6780), .C(n6781) );
  CKBD0 U6664 ( .CLK(n6781), .C(n6782) );
  CKBD0 U6665 ( .CLK(n6782), .C(n6783) );
  CKBD0 U6666 ( .CLK(n6783), .C(n6784) );
  CKBD0 U6667 ( .CLK(n6784), .C(n6785) );
  BUFFD0 U6668 ( .I(n6785), .Z(n6786) );
  CKBD0 U6669 ( .CLK(n6786), .C(n6787) );
  CKBD0 U6670 ( .CLK(n6787), .C(n6788) );
  CKBD0 U6671 ( .CLK(n6788), .C(n6789) );
  CKBD0 U6672 ( .CLK(n6789), .C(n6790) );
  CKBD0 U6673 ( .CLK(n6790), .C(n6791) );
  CKBD0 U6674 ( .CLK(n6791), .C(n6792) );
  CKBD0 U6675 ( .CLK(n6792), .C(n6793) );
  CKBD0 U6676 ( .CLK(n6793), .C(n6794) );
  CKBD0 U6677 ( .CLK(n6794), .C(n6795) );
  CKBD0 U6678 ( .CLK(n6795), .C(n6796) );
  BUFFD0 U6679 ( .I(n6796), .Z(n6797) );
  CKBD0 U6680 ( .CLK(n6797), .C(n6798) );
  CKBD0 U6681 ( .CLK(n6798), .C(n6799) );
  CKBD0 U6682 ( .CLK(n6799), .C(n6800) );
  CKBD0 U6683 ( .CLK(n6800), .C(n6801) );
  CKBD0 U6684 ( .CLK(n6801), .C(n6802) );
  CKBD0 U6685 ( .CLK(n6802), .C(n6803) );
  CKBD0 U6686 ( .CLK(n6803), .C(n6804) );
  CKBD0 U6687 ( .CLK(n6804), .C(n6805) );
  CKBD0 U6688 ( .CLK(n6805), .C(n6806) );
  CKBD0 U6689 ( .CLK(n6806), .C(n6807) );
  BUFFD0 U6690 ( .I(n6807), .Z(n6808) );
  CKBD0 U6691 ( .CLK(n6808), .C(n6809) );
  CKBD0 U6692 ( .CLK(n6809), .C(n6810) );
  CKBD0 U6693 ( .CLK(n6810), .C(n6811) );
  CKBD0 U6694 ( .CLK(n6811), .C(n6812) );
  CKBD0 U6695 ( .CLK(n6812), .C(n6813) );
  BUFFD0 U6696 ( .I(n6813), .Z(n6814) );
  CKBD0 U6697 ( .CLK(n6814), .C(n6815) );
  BUFFD0 U6698 ( .I(n6815), .Z(n6816) );
  CKBD0 U6699 ( .CLK(n6816), .C(n6817) );
  BUFFD0 U6700 ( .I(n6817), .Z(n6818) );
  CKBD0 U6701 ( .CLK(n6818), .C(n6819) );
  BUFFD0 U6702 ( .I(n6819), .Z(n6820) );
  CKBD0 U6703 ( .CLK(n6820), .C(n6821) );
  BUFFD0 U6704 ( .I(n6821), .Z(n6822) );
  CKBD0 U6705 ( .CLK(n6822), .C(n6823) );
  BUFFD0 U6706 ( .I(n6823), .Z(n6824) );
  CKBD0 U6707 ( .CLK(n6824), .C(n6825) );
  BUFFD0 U6708 ( .I(n6825), .Z(n6826) );
  CKBD0 U6709 ( .CLK(n6826), .C(n6827) );
  BUFFD0 U6710 ( .I(n6827), .Z(n6828) );
  BUFFD0 U6711 ( .I(n9199), .Z(n6829) );
  BUFFD0 U6712 ( .I(n6831), .Z(n6830) );
  BUFFD0 U6713 ( .I(n6832), .Z(n6831) );
  BUFFD0 U6714 ( .I(Decoder[0]), .Z(n6832) );
  CKBD0 U6715 ( .CLK(n938), .C(n6833) );
  CKBD0 U6716 ( .CLK(n6833), .C(n6834) );
  CKBD0 U6717 ( .CLK(n6834), .C(n6835) );
  BUFFD0 U6718 ( .I(n6835), .Z(n6836) );
  CKBD0 U6719 ( .CLK(n6836), .C(n6837) );
  CKBD0 U6720 ( .CLK(n6837), .C(n6838) );
  CKBD0 U6721 ( .CLK(n6838), .C(n6839) );
  CKBD0 U6722 ( .CLK(n6839), .C(n6840) );
  CKBD0 U6723 ( .CLK(n6840), .C(n6841) );
  CKBD0 U6724 ( .CLK(n6841), .C(n6842) );
  CKBD0 U6725 ( .CLK(n6842), .C(n6843) );
  CKBD0 U6726 ( .CLK(n6843), .C(n6844) );
  CKBD0 U6727 ( .CLK(n6844), .C(n6845) );
  CKBD0 U6728 ( .CLK(n6845), .C(n6846) );
  BUFFD0 U6729 ( .I(n6846), .Z(n6847) );
  CKBD0 U6730 ( .CLK(n6847), .C(n6848) );
  CKBD0 U6731 ( .CLK(n6848), .C(n6849) );
  CKBD0 U6732 ( .CLK(n6849), .C(n6850) );
  CKBD0 U6733 ( .CLK(n6850), .C(n6851) );
  CKBD0 U6734 ( .CLK(n6851), .C(n6852) );
  CKBD0 U6735 ( .CLK(n6852), .C(n6853) );
  CKBD0 U6736 ( .CLK(n6853), .C(n6854) );
  CKBD0 U6737 ( .CLK(n6854), .C(n6855) );
  CKBD0 U6738 ( .CLK(n6855), .C(n6856) );
  CKBD0 U6739 ( .CLK(n6856), .C(n6857) );
  BUFFD0 U6740 ( .I(n6857), .Z(n6858) );
  CKBD0 U6741 ( .CLK(n6858), .C(n6859) );
  CKBD0 U6742 ( .CLK(n6859), .C(n6860) );
  CKBD0 U6743 ( .CLK(n6860), .C(n6861) );
  CKBD0 U6744 ( .CLK(n6861), .C(n6862) );
  CKBD0 U6745 ( .CLK(n6862), .C(n6863) );
  CKBD0 U6746 ( .CLK(n6863), .C(n6864) );
  CKBD0 U6747 ( .CLK(n6864), .C(n6865) );
  CKBD0 U6748 ( .CLK(n6865), .C(n6866) );
  CKBD0 U6749 ( .CLK(n6866), .C(n6867) );
  CKBD0 U6750 ( .CLK(n6867), .C(n6868) );
  BUFFD0 U6751 ( .I(n6868), .Z(n6869) );
  CKBD0 U6752 ( .CLK(n6869), .C(n6870) );
  CKBD0 U6753 ( .CLK(n6870), .C(n6871) );
  CKBD0 U6754 ( .CLK(n6871), .C(n6872) );
  CKBD0 U6755 ( .CLK(n6872), .C(n6873) );
  CKBD0 U6756 ( .CLK(n6873), .C(n6874) );
  CKBD0 U6757 ( .CLK(n6874), .C(n6875) );
  CKBD0 U6758 ( .CLK(n6875), .C(n6876) );
  CKBD0 U6759 ( .CLK(n6876), .C(n6877) );
  CKBD0 U6760 ( .CLK(n6877), .C(n6878) );
  BUFFD0 U6761 ( .I(n6878), .Z(n6879) );
  CKBD0 U6762 ( .CLK(n6879), .C(n6880) );
  CKBD0 U6763 ( .CLK(n6880), .C(n6881) );
  CKBD0 U6764 ( .CLK(n6881), .C(n6882) );
  CKBD0 U6765 ( .CLK(n6882), .C(n6883) );
  CKBD0 U6766 ( .CLK(n6883), .C(n6884) );
  CKBD0 U6767 ( .CLK(n6884), .C(n6885) );
  CKBD0 U6768 ( .CLK(n6885), .C(n6886) );
  CKBD0 U6769 ( .CLK(n6886), .C(n6887) );
  CKBD0 U6770 ( .CLK(n6887), .C(n6888) );
  CKBD0 U6771 ( .CLK(n6888), .C(n6889) );
  CKBD0 U6772 ( .CLK(n6889), .C(n6890) );
  BUFFD0 U6773 ( .I(n6890), .Z(n6891) );
  CKBD0 U6774 ( .CLK(n6891), .C(n6892) );
  CKBD0 U6775 ( .CLK(n6892), .C(n6893) );
  CKBD0 U6776 ( .CLK(n6893), .C(n6894) );
  CKBD0 U6777 ( .CLK(n6894), .C(n6895) );
  CKBD0 U6778 ( .CLK(n6895), .C(n6896) );
  CKBD0 U6779 ( .CLK(n6896), .C(n6897) );
  CKBD0 U6780 ( .CLK(n6897), .C(n6898) );
  CKBD0 U6781 ( .CLK(n6898), .C(n6899) );
  CKBD0 U6782 ( .CLK(n6899), .C(n6900) );
  BUFFD0 U6783 ( .I(n6900), .Z(n6901) );
  CKBD0 U6784 ( .CLK(n6901), .C(n6902) );
  CKBD0 U6785 ( .CLK(n6902), .C(n6903) );
  CKBD0 U6786 ( .CLK(n6903), .C(n6904) );
  CKBD0 U6787 ( .CLK(n6904), .C(n6905) );
  CKBD0 U6788 ( .CLK(n6905), .C(n6906) );
  CKBD0 U6789 ( .CLK(n6906), .C(n6907) );
  CKBD0 U6790 ( .CLK(n6907), .C(n6908) );
  CKBD0 U6791 ( .CLK(n6908), .C(n6909) );
  CKBD0 U6792 ( .CLK(n6909), .C(n6910) );
  CKBD0 U6793 ( .CLK(n6910), .C(n6911) );
  BUFFD0 U6794 ( .I(n6911), .Z(n6912) );
  CKBD0 U6795 ( .CLK(n6912), .C(n6913) );
  CKBD0 U6796 ( .CLK(n6913), .C(n6914) );
  CKBD0 U6797 ( .CLK(n6914), .C(n6915) );
  CKBD0 U6798 ( .CLK(n6915), .C(n6916) );
  CKBD0 U6799 ( .CLK(n6916), .C(n6917) );
  CKBD0 U6800 ( .CLK(n6917), .C(n6918) );
  CKBD0 U6801 ( .CLK(n6918), .C(n6919) );
  CKBD0 U6802 ( .CLK(n6919), .C(n6920) );
  CKBD0 U6803 ( .CLK(n6920), .C(n6921) );
  CKBD0 U6804 ( .CLK(n6921), .C(n6922) );
  BUFFD0 U6805 ( .I(n6922), .Z(n6923) );
  CKBD0 U6806 ( .CLK(n6923), .C(n6924) );
  CKBD0 U6807 ( .CLK(n6924), .C(n6925) );
  CKBD0 U6808 ( .CLK(n6925), .C(n6926) );
  CKBD0 U6809 ( .CLK(n6926), .C(n6927) );
  CKBD0 U6810 ( .CLK(n6927), .C(n6928) );
  CKBD0 U6811 ( .CLK(n6928), .C(n6929) );
  CKBD0 U6812 ( .CLK(n6929), .C(n6930) );
  CKBD0 U6813 ( .CLK(n6930), .C(n6931) );
  CKBD0 U6814 ( .CLK(n6931), .C(n6932) );
  CKBD0 U6815 ( .CLK(n6932), .C(n6933) );
  BUFFD0 U6816 ( .I(n6933), .Z(n6934) );
  CKBD0 U6817 ( .CLK(n6934), .C(n6935) );
  CKBD0 U6818 ( .CLK(n6935), .C(n6936) );
  CKBD0 U6819 ( .CLK(n6936), .C(n6937) );
  CKBD0 U6820 ( .CLK(n6937), .C(n6938) );
  CKBD0 U6821 ( .CLK(n6938), .C(n6939) );
  CKBD0 U6822 ( .CLK(n6939), .C(n6940) );
  CKBD0 U6823 ( .CLK(n6940), .C(n6941) );
  CKBD0 U6824 ( .CLK(n6941), .C(n6942) );
  CKBD0 U6825 ( .CLK(n6942), .C(n6943) );
  CKBD0 U6826 ( .CLK(n6943), .C(n6944) );
  BUFFD0 U6827 ( .I(n6944), .Z(n6945) );
  CKBD0 U6828 ( .CLK(n6945), .C(n6946) );
  CKBD0 U6829 ( .CLK(n6946), .C(n6947) );
  CKBD0 U6830 ( .CLK(n6947), .C(n6948) );
  CKBD0 U6831 ( .CLK(n6948), .C(n6949) );
  CKBD0 U6832 ( .CLK(n6949), .C(n6950) );
  BUFFD0 U6833 ( .I(n6950), .Z(n6951) );
  CKBD0 U6834 ( .CLK(n6951), .C(n6952) );
  BUFFD0 U6835 ( .I(n6952), .Z(n6953) );
  CKBD0 U6836 ( .CLK(n6953), .C(n6954) );
  BUFFD0 U6837 ( .I(n6954), .Z(n6955) );
  CKBD0 U6838 ( .CLK(n6955), .C(n6956) );
  BUFFD0 U6839 ( .I(n6956), .Z(n6957) );
  CKBD0 U6840 ( .CLK(n6957), .C(n6958) );
  BUFFD0 U6841 ( .I(n6958), .Z(n6959) );
  CKBD0 U6842 ( .CLK(n6959), .C(n6960) );
  BUFFD0 U6843 ( .I(n6960), .Z(n6961) );
  CKBD0 U6844 ( .CLK(n6961), .C(n6962) );
  BUFFD0 U6845 ( .I(n6962), .Z(n6963) );
  CKBD0 U6846 ( .CLK(n6963), .C(n6964) );
  BUFFD0 U6847 ( .I(n6964), .Z(n6965) );
  BUFFD0 U6848 ( .I(n6967), .Z(n6966) );
  BUFFD0 U6849 ( .I(n9233), .Z(n6967) );
  CKND2D0 U6850 ( .A1(n9165), .A2(ParValidTimer[0]), .ZN(n9288) );
  XOR2D0 U6851 ( .A1(n9020), .A2(n9288), .Z(n9287) );
  BUFFD0 U6852 ( .I(N39), .Z(n6968) );
  CKBD0 U6853 ( .CLK(Count32[0]), .C(n6977) );
  BUFFD0 U6854 ( .I(Count32[1]), .Z(n6969) );
  BUFFD0 U6855 ( .I(n9232), .Z(n6970) );
  BUFFD0 U6856 ( .I(n9286), .Z(n6971) );
  CKXOR2D0 U6857 ( .A1(n9165), .A2(n9292), .Z(n9286) );
  BUFFD0 U6858 ( .I(n6973), .Z(n6972) );
  BUFFD0 U6859 ( .I(N41), .Z(n6973) );
  BUFFD0 U6860 ( .I(n6975), .Z(n6974) );
  BUFFD0 U6861 ( .I(N40), .Z(n6975) );
  BUFFD0 U6862 ( .I(N38), .Z(n6976) );
  BUFFD0 U6863 ( .I(n6979), .Z(n6978) );
  BUFFD0 U6864 ( .I(n6980), .Z(n6979) );
  BUFFD0 U6865 ( .I(n6981), .Z(n6980) );
  BUFFD0 U6866 ( .I(n9202), .Z(n6981) );
  IOA22D0 U6867 ( .B1(n9127), .B2(n9239), .A1(n1), .A2(Decoder[2]), .ZN(n9202)
         );
  BUFFD0 U6868 ( .I(n6983), .Z(n6982) );
  BUFFD0 U6869 ( .I(n6984), .Z(n6983) );
  BUFFD0 U6870 ( .I(n6985), .Z(n6984) );
  BUFFD0 U6871 ( .I(n9201), .Z(n6985) );
  IOA22D0 U6872 ( .B1(n9127), .B2(n9238), .A1(n1), .A2(Decoder[1]), .ZN(n9201)
         );
  BUFFD0 U6873 ( .I(n6987), .Z(n6986) );
  BUFFD0 U6874 ( .I(N37), .Z(n6987) );
  BUFFD0 U6875 ( .I(n6989), .Z(n6988) );
  BUFFD0 U6876 ( .I(N43), .Z(n6989) );
  BUFFD0 U6877 ( .I(n6991), .Z(n6990) );
  BUFFD0 U6878 ( .I(n6992), .Z(n6991) );
  BUFFD0 U6879 ( .I(n6993), .Z(n6992) );
  BUFFD0 U6880 ( .I(n9200), .Z(n6993) );
  IOA22D0 U6881 ( .B1(n9128), .B2(n9237), .A1(n1), .A2(Decoder[0]), .ZN(n9200)
         );
  BUFFD0 U6882 ( .I(n6995), .Z(n6994) );
  BUFFD0 U6883 ( .I(n6996), .Z(n6995) );
  BUFFD0 U6884 ( .I(n6997), .Z(n6996) );
  BUFFD0 U6885 ( .I(n9205), .Z(n6997) );
  IOA22D0 U6886 ( .B1(n9127), .B2(n9242), .A1(n1), .A2(Decoder[5]), .ZN(n9205)
         );
  CKBD0 U6887 ( .CLK(n9212), .C(n7001) );
  BUFFD0 U6888 ( .I(n6999), .Z(n6998) );
  BUFFD0 U6889 ( .I(n7000), .Z(n6999) );
  BUFFD0 U6890 ( .I(n7001), .Z(n7000) );
  CKBD0 U6891 ( .CLK(n9219), .C(n7005) );
  BUFFD0 U6892 ( .I(n7003), .Z(n7002) );
  BUFFD0 U6893 ( .I(n7004), .Z(n7003) );
  BUFFD0 U6894 ( .I(n7005), .Z(n7004) );
  CKBD0 U6895 ( .CLK(n9206), .C(n7009) );
  MOAI22D1 U6896 ( .A1(n9127), .A2(n9243), .B1(n9129), .B2(Decoder[6]), .ZN(
        n9206) );
  BUFFD0 U6897 ( .I(n7007), .Z(n7006) );
  BUFFD0 U6898 ( .I(n7008), .Z(n7007) );
  BUFFD0 U6899 ( .I(n7009), .Z(n7008) );
  IOA22D4 U6900 ( .B1(n9127), .B2(n9246), .A1(n9129), .A2(Decoder[9]), .ZN(
        n9209) );
  BUFFD0 U6901 ( .I(n7011), .Z(n7010) );
  BUFFD0 U6902 ( .I(n7012), .Z(n7011) );
  BUFFD0 U6903 ( .I(n7013), .Z(n7012) );
  BUFFD0 U6904 ( .I(n9209), .Z(n7013) );
  IOA22D4 U6905 ( .B1(n9127), .B2(n9250), .A1(n9129), .A2(Decoder[13]), .ZN(
        n9213) );
  BUFFD0 U6906 ( .I(n7015), .Z(n7014) );
  BUFFD0 U6907 ( .I(n7016), .Z(n7015) );
  BUFFD0 U6908 ( .I(n7017), .Z(n7016) );
  BUFFD0 U6909 ( .I(n9213), .Z(n7017) );
  IOA22D4 U6910 ( .B1(n9128), .B2(n9253), .A1(n9129), .A2(Decoder[16]), .ZN(
        n9216) );
  BUFFD0 U6911 ( .I(n7019), .Z(n7018) );
  BUFFD0 U6912 ( .I(n7020), .Z(n7019) );
  BUFFD0 U6913 ( .I(n7021), .Z(n7020) );
  BUFFD0 U6914 ( .I(n9216), .Z(n7021) );
  IOA22D4 U6915 ( .B1(n9128), .B2(n9257), .A1(n9128), .A2(Decoder[20]), .ZN(
        n9220) );
  BUFFD0 U6916 ( .I(n7023), .Z(n7022) );
  BUFFD0 U6917 ( .I(n7024), .Z(n7023) );
  BUFFD0 U6918 ( .I(n7025), .Z(n7024) );
  BUFFD0 U6919 ( .I(n9220), .Z(n7025) );
  IOA22D4 U6920 ( .B1(n9128), .B2(n9260), .A1(n9129), .A2(Decoder[23]), .ZN(
        n9223) );
  BUFFD0 U6921 ( .I(n7027), .Z(n7026) );
  BUFFD0 U6922 ( .I(n7028), .Z(n7027) );
  BUFFD0 U6923 ( .I(n7029), .Z(n7028) );
  BUFFD0 U6924 ( .I(n9223), .Z(n7029) );
  IOA22D4 U6925 ( .B1(n9128), .B2(n9261), .A1(n9129), .A2(Decoder[24]), .ZN(
        n9224) );
  BUFFD0 U6926 ( .I(n7031), .Z(n7030) );
  BUFFD0 U6927 ( .I(n7032), .Z(n7031) );
  BUFFD0 U6928 ( .I(n7033), .Z(n7032) );
  BUFFD0 U6929 ( .I(n9224), .Z(n7033) );
  IOA22D4 U6930 ( .B1(n9128), .B2(n9264), .A1(n9129), .A2(Decoder[27]), .ZN(
        n9227) );
  BUFFD0 U6931 ( .I(n7035), .Z(n7034) );
  BUFFD0 U6932 ( .I(n7036), .Z(n7035) );
  BUFFD0 U6933 ( .I(n7037), .Z(n7036) );
  BUFFD0 U6934 ( .I(n9227), .Z(n7037) );
  IOA22D4 U6935 ( .B1(n9128), .B2(n9265), .A1(n1), .A2(Decoder[28]), .ZN(n9228) );
  BUFFD0 U6936 ( .I(n7039), .Z(n7038) );
  BUFFD0 U6937 ( .I(n7040), .Z(n7039) );
  BUFFD0 U6938 ( .I(n7041), .Z(n7040) );
  BUFFD0 U6939 ( .I(n9228), .Z(n7041) );
  BUFFD0 U6940 ( .I(n7043), .Z(n7042) );
  BUFFD0 U6941 ( .I(n7044), .Z(n7043) );
  BUFFD0 U6942 ( .I(n7045), .Z(n7044) );
  BUFFD0 U6943 ( .I(n9231), .Z(n7045) );
  BUFFD0 U6944 ( .I(n7047), .Z(n7046) );
  BUFFD0 U6945 ( .I(n7048), .Z(n7047) );
  BUFFD0 U6946 ( .I(n7049), .Z(n7048) );
  BUFFD0 U6947 ( .I(n9203), .Z(n7049) );
  IOA22D0 U6948 ( .B1(n9127), .B2(n9240), .A1(n1), .A2(Decoder[3]), .ZN(n9203)
         );
  BUFFD0 U6949 ( .I(n7051), .Z(n7050) );
  BUFFD0 U6950 ( .I(n7052), .Z(n7051) );
  BUFFD0 U6951 ( .I(n7053), .Z(n7052) );
  BUFFD0 U6952 ( .I(n9204), .Z(n7053) );
  IOA22D0 U6953 ( .B1(n9127), .B2(n9241), .A1(n1), .A2(Decoder[4]), .ZN(n9204)
         );
  IOA22D4 U6954 ( .B1(n9127), .B2(n9247), .A1(n9129), .A2(Decoder[10]), .ZN(
        n9210) );
  BUFFD0 U6955 ( .I(n7055), .Z(n7054) );
  BUFFD0 U6956 ( .I(n7056), .Z(n7055) );
  BUFFD0 U6957 ( .I(n7057), .Z(n7056) );
  BUFFD0 U6958 ( .I(n9210), .Z(n7057) );
  IOA22D4 U6959 ( .B1(n9127), .B2(n9248), .A1(n9129), .A2(Decoder[11]), .ZN(
        n9211) );
  BUFFD0 U6960 ( .I(n7059), .Z(n7058) );
  BUFFD0 U6961 ( .I(n7060), .Z(n7059) );
  BUFFD0 U6962 ( .I(n7061), .Z(n7060) );
  BUFFD0 U6963 ( .I(n9211), .Z(n7061) );
  IOA22D4 U6964 ( .B1(n9128), .B2(n9254), .A1(n9129), .A2(Decoder[17]), .ZN(
        n9217) );
  BUFFD0 U6965 ( .I(n7063), .Z(n7062) );
  BUFFD0 U6966 ( .I(n7064), .Z(n7063) );
  BUFFD0 U6967 ( .I(n7065), .Z(n7064) );
  BUFFD0 U6968 ( .I(n9217), .Z(n7065) );
  IOA22D4 U6969 ( .B1(n9128), .B2(n9255), .A1(n9129), .A2(Decoder[18]), .ZN(
        n9218) );
  BUFFD0 U6970 ( .I(n7067), .Z(n7066) );
  BUFFD0 U6971 ( .I(n7068), .Z(n7067) );
  BUFFD0 U6972 ( .I(n7069), .Z(n7068) );
  BUFFD0 U6973 ( .I(n9218), .Z(n7069) );
  IOA22D4 U6974 ( .B1(n9127), .B2(n9244), .A1(n1), .A2(Decoder[7]), .ZN(n9207)
         );
  BUFFD0 U6975 ( .I(n7071), .Z(n7070) );
  BUFFD0 U6976 ( .I(n7072), .Z(n7071) );
  BUFFD0 U6977 ( .I(n7073), .Z(n7072) );
  BUFFD0 U6978 ( .I(n9207), .Z(n7073) );
  IOA22D4 U6979 ( .B1(n9127), .B2(n9245), .A1(n9129), .A2(Decoder[8]), .ZN(
        n9208) );
  BUFFD0 U6980 ( .I(n7075), .Z(n7074) );
  BUFFD0 U6981 ( .I(n7076), .Z(n7075) );
  BUFFD0 U6982 ( .I(n7077), .Z(n7076) );
  BUFFD0 U6983 ( .I(n9208), .Z(n7077) );
  IOA22D4 U6984 ( .B1(n9128), .B2(n9251), .A1(n9129), .A2(Decoder[14]), .ZN(
        n9214) );
  BUFFD0 U6985 ( .I(n7079), .Z(n7078) );
  BUFFD0 U6986 ( .I(n7080), .Z(n7079) );
  BUFFD0 U6987 ( .I(n7081), .Z(n7080) );
  BUFFD0 U6988 ( .I(n9214), .Z(n7081) );
  IOA22D4 U6989 ( .B1(n9128), .B2(n9252), .A1(n9129), .A2(Decoder[15]), .ZN(
        n9215) );
  BUFFD0 U6990 ( .I(n7083), .Z(n7082) );
  BUFFD0 U6991 ( .I(n7084), .Z(n7083) );
  BUFFD0 U6992 ( .I(n7085), .Z(n7084) );
  BUFFD0 U6993 ( .I(n9215), .Z(n7085) );
  IOA22D4 U6994 ( .B1(n9128), .B2(n9258), .A1(n9129), .A2(Decoder[21]), .ZN(
        n9221) );
  BUFFD0 U6995 ( .I(n7087), .Z(n7086) );
  BUFFD0 U6996 ( .I(n7088), .Z(n7087) );
  BUFFD0 U6997 ( .I(n7089), .Z(n7088) );
  BUFFD0 U6998 ( .I(n9221), .Z(n7089) );
  IOA22D4 U6999 ( .B1(n9128), .B2(n9259), .A1(n9129), .A2(Decoder[22]), .ZN(
        n9222) );
  BUFFD0 U7000 ( .I(n7091), .Z(n7090) );
  BUFFD0 U7001 ( .I(n7092), .Z(n7091) );
  BUFFD0 U7002 ( .I(n7093), .Z(n7092) );
  BUFFD0 U7003 ( .I(n9222), .Z(n7093) );
  IOA22D4 U7004 ( .B1(n9128), .B2(n9262), .A1(n9129), .A2(Decoder[25]), .ZN(
        n9225) );
  BUFFD0 U7005 ( .I(n7095), .Z(n7094) );
  BUFFD0 U7006 ( .I(n7096), .Z(n7095) );
  BUFFD0 U7007 ( .I(n7097), .Z(n7096) );
  BUFFD0 U7008 ( .I(n9225), .Z(n7097) );
  IOA22D4 U7009 ( .B1(n9128), .B2(n9263), .A1(n9129), .A2(Decoder[26]), .ZN(
        n9226) );
  BUFFD0 U7010 ( .I(n7099), .Z(n7098) );
  BUFFD0 U7011 ( .I(n7100), .Z(n7099) );
  BUFFD0 U7012 ( .I(n7101), .Z(n7100) );
  BUFFD0 U7013 ( .I(n9226), .Z(n7101) );
  IOA22D4 U7014 ( .B1(n9128), .B2(n9266), .A1(n1), .A2(Decoder[29]), .ZN(n9229) );
  BUFFD0 U7015 ( .I(n7103), .Z(n7102) );
  BUFFD0 U7016 ( .I(n7104), .Z(n7103) );
  BUFFD0 U7017 ( .I(n7105), .Z(n7104) );
  BUFFD0 U7018 ( .I(n9229), .Z(n7105) );
  IOA22D4 U7019 ( .B1(n9128), .B2(n9267), .A1(n1), .A2(Decoder[30]), .ZN(n9230) );
  BUFFD0 U7020 ( .I(n7107), .Z(n7106) );
  BUFFD0 U7021 ( .I(n7108), .Z(n7107) );
  BUFFD0 U7022 ( .I(n7109), .Z(n7108) );
  BUFFD0 U7023 ( .I(n9230), .Z(n7109) );
  OAI21D0 U7024 ( .A1(n9293), .A2(n9269), .B(n9166), .ZN(n9236) );
  BUFFD0 U7025 ( .I(n7111), .Z(n7110) );
  BUFFD0 U7026 ( .I(n7112), .Z(n7111) );
  BUFFD0 U7027 ( .I(n7113), .Z(n7112) );
  BUFFD0 U7028 ( .I(n9236), .Z(n7113) );
  NR2D0 U7029 ( .A1(n9283), .A2(n9284), .ZN(N47) );
  CKBD0 U7030 ( .CLK(n1900), .C(n7114) );
  CKBD0 U7031 ( .CLK(n1692), .C(n7115) );
  CKBD0 U7032 ( .CLK(n1906), .C(n7116) );
  CKBD0 U7033 ( .CLK(n1696), .C(n7117) );
  CKBD0 U7034 ( .CLK(n1903), .C(n7118) );
  CKBD0 U7035 ( .CLK(n1910), .C(n7119) );
  CKBD0 U7036 ( .CLK(n2207), .C(n7120) );
  CKBD0 U7037 ( .CLK(n2108), .C(n7121) );
  CKBD0 U7038 ( .CLK(n2306), .C(n7122) );
  CKBD0 U7039 ( .CLK(n1392), .C(n7123) );
  CKBD0 U7040 ( .CLK(n1689), .C(n7124) );
  CKBD0 U7041 ( .CLK(n2009), .C(n7125) );
  CKBD0 U7042 ( .CLK(n2405), .C(n7126) );
  CKBD0 U7043 ( .CLK(n1377), .C(n7127) );
  CKBD0 U7044 ( .CLK(n1263), .C(n7128) );
  CKBD0 U7045 ( .CLK(n936), .C(n7129) );
  CKBD0 U7046 ( .CLK(n932), .C(n7130) );
  BUFFD0 U7047 ( .I(n229), .Z(n7131) );
  CKBD0 U7048 ( .CLK(n1590), .C(n7132) );
  CKBD0 U7049 ( .CLK(n1895), .C(n7133) );
  CKBD0 U7050 ( .CLK(n832), .C(n7134) );
  BUFFD0 U7051 ( .I(n1049), .Z(n7135) );
  CKBD0 U7052 ( .CLK(n1149), .C(n7136) );
  BUFFD0 U7053 ( .I(n1795), .Z(n7137) );
  BUFFD0 U7054 ( .I(n730), .Z(n7138) );
  CKBD0 U7055 ( .CLK(n531), .C(n7139) );
  CKBD0 U7056 ( .CLK(n431), .C(n7140) );
  BUFFD0 U7057 ( .I(n2603), .Z(n7141) );
  CKBD0 U7058 ( .CLK(n332), .C(n7142) );
  CKBD0 U7059 ( .CLK(n630), .C(n7143) );
  CKBD0 U7060 ( .CLK(n2504), .C(n7144) );
  CKBD0 U7061 ( .CLK(n1491), .C(n7145) );
  CKBD0 U7062 ( .CLK(n7114), .C(n7146) );
  CKBD0 U7063 ( .CLK(n7115), .C(n7147) );
  CKBD0 U7064 ( .CLK(n7116), .C(n7148) );
  CKBD0 U7065 ( .CLK(n7117), .C(n7149) );
  CKBD0 U7066 ( .CLK(n7118), .C(n7150) );
  CKBD0 U7067 ( .CLK(n7119), .C(n7151) );
  CKBD0 U7068 ( .CLK(n7120), .C(n7152) );
  CKBD0 U7069 ( .CLK(n7121), .C(n7153) );
  CKBD0 U7070 ( .CLK(n7122), .C(n7154) );
  CKBD0 U7071 ( .CLK(n7123), .C(n7155) );
  CKBD0 U7072 ( .CLK(n7124), .C(n7156) );
  CKBD0 U7073 ( .CLK(n7125), .C(n7157) );
  CKBD0 U7074 ( .CLK(n7126), .C(n7158) );
  CKBD0 U7075 ( .CLK(n7127), .C(n7159) );
  CKBD0 U7076 ( .CLK(n7128), .C(n7160) );
  CKBD0 U7077 ( .CLK(n7130), .C(n7161) );
  CKBD0 U7078 ( .CLK(n7129), .C(n7162) );
  CKBD0 U7079 ( .CLK(n7131), .C(n7163) );
  CKBD0 U7080 ( .CLK(n7132), .C(n7164) );
  CKBD0 U7081 ( .CLK(n7133), .C(n7165) );
  CKBD0 U7082 ( .CLK(n7134), .C(n7166) );
  CKBD0 U7083 ( .CLK(n7135), .C(n7167) );
  CKBD0 U7084 ( .CLK(n7136), .C(n7168) );
  CKBD0 U7085 ( .CLK(n7137), .C(n7169) );
  CKBD0 U7086 ( .CLK(n7138), .C(n7170) );
  CKBD0 U7087 ( .CLK(n7139), .C(n7171) );
  CKBD0 U7088 ( .CLK(n7140), .C(n7172) );
  CKBD0 U7089 ( .CLK(n7141), .C(n7173) );
  CKBD0 U7090 ( .CLK(n7142), .C(n7174) );
  CKBD0 U7091 ( .CLK(n7143), .C(n7175) );
  CKBD0 U7092 ( .CLK(n7144), .C(n7176) );
  CKBD0 U7093 ( .CLK(n7145), .C(n7177) );
  CKBD0 U7094 ( .CLK(n7146), .C(n7178) );
  CKBD0 U7095 ( .CLK(n7147), .C(n7179) );
  CKBD0 U7096 ( .CLK(n7148), .C(n7180) );
  CKBD0 U7097 ( .CLK(n7149), .C(n7181) );
  CKBD0 U7098 ( .CLK(n7150), .C(n7182) );
  CKBD0 U7099 ( .CLK(n7151), .C(n7183) );
  CKBD0 U7100 ( .CLK(n7152), .C(n7184) );
  BUFFD0 U7101 ( .I(n7155), .Z(n7185) );
  CKBD0 U7102 ( .CLK(n7153), .C(n7186) );
  CKBD0 U7103 ( .CLK(n7154), .C(n7187) );
  BUFFD0 U7104 ( .I(n7156), .Z(n7188) );
  CKBD0 U7105 ( .CLK(n7157), .C(n7189) );
  CKBD0 U7106 ( .CLK(n7158), .C(n7190) );
  CKBD0 U7107 ( .CLK(n7159), .C(n7191) );
  CKBD0 U7108 ( .CLK(n7160), .C(n7192) );
  CKBD0 U7109 ( .CLK(n7161), .C(n7193) );
  CKBD0 U7110 ( .CLK(n7162), .C(n7194) );
  CKBD0 U7111 ( .CLK(n7163), .C(n7195) );
  CKBD0 U7112 ( .CLK(n7164), .C(n7196) );
  CKBD0 U7113 ( .CLK(n7165), .C(n7197) );
  CKBD0 U7114 ( .CLK(n7166), .C(n7198) );
  CKBD0 U7115 ( .CLK(n7167), .C(n7199) );
  CKBD0 U7116 ( .CLK(n7168), .C(n7200) );
  CKBD0 U7117 ( .CLK(n7169), .C(n7201) );
  CKBD0 U7118 ( .CLK(n7170), .C(n7202) );
  CKBD0 U7119 ( .CLK(n7171), .C(n7203) );
  CKBD0 U7120 ( .CLK(n7173), .C(n7204) );
  CKBD0 U7121 ( .CLK(n7174), .C(n7205) );
  CKBD0 U7122 ( .CLK(n7172), .C(n7206) );
  CKBD0 U7123 ( .CLK(n7175), .C(n7207) );
  CKBD0 U7124 ( .CLK(n7176), .C(n7208) );
  CKBD0 U7125 ( .CLK(n7177), .C(n7209) );
  CKBD0 U7126 ( .CLK(n7178), .C(n7210) );
  CKBD0 U7127 ( .CLK(n7179), .C(n7211) );
  CKBD0 U7128 ( .CLK(n7180), .C(n7212) );
  CKBD0 U7129 ( .CLK(n7181), .C(n7213) );
  CKBD0 U7130 ( .CLK(n7182), .C(n7214) );
  CKBD0 U7131 ( .CLK(n7183), .C(n7215) );
  CKBD0 U7132 ( .CLK(n7184), .C(n7216) );
  CKBD0 U7133 ( .CLK(n7185), .C(n7217) );
  CKBD0 U7134 ( .CLK(n7186), .C(n7218) );
  CKBD0 U7135 ( .CLK(n7187), .C(n7219) );
  CKBD0 U7136 ( .CLK(n7188), .C(n7220) );
  CKBD0 U7137 ( .CLK(n7189), .C(n7221) );
  CKBD0 U7138 ( .CLK(n7190), .C(n7222) );
  CKBD0 U7139 ( .CLK(n7191), .C(n7223) );
  BUFFD0 U7140 ( .I(n7192), .Z(n7224) );
  CKBD0 U7141 ( .CLK(n7193), .C(n7225) );
  CKBD0 U7142 ( .CLK(n7195), .C(n7226) );
  CKBD0 U7143 ( .CLK(n7194), .C(n7227) );
  CKBD0 U7144 ( .CLK(n7196), .C(n7228) );
  CKBD0 U7145 ( .CLK(n7197), .C(n7229) );
  CKBD0 U7146 ( .CLK(n7198), .C(n7230) );
  CKBD0 U7147 ( .CLK(n7199), .C(n7231) );
  CKBD0 U7148 ( .CLK(n7200), .C(n7232) );
  CKBD0 U7149 ( .CLK(n7201), .C(n7233) );
  CKBD0 U7150 ( .CLK(n7202), .C(n7234) );
  CKBD0 U7151 ( .CLK(n7203), .C(n7235) );
  CKBD0 U7152 ( .CLK(n7205), .C(n7236) );
  CKBD0 U7153 ( .CLK(n7204), .C(n7237) );
  CKBD0 U7154 ( .CLK(n7206), .C(n7238) );
  CKBD0 U7155 ( .CLK(n7207), .C(n7239) );
  BUFFD0 U7156 ( .I(n7210), .Z(n7240) );
  CKBD0 U7157 ( .CLK(n7208), .C(n7241) );
  CKBD0 U7158 ( .CLK(n7209), .C(n7242) );
  CKBD0 U7159 ( .CLK(n7211), .C(n7243) );
  CKBD0 U7160 ( .CLK(n7212), .C(n7244) );
  CKBD0 U7161 ( .CLK(n7213), .C(n7245) );
  BUFFD0 U7162 ( .I(n7214), .Z(n7246) );
  CKBD0 U7163 ( .CLK(n7215), .C(n7247) );
  CKBD0 U7164 ( .CLK(n7216), .C(n7248) );
  CKBD0 U7165 ( .CLK(n7218), .C(n7249) );
  CKBD0 U7166 ( .CLK(n7217), .C(n7250) );
  CKBD0 U7167 ( .CLK(n7219), .C(n7251) );
  CKBD0 U7168 ( .CLK(n7220), .C(n7252) );
  CKBD0 U7169 ( .CLK(n7221), .C(n7253) );
  CKBD0 U7170 ( .CLK(n7222), .C(n7254) );
  CKBD0 U7171 ( .CLK(n7223), .C(n7255) );
  CKBD0 U7172 ( .CLK(n7224), .C(n7256) );
  CKBD0 U7173 ( .CLK(n7225), .C(n7257) );
  CKBD0 U7174 ( .CLK(n7229), .C(n7258) );
  CKBD0 U7175 ( .CLK(n7227), .C(n7259) );
  CKBD0 U7176 ( .CLK(n7226), .C(n7260) );
  CKBD0 U7177 ( .CLK(n7228), .C(n7261) );
  CKBD0 U7178 ( .CLK(n7230), .C(n7262) );
  CKBD0 U7179 ( .CLK(n7231), .C(n7263) );
  CKBD0 U7180 ( .CLK(n7232), .C(n7264) );
  CKBD0 U7181 ( .CLK(n7233), .C(n7265) );
  CKBD0 U7182 ( .CLK(n7234), .C(n7266) );
  CKBD0 U7183 ( .CLK(n7235), .C(n7267) );
  BUFFD0 U7184 ( .I(n7236), .Z(n7268) );
  CKBD0 U7185 ( .CLK(n7237), .C(n7269) );
  CKBD0 U7186 ( .CLK(n7238), .C(n7270) );
  CKBD0 U7187 ( .CLK(n7239), .C(n7271) );
  CKBD0 U7188 ( .CLK(n7240), .C(n7272) );
  CKBD0 U7189 ( .CLK(n7241), .C(n7273) );
  CKBD0 U7190 ( .CLK(n7242), .C(n7274) );
  BUFFD0 U7191 ( .I(n7243), .Z(n7275) );
  BUFFD0 U7192 ( .I(n7244), .Z(n7276) );
  CKBD0 U7193 ( .CLK(n7245), .C(n7277) );
  CKBD0 U7194 ( .CLK(n7246), .C(n7278) );
  CKBD0 U7195 ( .CLK(n7247), .C(n7279) );
  CKBD0 U7196 ( .CLK(n7248), .C(n7280) );
  BUFFD0 U7197 ( .I(n7249), .Z(n7281) );
  BUFFD0 U7198 ( .I(n7251), .Z(n7282) );
  CKBD0 U7199 ( .CLK(n7250), .C(n7283) );
  CKBD0 U7200 ( .CLK(n7253), .C(n7284) );
  CKBD0 U7201 ( .CLK(n7252), .C(n7285) );
  CKBD0 U7202 ( .CLK(n7254), .C(n7286) );
  CKBD0 U7203 ( .CLK(n7255), .C(n7287) );
  BUFFD0 U7204 ( .I(n7259), .Z(n7288) );
  CKBD0 U7205 ( .CLK(n7256), .C(n7289) );
  CKBD0 U7206 ( .CLK(n7257), .C(n7290) );
  BUFFD0 U7207 ( .I(n7258), .Z(n7291) );
  CKBD0 U7208 ( .CLK(n7260), .C(n7292) );
  CKBD0 U7209 ( .CLK(n7261), .C(n7293) );
  CKBD0 U7210 ( .CLK(n7262), .C(n7294) );
  CKBD0 U7211 ( .CLK(n7264), .C(n7295) );
  CKBD0 U7212 ( .CLK(n7263), .C(n7296) );
  CKBD0 U7213 ( .CLK(n7265), .C(n7297) );
  CKBD0 U7214 ( .CLK(n7266), .C(n7298) );
  CKBD0 U7215 ( .CLK(n7267), .C(n7299) );
  CKBD0 U7216 ( .CLK(n7268), .C(n7300) );
  CKBD0 U7217 ( .CLK(n7269), .C(n7301) );
  CKBD0 U7218 ( .CLK(n7270), .C(n7302) );
  CKBD0 U7219 ( .CLK(n7271), .C(n7303) );
  CKBD0 U7220 ( .CLK(n7272), .C(n7304) );
  CKBD0 U7221 ( .CLK(n7273), .C(n7305) );
  CKBD0 U7222 ( .CLK(n7274), .C(n7306) );
  CKBD0 U7223 ( .CLK(n7275), .C(n7307) );
  CKBD0 U7224 ( .CLK(n7276), .C(n7308) );
  BUFFD0 U7225 ( .I(n7277), .Z(n7309) );
  CKBD0 U7226 ( .CLK(n7278), .C(n7310) );
  CKBD0 U7227 ( .CLK(n7279), .C(n7311) );
  CKBD0 U7228 ( .CLK(n7280), .C(n7312) );
  CKBD0 U7229 ( .CLK(n7281), .C(n7313) );
  CKBD0 U7230 ( .CLK(n7282), .C(n7314) );
  CKBD0 U7231 ( .CLK(n7283), .C(n7315) );
  CKBD0 U7232 ( .CLK(n7285), .C(n7316) );
  BUFFD0 U7233 ( .I(n7284), .Z(n7317) );
  CKBD0 U7234 ( .CLK(n7286), .C(n7318) );
  CKBD0 U7235 ( .CLK(n7287), .C(n7319) );
  CKBD0 U7236 ( .CLK(n7289), .C(n7320) );
  CKBD0 U7237 ( .CLK(n7288), .C(n7321) );
  CKBD0 U7238 ( .CLK(n7290), .C(n7322) );
  CKBD0 U7239 ( .CLK(n7291), .C(n7323) );
  CKBD0 U7240 ( .CLK(n7292), .C(n7324) );
  CKBD0 U7241 ( .CLK(n7293), .C(n7325) );
  BUFFD0 U7242 ( .I(n7294), .Z(n7326) );
  BUFFD0 U7243 ( .I(n7295), .Z(n7327) );
  CKBD0 U7244 ( .CLK(n7296), .C(n7328) );
  CKBD0 U7245 ( .CLK(n7297), .C(n7329) );
  CKBD0 U7246 ( .CLK(n7298), .C(n7330) );
  CKBD0 U7247 ( .CLK(n7299), .C(n7331) );
  CKBD0 U7248 ( .CLK(n7300), .C(n7332) );
  CKBD0 U7249 ( .CLK(n7301), .C(n7333) );
  CKBD0 U7250 ( .CLK(n7302), .C(n7334) );
  CKBD0 U7251 ( .CLK(n7303), .C(n7335) );
  CKBD0 U7252 ( .CLK(n7304), .C(n7336) );
  CKBD0 U7253 ( .CLK(n7305), .C(n7337) );
  CKBD0 U7254 ( .CLK(n7306), .C(n7338) );
  CKBD0 U7255 ( .CLK(n7307), .C(n7339) );
  CKBD0 U7256 ( .CLK(n7308), .C(n7340) );
  CKBD0 U7257 ( .CLK(n7309), .C(n7341) );
  CKBD0 U7258 ( .CLK(n7310), .C(n7342) );
  BUFFD0 U7259 ( .I(n7311), .Z(n7343) );
  BUFFD0 U7260 ( .I(n7312), .Z(n7344) );
  CKBD0 U7261 ( .CLK(n7313), .C(n7345) );
  CKBD0 U7262 ( .CLK(n7314), .C(n7346) );
  CKBD0 U7263 ( .CLK(n7315), .C(n7347) );
  CKBD0 U7264 ( .CLK(n7316), .C(n7348) );
  CKBD0 U7265 ( .CLK(n7317), .C(n7349) );
  CKBD0 U7266 ( .CLK(n7318), .C(n7350) );
  CKBD0 U7267 ( .CLK(n7319), .C(n7351) );
  CKBD0 U7268 ( .CLK(n7320), .C(n7352) );
  CKBD0 U7269 ( .CLK(n7321), .C(n7353) );
  CKBD0 U7270 ( .CLK(n7322), .C(n7354) );
  CKBD0 U7271 ( .CLK(n7323), .C(n7355) );
  CKBD0 U7272 ( .CLK(n7324), .C(n7356) );
  CKBD0 U7273 ( .CLK(n7325), .C(n7357) );
  CKBD0 U7274 ( .CLK(n7326), .C(n7358) );
  CKBD0 U7275 ( .CLK(n7327), .C(n7359) );
  CKBD0 U7276 ( .CLK(n7328), .C(n7360) );
  CKBD0 U7277 ( .CLK(n7329), .C(n7361) );
  CKBD0 U7278 ( .CLK(n7330), .C(n7362) );
  CKBD0 U7279 ( .CLK(n7331), .C(n7363) );
  CKBD0 U7280 ( .CLK(n7332), .C(n7364) );
  CKBD0 U7281 ( .CLK(n7333), .C(n7365) );
  CKBD0 U7282 ( .CLK(n7334), .C(n7366) );
  CKBD0 U7283 ( .CLK(n7335), .C(n7367) );
  CKBD0 U7284 ( .CLK(n7336), .C(n7368) );
  CKBD0 U7285 ( .CLK(n7337), .C(n7369) );
  CKBD0 U7286 ( .CLK(n7338), .C(n7370) );
  CKBD0 U7287 ( .CLK(n7339), .C(n7371) );
  CKBD0 U7288 ( .CLK(n7340), .C(n7372) );
  CKBD0 U7289 ( .CLK(n7341), .C(n7373) );
  CKBD0 U7290 ( .CLK(n7342), .C(n7374) );
  CKBD0 U7291 ( .CLK(n7343), .C(n7375) );
  CKBD0 U7292 ( .CLK(n7344), .C(n7376) );
  CKBD0 U7293 ( .CLK(n7345), .C(n7377) );
  CKBD0 U7294 ( .CLK(n7346), .C(n7378) );
  CKBD0 U7295 ( .CLK(n7347), .C(n7379) );
  CKBD0 U7296 ( .CLK(n7348), .C(n7380) );
  CKBD0 U7297 ( .CLK(n7349), .C(n7381) );
  CKBD0 U7298 ( .CLK(n7351), .C(n7382) );
  BUFFD0 U7299 ( .I(n7350), .Z(n7383) );
  CKBD0 U7300 ( .CLK(n7352), .C(n7384) );
  CKBD0 U7301 ( .CLK(n7353), .C(n7385) );
  BUFFD0 U7302 ( .I(n7354), .Z(n7386) );
  CKBD0 U7303 ( .CLK(n7357), .C(n7387) );
  CKBD0 U7304 ( .CLK(n7355), .C(n7388) );
  CKBD0 U7305 ( .CLK(n7356), .C(n7389) );
  CKBD0 U7306 ( .CLK(n7358), .C(n7390) );
  CKBD0 U7307 ( .CLK(n7359), .C(n7391) );
  CKBD0 U7308 ( .CLK(n7360), .C(n7392) );
  CKBD0 U7309 ( .CLK(n7361), .C(n7393) );
  CKBD0 U7310 ( .CLK(n7362), .C(n7394) );
  CKBD0 U7311 ( .CLK(n7363), .C(n7395) );
  CKBD0 U7312 ( .CLK(n7364), .C(n7396) );
  CKBD0 U7313 ( .CLK(n7365), .C(n7397) );
  BUFFD0 U7314 ( .I(n7367), .Z(n7398) );
  CKBD0 U7315 ( .CLK(n7366), .C(n7399) );
  BUFFD0 U7316 ( .I(n7369), .Z(n7400) );
  CKBD0 U7317 ( .CLK(n7368), .C(n7401) );
  CKBD0 U7318 ( .CLK(n7370), .C(n7402) );
  CKBD0 U7319 ( .CLK(n7371), .C(n7403) );
  CKBD0 U7320 ( .CLK(n7372), .C(n7404) );
  CKBD0 U7321 ( .CLK(n7373), .C(n7405) );
  CKBD0 U7322 ( .CLK(n7374), .C(n7406) );
  CKBD0 U7323 ( .CLK(n7375), .C(n7407) );
  CKBD0 U7324 ( .CLK(n7376), .C(n7408) );
  CKBD0 U7325 ( .CLK(n7377), .C(n7409) );
  CKBD0 U7326 ( .CLK(n7378), .C(n7410) );
  CKBD0 U7327 ( .CLK(n7379), .C(n7411) );
  CKBD0 U7328 ( .CLK(n7380), .C(n7412) );
  CKBD0 U7329 ( .CLK(n7381), .C(n7413) );
  CKBD0 U7330 ( .CLK(n7383), .C(n7414) );
  BUFFD0 U7331 ( .I(n7382), .Z(n7415) );
  CKBD0 U7332 ( .CLK(n7384), .C(n7416) );
  CKBD0 U7333 ( .CLK(n7385), .C(n7417) );
  CKBD0 U7334 ( .CLK(n7386), .C(n7418) );
  BUFFD0 U7335 ( .I(n7387), .Z(n7419) );
  CKBD0 U7336 ( .CLK(n7388), .C(n7420) );
  CKBD0 U7337 ( .CLK(n7389), .C(n7421) );
  CKBD0 U7338 ( .CLK(n7390), .C(n7422) );
  CKBD0 U7339 ( .CLK(n7391), .C(n7423) );
  CKBD0 U7340 ( .CLK(n7392), .C(n7424) );
  CKBD0 U7341 ( .CLK(n7393), .C(n7425) );
  CKBD0 U7342 ( .CLK(n7394), .C(n7426) );
  BUFFD0 U7343 ( .I(n7395), .Z(n7427) );
  CKBD0 U7344 ( .CLK(n7397), .C(n7428) );
  CKBD0 U7345 ( .CLK(n7396), .C(n7429) );
  CKBD0 U7346 ( .CLK(n7398), .C(n7430) );
  CKBD0 U7347 ( .CLK(n7399), .C(n7431) );
  CKBD0 U7348 ( .CLK(n7400), .C(n7432) );
  BUFFD0 U7349 ( .I(n7402), .Z(n7433) );
  CKBD0 U7350 ( .CLK(n7401), .C(n7434) );
  CKBD0 U7351 ( .CLK(n7403), .C(n7435) );
  CKBD0 U7352 ( .CLK(n7404), .C(n7436) );
  CKBD0 U7353 ( .CLK(n7405), .C(n7437) );
  CKBD0 U7354 ( .CLK(n7406), .C(n7438) );
  CKBD0 U7355 ( .CLK(n7407), .C(n7439) );
  CKBD0 U7356 ( .CLK(n7408), .C(n7440) );
  CKBD0 U7357 ( .CLK(n7409), .C(n7441) );
  CKBD0 U7358 ( .CLK(n7410), .C(n7442) );
  CKBD0 U7359 ( .CLK(n7411), .C(n7443) );
  CKBD0 U7360 ( .CLK(n7412), .C(n7444) );
  CKBD0 U7361 ( .CLK(n7413), .C(n7445) );
  CKBD0 U7362 ( .CLK(n7414), .C(n7446) );
  CKBD0 U7363 ( .CLK(n7415), .C(n7447) );
  CKBD0 U7364 ( .CLK(n7416), .C(n7448) );
  CKBD0 U7365 ( .CLK(n7417), .C(n7449) );
  CKBD0 U7366 ( .CLK(n7418), .C(n7450) );
  CKBD0 U7367 ( .CLK(n7421), .C(n7451) );
  CKBD0 U7368 ( .CLK(n7419), .C(n7452) );
  CKBD0 U7369 ( .CLK(n7420), .C(n7453) );
  CKBD0 U7370 ( .CLK(n7422), .C(n7454) );
  CKBD0 U7371 ( .CLK(n7424), .C(n7455) );
  CKBD0 U7372 ( .CLK(n7423), .C(n7456) );
  BUFFD0 U7373 ( .I(n7425), .Z(n7457) );
  CKBD0 U7374 ( .CLK(n7426), .C(n7458) );
  CKBD0 U7375 ( .CLK(n7427), .C(n7459) );
  BUFFD0 U7376 ( .I(n7428), .Z(n7460) );
  CKBD0 U7377 ( .CLK(n7429), .C(n7461) );
  CKBD0 U7378 ( .CLK(n7430), .C(n7462) );
  CKBD0 U7379 ( .CLK(n7431), .C(n7463) );
  CKBD0 U7380 ( .CLK(n7432), .C(n7464) );
  CKBD0 U7381 ( .CLK(n7433), .C(n7465) );
  CKBD0 U7382 ( .CLK(n7434), .C(n7466) );
  CKBD0 U7383 ( .CLK(n7435), .C(n7467) );
  CKBD0 U7384 ( .CLK(n7436), .C(n7468) );
  CKBD0 U7385 ( .CLK(n7437), .C(n7469) );
  CKBD0 U7386 ( .CLK(n7438), .C(n7470) );
  CKBD0 U7387 ( .CLK(n7439), .C(n7471) );
  CKBD0 U7388 ( .CLK(n7440), .C(n7472) );
  CKBD0 U7389 ( .CLK(n7441), .C(n7473) );
  CKBD0 U7390 ( .CLK(n7442), .C(n7474) );
  CKBD0 U7391 ( .CLK(n7443), .C(n7475) );
  CKBD0 U7392 ( .CLK(n7444), .C(n7476) );
  CKBD0 U7393 ( .CLK(n7445), .C(n7477) );
  CKBD0 U7394 ( .CLK(n7446), .C(n7478) );
  CKBD0 U7395 ( .CLK(n7447), .C(n7479) );
  CKBD0 U7396 ( .CLK(n7448), .C(n7480) );
  CKBD0 U7397 ( .CLK(n7449), .C(n7481) );
  CKBD0 U7398 ( .CLK(n7450), .C(n7482) );
  BUFFD0 U7399 ( .I(n7451), .Z(n7483) );
  CKBD0 U7400 ( .CLK(n7452), .C(n7484) );
  CKBD0 U7401 ( .CLK(n7453), .C(n7485) );
  CKBD0 U7402 ( .CLK(n7454), .C(n7486) );
  BUFFD0 U7403 ( .I(n7455), .Z(n7487) );
  CKBD0 U7404 ( .CLK(n7456), .C(n7488) );
  CKBD0 U7405 ( .CLK(n7457), .C(n7489) );
  CKBD0 U7406 ( .CLK(n7458), .C(n7490) );
  CKBD0 U7407 ( .CLK(n7459), .C(n7491) );
  CKBD0 U7408 ( .CLK(n7460), .C(n7492) );
  CKBD0 U7409 ( .CLK(n7461), .C(n7493) );
  CKBD0 U7410 ( .CLK(n7462), .C(n7494) );
  CKBD0 U7411 ( .CLK(n7463), .C(n7495) );
  CKBD0 U7412 ( .CLK(n7464), .C(n7496) );
  CKBD0 U7413 ( .CLK(n7465), .C(n7497) );
  CKBD0 U7414 ( .CLK(n7466), .C(n7498) );
  CKBD0 U7415 ( .CLK(n7467), .C(n7499) );
  CKBD0 U7416 ( .CLK(n7468), .C(n7500) );
  CKBD0 U7417 ( .CLK(n7469), .C(n7501) );
  CKBD0 U7418 ( .CLK(n7470), .C(n7502) );
  CKBD0 U7419 ( .CLK(n7471), .C(n7503) );
  CKBD0 U7420 ( .CLK(n7472), .C(n7504) );
  CKBD0 U7421 ( .CLK(n7473), .C(n7505) );
  CKBD0 U7422 ( .CLK(n7474), .C(n7506) );
  CKBD0 U7423 ( .CLK(n7475), .C(n7507) );
  CKBD0 U7424 ( .CLK(n7476), .C(n7508) );
  CKBD0 U7425 ( .CLK(n7477), .C(n7509) );
  CKBD0 U7426 ( .CLK(n7478), .C(n7510) );
  CKBD0 U7427 ( .CLK(n7479), .C(n7511) );
  CKBD0 U7428 ( .CLK(n7480), .C(n7512) );
  CKBD0 U7429 ( .CLK(n7482), .C(n7513) );
  CKBD0 U7430 ( .CLK(n7481), .C(n7514) );
  CKBD0 U7431 ( .CLK(n7483), .C(n7515) );
  CKBD0 U7432 ( .CLK(n7484), .C(n7516) );
  CKBD0 U7433 ( .CLK(n7485), .C(n7517) );
  CKBD0 U7434 ( .CLK(n7486), .C(n7518) );
  CKBD0 U7435 ( .CLK(n7487), .C(n7519) );
  CKBD0 U7436 ( .CLK(n7488), .C(n7520) );
  CKBD0 U7437 ( .CLK(n7489), .C(n7521) );
  BUFFD0 U7438 ( .I(n7490), .Z(n7522) );
  CKBD0 U7439 ( .CLK(n7491), .C(n7523) );
  CKBD0 U7440 ( .CLK(n7492), .C(n7524) );
  CKBD0 U7441 ( .CLK(n7493), .C(n7525) );
  CKBD0 U7442 ( .CLK(n7494), .C(n7526) );
  CKBD0 U7443 ( .CLK(n7495), .C(n7527) );
  CKBD0 U7444 ( .CLK(n7496), .C(n7528) );
  CKBD0 U7445 ( .CLK(n7497), .C(n7529) );
  CKBD0 U7446 ( .CLK(n7498), .C(n7530) );
  CKBD0 U7447 ( .CLK(n7499), .C(n7531) );
  CKBD0 U7448 ( .CLK(n7500), .C(n7532) );
  CKBD0 U7449 ( .CLK(n7501), .C(n7533) );
  CKBD0 U7450 ( .CLK(n7502), .C(n7534) );
  CKBD0 U7451 ( .CLK(n7503), .C(n7535) );
  CKBD0 U7452 ( .CLK(n7504), .C(n7536) );
  CKBD0 U7453 ( .CLK(n7505), .C(n7537) );
  CKBD0 U7454 ( .CLK(n7506), .C(n7538) );
  CKBD0 U7455 ( .CLK(n7508), .C(n7539) );
  CKBD0 U7456 ( .CLK(n7509), .C(n7540) );
  CKBD0 U7457 ( .CLK(n7507), .C(n7541) );
  CKBD0 U7458 ( .CLK(n7510), .C(n7542) );
  CKBD0 U7459 ( .CLK(n7511), .C(n7543) );
  CKBD0 U7460 ( .CLK(n7512), .C(n7544) );
  CKBD0 U7461 ( .CLK(n7513), .C(n7545) );
  CKBD0 U7462 ( .CLK(n7514), .C(n7546) );
  CKBD0 U7463 ( .CLK(n7515), .C(n7547) );
  CKBD0 U7464 ( .CLK(n7516), .C(n7548) );
  CKBD0 U7465 ( .CLK(n7517), .C(n7549) );
  CKBD0 U7466 ( .CLK(n7518), .C(n7550) );
  CKBD0 U7467 ( .CLK(n7519), .C(n7551) );
  CKBD0 U7468 ( .CLK(n7520), .C(n7552) );
  CKBD0 U7469 ( .CLK(n7521), .C(n7553) );
  CKBD0 U7470 ( .CLK(n7522), .C(n7554) );
  CKBD0 U7471 ( .CLK(n7523), .C(n7555) );
  CKBD0 U7472 ( .CLK(n7524), .C(n7556) );
  CKBD0 U7473 ( .CLK(n7525), .C(n7557) );
  BUFFD0 U7474 ( .I(n7527), .Z(n7558) );
  CKBD0 U7475 ( .CLK(n7526), .C(n7559) );
  BUFFD0 U7476 ( .I(n7530), .Z(n7560) );
  CKBD0 U7477 ( .CLK(n7528), .C(n7561) );
  CKBD0 U7478 ( .CLK(n7529), .C(n7562) );
  BUFFD0 U7479 ( .I(n7531), .Z(n7563) );
  BUFFD0 U7480 ( .I(n7532), .Z(n7564) );
  CKBD0 U7481 ( .CLK(n7533), .C(n7565) );
  BUFFD0 U7482 ( .I(n7534), .Z(n7566) );
  CKBD0 U7483 ( .CLK(n7535), .C(n7567) );
  CKBD0 U7484 ( .CLK(n7536), .C(n7568) );
  CKBD0 U7485 ( .CLK(n7537), .C(n7569) );
  CKBD0 U7486 ( .CLK(n7538), .C(n7570) );
  BUFFD0 U7487 ( .I(n7539), .Z(n7571) );
  CKBD0 U7488 ( .CLK(n7541), .C(n7572) );
  CKBD0 U7489 ( .CLK(n7540), .C(n7573) );
  CKBD0 U7490 ( .CLK(n7542), .C(n7574) );
  CKBD0 U7491 ( .CLK(n7543), .C(n7575) );
  BUFFD0 U7492 ( .I(n7544), .Z(n7576) );
  CKBD0 U7493 ( .CLK(n7545), .C(n7577) );
  CKBD0 U7494 ( .CLK(n7547), .C(n7578) );
  CKBD0 U7495 ( .CLK(n7546), .C(n7579) );
  CKBD0 U7496 ( .CLK(n7548), .C(n7580) );
  CKBD0 U7497 ( .CLK(n7549), .C(n7581) );
  CKBD0 U7498 ( .CLK(n7550), .C(n7582) );
  CKBD0 U7499 ( .CLK(n7551), .C(n7583) );
  CKBD0 U7500 ( .CLK(n7552), .C(n7584) );
  CKBD0 U7501 ( .CLK(n7553), .C(n7585) );
  CKBD0 U7502 ( .CLK(n7554), .C(n7586) );
  CKBD0 U7503 ( .CLK(n7555), .C(n7587) );
  CKBD0 U7504 ( .CLK(n7556), .C(n7588) );
  CKBD0 U7505 ( .CLK(n7557), .C(n7589) );
  CKBD0 U7506 ( .CLK(n7558), .C(n7590) );
  CKBD0 U7507 ( .CLK(n7559), .C(n7591) );
  CKBD0 U7508 ( .CLK(n7560), .C(n7592) );
  CKBD0 U7509 ( .CLK(n7561), .C(n7593) );
  CKBD0 U7510 ( .CLK(n7562), .C(n7594) );
  CKBD0 U7511 ( .CLK(n7563), .C(n7595) );
  CKBD0 U7512 ( .CLK(n7564), .C(n7596) );
  CKBD0 U7513 ( .CLK(n7565), .C(n7597) );
  CKBD0 U7514 ( .CLK(n7566), .C(n7598) );
  CKBD0 U7515 ( .CLK(n7567), .C(n7599) );
  CKBD0 U7516 ( .CLK(n7568), .C(n7600) );
  CKBD0 U7517 ( .CLK(n7569), .C(n7601) );
  CKBD0 U7518 ( .CLK(n7570), .C(n7602) );
  BUFFD0 U7519 ( .I(n7572), .Z(n7603) );
  CKBD0 U7520 ( .CLK(n7571), .C(n7604) );
  CKBD0 U7521 ( .CLK(n7573), .C(n7605) );
  CKBD0 U7522 ( .CLK(n7574), .C(n7606) );
  CKBD0 U7523 ( .CLK(n7575), .C(n7607) );
  CKBD0 U7524 ( .CLK(n7576), .C(n7608) );
  CKBD0 U7525 ( .CLK(n7577), .C(n7609) );
  CKBD0 U7526 ( .CLK(n7581), .C(n7610) );
  CKBD0 U7527 ( .CLK(n7578), .C(n7611) );
  CKBD0 U7528 ( .CLK(n7580), .C(n7612) );
  CKBD0 U7529 ( .CLK(n7579), .C(n7613) );
  CKBD0 U7530 ( .CLK(n7582), .C(n7614) );
  CKBD0 U7531 ( .CLK(n7583), .C(n7615) );
  CKBD0 U7532 ( .CLK(n7584), .C(n7616) );
  CKBD0 U7533 ( .CLK(n7585), .C(n7617) );
  CKBD0 U7534 ( .CLK(n7586), .C(n7618) );
  CKBD0 U7535 ( .CLK(n7587), .C(n7619) );
  CKBD0 U7536 ( .CLK(n7589), .C(n7620) );
  CKBD0 U7537 ( .CLK(n7588), .C(n7621) );
  CKBD0 U7538 ( .CLK(n7590), .C(n7622) );
  CKBD0 U7539 ( .CLK(n7591), .C(n7623) );
  CKBD0 U7540 ( .CLK(n7592), .C(n7624) );
  CKBD0 U7541 ( .CLK(n7593), .C(n7625) );
  CKBD0 U7542 ( .CLK(n7594), .C(n7626) );
  CKBD0 U7543 ( .CLK(n7595), .C(n7627) );
  CKBD0 U7544 ( .CLK(n7596), .C(n7628) );
  CKBD0 U7545 ( .CLK(n7597), .C(n7629) );
  CKBD0 U7546 ( .CLK(n7598), .C(n7630) );
  BUFFD0 U7547 ( .I(n7599), .Z(n7631) );
  CKBD0 U7548 ( .CLK(n7600), .C(n7632) );
  BUFFD0 U7549 ( .I(n7601), .Z(n7633) );
  BUFFD0 U7550 ( .I(n7602), .Z(n7634) );
  CKBD0 U7551 ( .CLK(n7604), .C(n7635) );
  CKBD0 U7552 ( .CLK(n7606), .C(n7636) );
  CKBD0 U7553 ( .CLK(n7605), .C(n7637) );
  CKBD0 U7554 ( .CLK(n7607), .C(n7638) );
  CKBD0 U7555 ( .CLK(n7608), .C(n7639) );
  CKBD0 U7556 ( .CLK(n7609), .C(n7640) );
  BUFFD0 U7557 ( .I(n7610), .Z(n7641) );
  CKBD0 U7558 ( .CLK(n7611), .C(n7642) );
  CKBD0 U7559 ( .CLK(n7612), .C(n7643) );
  CKBD0 U7560 ( .CLK(n7614), .C(n7644) );
  CKBD0 U7561 ( .CLK(n7616), .C(n7645) );
  CKBD0 U7562 ( .CLK(n7615), .C(n7646) );
  CKBD0 U7563 ( .CLK(n7617), .C(n7647) );
  CKBD0 U7564 ( .CLK(n7618), .C(n7648) );
  CKBD0 U7565 ( .CLK(n7619), .C(n7649) );
  BUFFD0 U7566 ( .I(n7620), .Z(n7650) );
  CKBD0 U7567 ( .CLK(n7621), .C(n7651) );
  CKBD0 U7568 ( .CLK(n7622), .C(n7652) );
  CKBD0 U7569 ( .CLK(n7623), .C(n7653) );
  CKBD0 U7570 ( .CLK(n7625), .C(n7654) );
  CKBD0 U7571 ( .CLK(n7626), .C(n7655) );
  CKBD0 U7572 ( .CLK(n7632), .C(n7656) );
  CKBD0 U7573 ( .CLK(n7633), .C(n7657) );
  CKBD0 U7574 ( .CLK(n7634), .C(n7658) );
  CKBD0 U7575 ( .CLK(n7637), .C(n7659) );
  CKBD0 U7576 ( .CLK(n7635), .C(n7660) );
  BUFFD0 U7577 ( .I(n7636), .Z(n7661) );
  CKBD0 U7578 ( .CLK(n7638), .C(n7662) );
  CKBD0 U7579 ( .CLK(n7639), .C(n7663) );
  CKBD0 U7580 ( .CLK(n7603), .C(n7664) );
  CKBD0 U7581 ( .CLK(n7613), .C(n7665) );
  CKBD0 U7582 ( .CLK(n7624), .C(n7666) );
  CKBD0 U7583 ( .CLK(n7627), .C(n7667) );
  CKBD0 U7584 ( .CLK(n7628), .C(n7668) );
  BUFFD0 U7585 ( .I(n7629), .Z(n7669) );
  CKBD0 U7586 ( .CLK(n7630), .C(n7670) );
  CKBD0 U7587 ( .CLK(n7640), .C(n7671) );
  CKBD0 U7588 ( .CLK(n7641), .C(n7672) );
  CKBD0 U7589 ( .CLK(n7642), .C(n7673) );
  CKBD0 U7590 ( .CLK(n7643), .C(n7674) );
  CKBD0 U7591 ( .CLK(n7631), .C(n7675) );
  CKBD0 U7592 ( .CLK(n7644), .C(n7676) );
  CKBD0 U7593 ( .CLK(n7664), .C(n7677) );
  BUFFD0 U7594 ( .I(n7665), .Z(n7678) );
  CKBD0 U7595 ( .CLK(n7666), .C(n7679) );
  CKBD0 U7596 ( .CLK(n7667), .C(n7680) );
  CKBD0 U7597 ( .CLK(n7668), .C(n7681) );
  CKBD0 U7598 ( .CLK(n7669), .C(n7682) );
  CKBD0 U7599 ( .CLK(n7670), .C(n7683) );
  BUFFD0 U7600 ( .I(n7645), .Z(n7684) );
  CKBD0 U7601 ( .CLK(n7646), .C(n7685) );
  CKBD0 U7602 ( .CLK(n7647), .C(n7686) );
  CKBD0 U7603 ( .CLK(n7648), .C(n7687) );
  CKBD0 U7604 ( .CLK(n7675), .C(n7688) );
  CKBD0 U7605 ( .CLK(n7649), .C(n7689) );
  CKBD0 U7606 ( .CLK(n7650), .C(n7690) );
  CKBD0 U7607 ( .CLK(n7651), .C(n7691) );
  CKBD0 U7608 ( .CLK(n7652), .C(n7692) );
  CKBD0 U7609 ( .CLK(n7653), .C(n7693) );
  CKBD0 U7610 ( .CLK(n7677), .C(n7694) );
  CKBD0 U7611 ( .CLK(n7654), .C(n7695) );
  CKBD0 U7612 ( .CLK(n7655), .C(n7696) );
  CKBD0 U7613 ( .CLK(n7678), .C(n7697) );
  CKBD0 U7614 ( .CLK(n7679), .C(n7698) );
  BUFFD0 U7615 ( .I(n7656), .Z(n7699) );
  CKBD0 U7616 ( .CLK(n7657), .C(n7700) );
  CKBD0 U7617 ( .CLK(n7658), .C(n7701) );
  CKBD0 U7618 ( .CLK(n7680), .C(n7702) );
  CKBD0 U7619 ( .CLK(n7681), .C(n7703) );
  CKBD0 U7620 ( .CLK(n7682), .C(n7704) );
  CKBD0 U7621 ( .CLK(n7683), .C(n7705) );
  CKBD0 U7622 ( .CLK(n7688), .C(n7706) );
  CKBD0 U7623 ( .CLK(n7694), .C(n7707) );
  CKBD0 U7624 ( .CLK(n7697), .C(n7708) );
  CKBD0 U7625 ( .CLK(n7698), .C(n7709) );
  CKBD0 U7626 ( .CLK(n7660), .C(n7710) );
  BUFFD0 U7627 ( .I(n7659), .Z(n7711) );
  CKBD0 U7628 ( .CLK(n7662), .C(n7712) );
  CKBD0 U7629 ( .CLK(n7661), .C(n7713) );
  CKBD0 U7630 ( .CLK(n7663), .C(n7714) );
  CKBD0 U7631 ( .CLK(n7702), .C(n7715) );
  CKBD0 U7632 ( .CLK(n7703), .C(n7716) );
  CKBD0 U7633 ( .CLK(n7704), .C(n7717) );
  CKBD0 U7634 ( .CLK(n7705), .C(n7718) );
  CKBD0 U7635 ( .CLK(n7706), .C(n7719) );
  CKBD0 U7636 ( .CLK(n7707), .C(n7720) );
  CKBD0 U7637 ( .CLK(n7708), .C(n7721) );
  CKBD0 U7638 ( .CLK(n7709), .C(n7722) );
  BUFFD0 U7639 ( .I(n7671), .Z(n7723) );
  CKBD0 U7640 ( .CLK(n7674), .C(n7724) );
  CKBD0 U7641 ( .CLK(n7672), .C(n7725) );
  CKBD0 U7642 ( .CLK(n7673), .C(n7726) );
  CKBD0 U7643 ( .CLK(n7715), .C(n7727) );
  BUFFD0 U7644 ( .I(n7676), .Z(n7728) );
  CKBD0 U7645 ( .CLK(n7716), .C(n7729) );
  CKBD0 U7646 ( .CLK(n7717), .C(n7730) );
  CKBD0 U7647 ( .CLK(n7718), .C(n7731) );
  CKBD0 U7648 ( .CLK(n7719), .C(n7732) );
  CKBD0 U7649 ( .CLK(n7720), .C(n7733) );
  CKBD0 U7650 ( .CLK(n7721), .C(n7734) );
  CKBD0 U7651 ( .CLK(n7722), .C(n7735) );
  CKBD0 U7652 ( .CLK(n7684), .C(n7736) );
  CKBD0 U7653 ( .CLK(n7685), .C(n7737) );
  CKBD0 U7654 ( .CLK(n7686), .C(n7738) );
  CKBD0 U7655 ( .CLK(n7687), .C(n7739) );
  CKBD0 U7656 ( .CLK(n7727), .C(n7740) );
  CKBD0 U7657 ( .CLK(n7729), .C(n7741) );
  CKBD0 U7658 ( .CLK(n7730), .C(n7742) );
  CKBD0 U7659 ( .CLK(n7731), .C(n7743) );
  CKBD0 U7660 ( .CLK(n7732), .C(n7744) );
  CKBD0 U7661 ( .CLK(n7733), .C(n7745) );
  CKBD0 U7662 ( .CLK(n7734), .C(n7746) );
  CKBD0 U7663 ( .CLK(n7735), .C(n7747) );
  CKBD0 U7664 ( .CLK(n7689), .C(n7748) );
  CKBD0 U7665 ( .CLK(n7690), .C(n7749) );
  CKBD0 U7666 ( .CLK(n7691), .C(n7750) );
  CKBD0 U7667 ( .CLK(n7692), .C(n7751) );
  CKBD0 U7668 ( .CLK(n7740), .C(n7752) );
  CKBD0 U7669 ( .CLK(n7741), .C(n7753) );
  CKBD0 U7670 ( .CLK(n7742), .C(n7754) );
  CKBD0 U7671 ( .CLK(n7743), .C(n7755) );
  CKBD0 U7672 ( .CLK(n7744), .C(n7756) );
  CKBD0 U7673 ( .CLK(n7745), .C(n7757) );
  CKBD0 U7674 ( .CLK(n7746), .C(n7758) );
  CKBD0 U7675 ( .CLK(n7747), .C(n7759) );
  BUFFD0 U7676 ( .I(n7695), .Z(n7760) );
  CKBD0 U7677 ( .CLK(n7693), .C(n7761) );
  CKBD0 U7678 ( .CLK(n7752), .C(n7762) );
  CKBD0 U7679 ( .CLK(n7753), .C(n7763) );
  CKBD0 U7680 ( .CLK(n7696), .C(n7764) );
  CKBD0 U7681 ( .CLK(n7754), .C(n7765) );
  CKBD0 U7682 ( .CLK(n7755), .C(n7766) );
  CKBD0 U7683 ( .CLK(n7756), .C(n7767) );
  CKBD0 U7684 ( .CLK(n7699), .C(n7768) );
  CKBD0 U7685 ( .CLK(n7757), .C(n7769) );
  CKBD0 U7686 ( .CLK(n7700), .C(n7770) );
  CKBD0 U7687 ( .CLK(n7701), .C(n7771) );
  CKBD0 U7688 ( .CLK(n7758), .C(n7772) );
  CKBD0 U7689 ( .CLK(n7710), .C(n7773) );
  CKBD0 U7690 ( .CLK(n7711), .C(n7774) );
  CKBD0 U7691 ( .CLK(n7713), .C(n7775) );
  BUFFD0 U7692 ( .I(n7712), .Z(n7776) );
  CKBD0 U7693 ( .CLK(n7714), .C(n7777) );
  CKBD0 U7694 ( .CLK(n7723), .C(n7778) );
  CKBD0 U7695 ( .CLK(n7759), .C(n7779) );
  CKBD0 U7696 ( .CLK(n7762), .C(n7780) );
  CKBD0 U7697 ( .CLK(n7763), .C(n7781) );
  CKBD0 U7698 ( .CLK(n7765), .C(n7782) );
  CKBD0 U7699 ( .CLK(n7766), .C(n7783) );
  CKBD0 U7700 ( .CLK(n7767), .C(n7784) );
  BUFFD0 U7701 ( .I(n7769), .Z(n7785) );
  CKBD0 U7702 ( .CLK(n7772), .C(n7786) );
  BUFFD0 U7703 ( .I(n7724), .Z(n7787) );
  CKBD0 U7704 ( .CLK(n7725), .C(n7788) );
  CKBD0 U7705 ( .CLK(n7726), .C(n7789) );
  BUFFD0 U7706 ( .I(n7779), .Z(n7790) );
  BUFFD0 U7707 ( .I(n7780), .Z(n7791) );
  BUFFD0 U7708 ( .I(n7781), .Z(n7792) );
  CKBD0 U7709 ( .CLK(n7782), .C(n7793) );
  CKBD0 U7710 ( .CLK(n7783), .C(n7794) );
  CKBD0 U7711 ( .CLK(n7784), .C(n7795) );
  CKBD0 U7712 ( .CLK(n7785), .C(n7796) );
  CKBD0 U7713 ( .CLK(n7728), .C(n7797) );
  CKBD0 U7714 ( .CLK(n7786), .C(n7798) );
  CKBD0 U7715 ( .CLK(n7736), .C(n7799) );
  CKBD0 U7716 ( .CLK(n7737), .C(n7800) );
  CKBD0 U7717 ( .CLK(n7790), .C(n7801) );
  CKBD0 U7718 ( .CLK(n7791), .C(n7802) );
  CKBD0 U7719 ( .CLK(n7792), .C(n7803) );
  BUFFD0 U7720 ( .I(n7793), .Z(n7804) );
  BUFFD0 U7721 ( .I(n7794), .Z(n7805) );
  CKBD0 U7722 ( .CLK(n7795), .C(n7806) );
  CKBD0 U7723 ( .CLK(n7796), .C(n7807) );
  BUFFD0 U7724 ( .I(n7798), .Z(n7808) );
  CKBD0 U7725 ( .CLK(n7801), .C(n7809) );
  CKBD0 U7726 ( .CLK(n7802), .C(n7810) );
  CKBD0 U7727 ( .CLK(n7803), .C(n7811) );
  CKBD0 U7728 ( .CLK(n7804), .C(n7812) );
  CKBD0 U7729 ( .CLK(n7805), .C(n7813) );
  BUFFD0 U7730 ( .I(n7806), .Z(n7814) );
  CKBD0 U7731 ( .CLK(n7807), .C(n7815) );
  CKBD0 U7732 ( .CLK(n7738), .C(n7816) );
  CKBD0 U7733 ( .CLK(n7739), .C(n7817) );
  CKBD0 U7734 ( .CLK(n7748), .C(n7818) );
  CKBD0 U7735 ( .CLK(n7749), .C(n7819) );
  CKBD0 U7736 ( .CLK(n7808), .C(n7820) );
  CKBD0 U7737 ( .CLK(n7750), .C(n7821) );
  CKBD0 U7738 ( .CLK(n7809), .C(n7822) );
  CKBD0 U7739 ( .CLK(n7810), .C(n7823) );
  CKBD0 U7740 ( .CLK(n7811), .C(n7824) );
  CKBD0 U7741 ( .CLK(n7812), .C(n7825) );
  CKBD0 U7742 ( .CLK(n7813), .C(n7826) );
  CKBD0 U7743 ( .CLK(n7814), .C(n7827) );
  CKBD0 U7744 ( .CLK(n7815), .C(n7828) );
  CKBD0 U7745 ( .CLK(n7751), .C(n7829) );
  CKBD0 U7746 ( .CLK(n7820), .C(n7830) );
  CKBD0 U7747 ( .CLK(n7760), .C(n7831) );
  CKBD0 U7748 ( .CLK(n7822), .C(n7832) );
  CKBD0 U7749 ( .CLK(n7823), .C(n7833) );
  CKBD0 U7750 ( .CLK(n7824), .C(n7834) );
  CKBD0 U7751 ( .CLK(n7825), .C(n7835) );
  CKBD0 U7752 ( .CLK(n7826), .C(n7836) );
  CKBD0 U7753 ( .CLK(n7827), .C(n7837) );
  CKBD0 U7754 ( .CLK(n7828), .C(n7838) );
  CKBD0 U7755 ( .CLK(n7761), .C(n7839) );
  CKBD0 U7756 ( .CLK(n7830), .C(n7840) );
  CKBD0 U7757 ( .CLK(n7832), .C(n7841) );
  CKBD0 U7758 ( .CLK(n7833), .C(n7842) );
  CKBD0 U7759 ( .CLK(n7834), .C(n7843) );
  CKBD0 U7760 ( .CLK(n7835), .C(n7844) );
  CKBD0 U7761 ( .CLK(n7836), .C(n7845) );
  CKBD0 U7762 ( .CLK(n7837), .C(n7846) );
  CKBD0 U7763 ( .CLK(n7838), .C(n7847) );
  CKBD0 U7764 ( .CLK(n7764), .C(n7848) );
  CKBD0 U7765 ( .CLK(n7840), .C(n7849) );
  CKBD0 U7766 ( .CLK(n7768), .C(n7850) );
  CKBD0 U7767 ( .CLK(n7841), .C(n7851) );
  CKBD0 U7768 ( .CLK(n7770), .C(n7852) );
  CKBD0 U7769 ( .CLK(n7771), .C(n7853) );
  CKBD0 U7770 ( .CLK(n7773), .C(n7854) );
  CKBD0 U7771 ( .CLK(n7774), .C(n7855) );
  CKBD0 U7772 ( .CLK(n7842), .C(n7856) );
  CKBD0 U7773 ( .CLK(n7843), .C(n7857) );
  CKBD0 U7774 ( .CLK(n7775), .C(n7858) );
  CKBD0 U7775 ( .CLK(n7776), .C(n7859) );
  CKBD0 U7776 ( .CLK(n7777), .C(n7860) );
  CKBD0 U7777 ( .CLK(n7844), .C(n7861) );
  CKBD0 U7778 ( .CLK(n7845), .C(n7862) );
  CKBD0 U7779 ( .CLK(n7846), .C(n7863) );
  CKBD0 U7780 ( .CLK(n7847), .C(n7864) );
  CKBD0 U7781 ( .CLK(n7849), .C(n7865) );
  CKBD0 U7782 ( .CLK(n7851), .C(n7866) );
  CKBD0 U7783 ( .CLK(n7778), .C(n7867) );
  CKBD0 U7784 ( .CLK(n7787), .C(n7868) );
  CKBD0 U7785 ( .CLK(n7788), .C(n7869) );
  CKBD0 U7786 ( .CLK(n7856), .C(n7870) );
  CKBD0 U7787 ( .CLK(n7789), .C(n7871) );
  CKBD0 U7788 ( .CLK(n7857), .C(n7872) );
  CKBD0 U7789 ( .CLK(n7861), .C(n7873) );
  CKBD0 U7790 ( .CLK(n7862), .C(n7874) );
  CKBD0 U7791 ( .CLK(n7863), .C(n7875) );
  CKBD0 U7792 ( .CLK(n7864), .C(n7876) );
  CKBD0 U7793 ( .CLK(n7865), .C(n7877) );
  CKBD0 U7794 ( .CLK(n7866), .C(n7878) );
  CKBD0 U7795 ( .CLK(n7797), .C(n7879) );
  CKBD0 U7796 ( .CLK(n7800), .C(n7880) );
  CKBD0 U7797 ( .CLK(n7799), .C(n7881) );
  CKBD0 U7798 ( .CLK(n7816), .C(n7882) );
  CKBD0 U7799 ( .CLK(n7870), .C(n7883) );
  CKBD0 U7800 ( .CLK(n7872), .C(n7884) );
  CKBD0 U7801 ( .CLK(n7817), .C(n7885) );
  CKBD0 U7802 ( .CLK(n7873), .C(n7886) );
  CKBD0 U7803 ( .CLK(n7874), .C(n7887) );
  CKBD0 U7804 ( .CLK(n7875), .C(n7888) );
  CKBD0 U7805 ( .CLK(n7876), .C(n7889) );
  CKBD0 U7806 ( .CLK(n7877), .C(n7890) );
  CKBD0 U7807 ( .CLK(n7878), .C(n7891) );
  CKBD0 U7808 ( .CLK(n7818), .C(n7892) );
  CKBD0 U7809 ( .CLK(n7821), .C(n7893) );
  CKBD0 U7810 ( .CLK(n7819), .C(n7894) );
  CKBD0 U7811 ( .CLK(n7883), .C(n7895) );
  CKBD0 U7812 ( .CLK(n7884), .C(n7896) );
  BUFFD0 U7813 ( .I(n7839), .Z(n7897) );
  CKBD0 U7814 ( .CLK(n7886), .C(n7898) );
  CKBD0 U7815 ( .CLK(n7887), .C(n7899) );
  CKBD0 U7816 ( .CLK(n7888), .C(n7900) );
  CKBD0 U7817 ( .CLK(n7889), .C(n7901) );
  CKBD0 U7818 ( .CLK(n7890), .C(n7902) );
  CKBD0 U7819 ( .CLK(n7891), .C(n7903) );
  CKBD0 U7820 ( .CLK(n7829), .C(n7904) );
  CKBD0 U7821 ( .CLK(n7895), .C(n7905) );
  CKBD0 U7822 ( .CLK(n7896), .C(n7906) );
  CKBD0 U7823 ( .CLK(n7898), .C(n7907) );
  CKBD0 U7824 ( .CLK(n7899), .C(n7908) );
  CKBD0 U7825 ( .CLK(n7900), .C(n7909) );
  BUFFD0 U7826 ( .I(n7901), .Z(n7910) );
  CKBD0 U7827 ( .CLK(n7902), .C(n7911) );
  CKBD0 U7828 ( .CLK(n7903), .C(n7912) );
  CKBD0 U7829 ( .CLK(n7831), .C(n7913) );
  BUFFD0 U7830 ( .I(n7905), .Z(n7914) );
  BUFFD0 U7831 ( .I(n7906), .Z(n7915) );
  CKBD0 U7832 ( .CLK(n7848), .C(n7916) );
  CKBD0 U7833 ( .CLK(n7907), .C(n7917) );
  BUFFD0 U7834 ( .I(n7908), .Z(n7918) );
  CKBD0 U7835 ( .CLK(n7909), .C(n7919) );
  CKBD0 U7836 ( .CLK(n7910), .C(n7920) );
  CKBD0 U7837 ( .CLK(n7850), .C(n7921) );
  CKBD0 U7838 ( .CLK(n7852), .C(n7922) );
  CKBD0 U7839 ( .CLK(n7853), .C(n7923) );
  CKBD0 U7840 ( .CLK(n7911), .C(n7924) );
  BUFFD0 U7841 ( .I(n7912), .Z(n7925) );
  CKBD0 U7842 ( .CLK(n7914), .C(n7926) );
  CKBD0 U7843 ( .CLK(n7915), .C(n7927) );
  CKBD0 U7844 ( .CLK(n7917), .C(n7928) );
  CKBD0 U7845 ( .CLK(n7918), .C(n7929) );
  BUFFD0 U7846 ( .I(n7919), .Z(n7930) );
  CKBD0 U7847 ( .CLK(n7920), .C(n7931) );
  BUFFD0 U7848 ( .I(n7854), .Z(n7932) );
  CKBD0 U7849 ( .CLK(n7855), .C(n7933) );
  CKBD0 U7850 ( .CLK(n7858), .C(n7934) );
  CKBD0 U7851 ( .CLK(n7859), .C(n7935) );
  BUFFD0 U7852 ( .I(n7860), .Z(n7936) );
  CKBD0 U7853 ( .CLK(n7924), .C(n7937) );
  CKBD0 U7854 ( .CLK(n7925), .C(n7938) );
  CKBD0 U7855 ( .CLK(n7926), .C(n7939) );
  CKBD0 U7856 ( .CLK(n7927), .C(n7940) );
  BUFFD0 U7857 ( .I(n7928), .Z(n7941) );
  CKBD0 U7858 ( .CLK(n7929), .C(n7942) );
  CKBD0 U7859 ( .CLK(n7930), .C(n7943) );
  CKBD0 U7860 ( .CLK(n7931), .C(n7944) );
  CKBD0 U7861 ( .CLK(n7867), .C(n7945) );
  CKBD0 U7862 ( .CLK(n7869), .C(n7946) );
  CKBD0 U7863 ( .CLK(n7871), .C(n7947) );
  CKBD0 U7864 ( .CLK(n7868), .C(n7948) );
  CKBD0 U7865 ( .CLK(n7879), .C(n7949) );
  BUFFD0 U7866 ( .I(n7937), .Z(n7950) );
  CKBD0 U7867 ( .CLK(n7938), .C(n7951) );
  CKBD0 U7868 ( .CLK(n7939), .C(n7952) );
  CKBD0 U7869 ( .CLK(n7940), .C(n7953) );
  CKBD0 U7870 ( .CLK(n7941), .C(n7954) );
  CKBD0 U7871 ( .CLK(n7942), .C(n7955) );
  CKBD0 U7872 ( .CLK(n7943), .C(n7956) );
  CKBD0 U7873 ( .CLK(n7944), .C(n7957) );
  CKBD0 U7874 ( .CLK(n7881), .C(n7958) );
  BUFFD0 U7875 ( .I(n7880), .Z(n7959) );
  CKBD0 U7876 ( .CLK(n7882), .C(n7960) );
  CKBD0 U7877 ( .CLK(n7885), .C(n7961) );
  BUFFD0 U7878 ( .I(n7892), .Z(n7962) );
  CKBD0 U7879 ( .CLK(n7950), .C(n7963) );
  CKBD0 U7880 ( .CLK(n7894), .C(n7964) );
  CKBD0 U7881 ( .CLK(n7951), .C(n7965) );
  CKBD0 U7882 ( .CLK(n7952), .C(n7966) );
  CKBD0 U7883 ( .CLK(n7953), .C(n7967) );
  CKBD0 U7884 ( .CLK(n7954), .C(n7968) );
  CKBD0 U7885 ( .CLK(n7955), .C(n7969) );
  CKBD0 U7886 ( .CLK(n7956), .C(n7970) );
  CKBD0 U7887 ( .CLK(n7957), .C(n7971) );
  BUFFD0 U7888 ( .I(n7893), .Z(n7972) );
  CKBD0 U7889 ( .CLK(n7897), .C(n7973) );
  CKBD0 U7890 ( .CLK(n7904), .C(n7974) );
  CKBD0 U7891 ( .CLK(n7963), .C(n7975) );
  CKBD0 U7892 ( .CLK(n7965), .C(n7976) );
  CKBD0 U7893 ( .CLK(n7966), .C(n7977) );
  CKBD0 U7894 ( .CLK(n7967), .C(n7978) );
  CKBD0 U7895 ( .CLK(n7968), .C(n7979) );
  CKBD0 U7896 ( .CLK(n7969), .C(n7980) );
  CKBD0 U7897 ( .CLK(n7970), .C(n7981) );
  CKBD0 U7898 ( .CLK(n7971), .C(n7982) );
  CKBD0 U7899 ( .CLK(n7913), .C(n7983) );
  BUFFD0 U7900 ( .I(n7916), .Z(n7984) );
  CKBD0 U7901 ( .CLK(n7975), .C(n7985) );
  CKBD0 U7902 ( .CLK(n7976), .C(n7986) );
  CKBD0 U7903 ( .CLK(n7921), .C(n7987) );
  CKBD0 U7904 ( .CLK(n7977), .C(n7988) );
  CKBD0 U7905 ( .CLK(n7978), .C(n7989) );
  BUFFD0 U7906 ( .I(n7922), .Z(n7990) );
  BUFFD0 U7907 ( .I(n7923), .Z(n7991) );
  CKBD0 U7908 ( .CLK(n7979), .C(n7992) );
  CKBD0 U7909 ( .CLK(n7932), .C(n7993) );
  CKBD0 U7910 ( .CLK(n7933), .C(n7994) );
  CKBD0 U7911 ( .CLK(n7934), .C(n7995) );
  CKBD0 U7912 ( .CLK(n7936), .C(n7996) );
  CKBD0 U7913 ( .CLK(n7935), .C(n7997) );
  CKBD0 U7914 ( .CLK(n7945), .C(n7998) );
  CKBD0 U7915 ( .CLK(n7980), .C(n7999) );
  BUFFD0 U7916 ( .I(n7946), .Z(n8000) );
  BUFFD0 U7917 ( .I(n7947), .Z(n8001) );
  CKBD0 U7918 ( .CLK(n7948), .C(n8002) );
  CKBD0 U7919 ( .CLK(n7949), .C(n8003) );
  BUFFD0 U7920 ( .I(n7958), .Z(n8004) );
  CKBD0 U7921 ( .CLK(n7981), .C(n8005) );
  CKBD0 U7922 ( .CLK(n7959), .C(n8006) );
  BUFFD0 U7923 ( .I(n7960), .Z(n8007) );
  BUFFD0 U7924 ( .I(n7961), .Z(n8008) );
  BUFFD0 U7925 ( .I(n8885), .Z(n8009) );
  CKBD0 U7926 ( .CLK(n7962), .C(n8010) );
  BUFFD0 U7927 ( .I(n7974), .Z(n8011) );
  CKBD0 U7928 ( .CLK(n7972), .C(n8012) );
  CKBD0 U7929 ( .CLK(n7973), .C(n8013) );
  CKBD0 U7930 ( .CLK(n7982), .C(n8014) );
  CKBD0 U7931 ( .CLK(n7983), .C(n8015) );
  CKBD0 U7932 ( .CLK(n7984), .C(n8016) );
  CKBD0 U7933 ( .CLK(n7985), .C(n8017) );
  CKBD0 U7934 ( .CLK(n7986), .C(n8018) );
  CKBD0 U7935 ( .CLK(n7988), .C(n8019) );
  CKBD0 U7936 ( .CLK(n7989), .C(n8020) );
  CKBD0 U7937 ( .CLK(n7992), .C(n8021) );
  CKBD0 U7938 ( .CLK(n7999), .C(n8022) );
  CKBD0 U7939 ( .CLK(n8005), .C(n8023) );
  CKBD0 U7940 ( .CLK(n8014), .C(n8024) );
  CKBD0 U7941 ( .CLK(n8017), .C(n8025) );
  BUFFD0 U7942 ( .I(n7987), .Z(n8026) );
  CKBD0 U7943 ( .CLK(n8018), .C(n8027) );
  CKBD0 U7944 ( .CLK(n7990), .C(n8028) );
  CKBD0 U7945 ( .CLK(n7991), .C(n8029) );
  CKBD0 U7946 ( .CLK(n8019), .C(n8030) );
  CKBD0 U7947 ( .CLK(n8020), .C(n8031) );
  CKBD0 U7948 ( .CLK(n8021), .C(n8032) );
  CKBD0 U7949 ( .CLK(n8022), .C(n8033) );
  CKBD0 U7950 ( .CLK(n8023), .C(n8034) );
  CKBD0 U7951 ( .CLK(n8024), .C(n8035) );
  CKBD0 U7952 ( .CLK(n8025), .C(n8036) );
  CKBD0 U7953 ( .CLK(n8027), .C(n8037) );
  CKBD0 U7954 ( .CLK(n8030), .C(n8038) );
  CKBD0 U7955 ( .CLK(n8031), .C(n8039) );
  CKBD0 U7956 ( .CLK(n8032), .C(n8040) );
  CKBD0 U7957 ( .CLK(n8033), .C(n8041) );
  CKBD0 U7958 ( .CLK(n8034), .C(n8042) );
  BUFFD0 U7959 ( .I(n8035), .Z(n8043) );
  CKBD0 U7960 ( .CLK(n8036), .C(n8044) );
  CKBD0 U7961 ( .CLK(n8037), .C(n8045) );
  CKBD0 U7962 ( .CLK(n8038), .C(n8046) );
  CKBD0 U7963 ( .CLK(n8039), .C(n8047) );
  CKBD0 U7964 ( .CLK(n8040), .C(n8048) );
  BUFFD0 U7965 ( .I(n8041), .Z(n8049) );
  CKBD0 U7966 ( .CLK(n8042), .C(n8050) );
  CKBD0 U7967 ( .CLK(n8043), .C(n8051) );
  CKBD0 U7968 ( .CLK(n8044), .C(n8052) );
  BUFFD0 U7969 ( .I(n8045), .Z(n8053) );
  BUFFD0 U7970 ( .I(n8046), .Z(n8054) );
  CKBD0 U7971 ( .CLK(n8047), .C(n8055) );
  CKBD0 U7972 ( .CLK(n8048), .C(n8056) );
  CKBD0 U7973 ( .CLK(n8049), .C(n8057) );
  CKBD0 U7974 ( .CLK(n8050), .C(n8058) );
  CKBD0 U7975 ( .CLK(n8051), .C(n8059) );
  CKBD0 U7976 ( .CLK(n8052), .C(n8060) );
  CKBD0 U7977 ( .CLK(n8053), .C(n8061) );
  CKBD0 U7978 ( .CLK(n8054), .C(n8062) );
  BUFFD0 U7979 ( .I(n8055), .Z(n8063) );
  CKBD0 U7980 ( .CLK(n8056), .C(n8064) );
  CKBD0 U7981 ( .CLK(n8057), .C(n8065) );
  CKBD0 U7982 ( .CLK(n8058), .C(n8066) );
  CKBD0 U7983 ( .CLK(n8059), .C(n8067) );
  BUFFD0 U7984 ( .I(n8060), .Z(n8068) );
  CKBD0 U7985 ( .CLK(n8061), .C(n8069) );
  CKBD0 U7986 ( .CLK(n8062), .C(n8070) );
  CKBD0 U7987 ( .CLK(n8063), .C(n8071) );
  CKBD0 U7988 ( .CLK(n8064), .C(n8072) );
  CKBD0 U7989 ( .CLK(n8065), .C(n8073) );
  BUFFD0 U7990 ( .I(n8066), .Z(n8074) );
  CKBD0 U7991 ( .CLK(n8067), .C(n8075) );
  BUFFD0 U7992 ( .I(n7993), .Z(n8076) );
  BUFFD0 U7993 ( .I(n7994), .Z(n8077) );
  CKBD0 U7994 ( .CLK(n7997), .C(n8078) );
  BUFFD0 U7995 ( .I(n7995), .Z(n8079) );
  BUFFD0 U7996 ( .I(n7996), .Z(n8080) );
  CKBD0 U7997 ( .CLK(n8068), .C(n8081) );
  CKBD0 U7998 ( .CLK(n8069), .C(n8082) );
  CKBD0 U7999 ( .CLK(n8070), .C(n8083) );
  CKBD0 U8000 ( .CLK(n8071), .C(n8084) );
  BUFFD0 U8001 ( .I(n8072), .Z(n8085) );
  CKBD0 U8002 ( .CLK(n8073), .C(n8086) );
  CKBD0 U8003 ( .CLK(n8074), .C(n8087) );
  CKBD0 U8004 ( .CLK(n8075), .C(n8088) );
  BUFFD0 U8005 ( .I(n7998), .Z(n8089) );
  CKBD0 U8006 ( .CLK(n8000), .C(n8090) );
  CKBD0 U8007 ( .CLK(n8002), .C(n8091) );
  CKBD0 U8008 ( .CLK(n8001), .C(n8092) );
  CKBD0 U8009 ( .CLK(n8081), .C(n8093) );
  BUFFD0 U8010 ( .I(n8003), .Z(n8094) );
  CKBD0 U8011 ( .CLK(n8082), .C(n8095) );
  CKBD0 U8012 ( .CLK(n8083), .C(n8096) );
  CKBD0 U8013 ( .CLK(n8084), .C(n8097) );
  CKBD0 U8014 ( .CLK(n8085), .C(n8098) );
  CKBD0 U8015 ( .CLK(n8086), .C(n8099) );
  CKBD0 U8016 ( .CLK(n8087), .C(n8100) );
  CKBD0 U8017 ( .CLK(n8088), .C(n8101) );
  CKBD0 U8018 ( .CLK(n8004), .C(n8102) );
  CKBD0 U8019 ( .CLK(n8006), .C(n8103) );
  CKBD0 U8020 ( .CLK(n8007), .C(n8104) );
  CKBD0 U8021 ( .CLK(n8008), .C(n8105) );
  CKBD0 U8022 ( .CLK(n8093), .C(n8106) );
  CKBD0 U8023 ( .CLK(n8095), .C(n8107) );
  CKBD0 U8024 ( .CLK(n8096), .C(n8108) );
  CKBD0 U8025 ( .CLK(n8097), .C(n8109) );
  CKBD0 U8026 ( .CLK(n8098), .C(n8110) );
  CKBD0 U8027 ( .CLK(n8099), .C(n8111) );
  CKBD0 U8028 ( .CLK(n8100), .C(n8112) );
  CKBD0 U8029 ( .CLK(n8101), .C(n8113) );
  CKBD0 U8030 ( .CLK(n8010), .C(n8114) );
  BUFFD0 U8031 ( .I(n7964), .Z(n8115) );
  CKBD0 U8032 ( .CLK(n8011), .C(n8116) );
  CKBD0 U8033 ( .CLK(n8012), .C(n8117) );
  CKBD0 U8034 ( .CLK(n8106), .C(n8118) );
  CKBD0 U8035 ( .CLK(n8107), .C(n8119) );
  CKBD0 U8036 ( .CLK(n8108), .C(n8120) );
  CKBD0 U8037 ( .CLK(n8109), .C(n8121) );
  CKBD0 U8038 ( .CLK(n8110), .C(n8122) );
  CKBD0 U8039 ( .CLK(n8111), .C(n8123) );
  CKBD0 U8040 ( .CLK(n8112), .C(n8124) );
  CKBD0 U8041 ( .CLK(n8113), .C(n8125) );
  CKBD0 U8042 ( .CLK(n8013), .C(n8126) );
  CKBD0 U8043 ( .CLK(n8016), .C(n8127) );
  CKBD0 U8044 ( .CLK(n8118), .C(n8128) );
  CKBD0 U8045 ( .CLK(n8015), .C(n8129) );
  CKBD0 U8046 ( .CLK(n8119), .C(n8130) );
  CKBD0 U8047 ( .CLK(n8120), .C(n8131) );
  CKBD0 U8048 ( .CLK(n8121), .C(n8132) );
  CKBD0 U8049 ( .CLK(n8122), .C(n8133) );
  CKBD0 U8050 ( .CLK(n8123), .C(n8134) );
  CKBD0 U8051 ( .CLK(n8124), .C(n8135) );
  CKBD0 U8052 ( .CLK(n8125), .C(n8136) );
  CKBD0 U8053 ( .CLK(n8128), .C(n8137) );
  CKBD0 U8054 ( .CLK(n8026), .C(n8138) );
  CKBD0 U8055 ( .CLK(n8130), .C(n8139) );
  BUFFD0 U8056 ( .I(n8991), .Z(n8140) );
  BUFFD0 U8057 ( .I(n8028), .Z(n8141) );
  CKBD0 U8058 ( .CLK(n8131), .C(n8142) );
  CKBD0 U8059 ( .CLK(n8132), .C(n8143) );
  CKBD0 U8060 ( .CLK(n8133), .C(n8144) );
  CKBD0 U8061 ( .CLK(n8134), .C(n8145) );
  CKBD0 U8062 ( .CLK(n8135), .C(n8146) );
  CKBD0 U8063 ( .CLK(n8136), .C(n8147) );
  CKBD0 U8064 ( .CLK(n8137), .C(n8148) );
  CKBD0 U8065 ( .CLK(n8139), .C(n8149) );
  CKBD0 U8066 ( .CLK(n8076), .C(n8150) );
  CKBD0 U8067 ( .CLK(n8077), .C(n8151) );
  BUFFD0 U8068 ( .I(n8547), .Z(n8152) );
  CKBD0 U8069 ( .CLK(n8079), .C(n8153) );
  CKBD0 U8070 ( .CLK(n8080), .C(n8154) );
  CKBD0 U8071 ( .CLK(n8142), .C(n8155) );
  CKBD0 U8072 ( .CLK(n8143), .C(n8156) );
  CKBD0 U8073 ( .CLK(n8089), .C(n8157) );
  BUFFD0 U8074 ( .I(n8090), .Z(n8158) );
  CKBD0 U8075 ( .CLK(n8092), .C(n8159) );
  BUFFD0 U8076 ( .I(n8091), .Z(n8160) );
  CKBD0 U8077 ( .CLK(n8094), .C(n8161) );
  BUFFD0 U8078 ( .I(n8207), .Z(n8162) );
  CKBD0 U8079 ( .CLK(n8144), .C(n8163) );
  CKBD0 U8080 ( .CLK(n8103), .C(n8164) );
  CKBD0 U8081 ( .CLK(n8104), .C(n8165) );
  BUFFD0 U8082 ( .I(n8116), .Z(n8166) );
  CKBD0 U8083 ( .CLK(n8105), .C(n8167) );
  CKBD0 U8084 ( .CLK(n8115), .C(n8168) );
  BUFFD0 U8085 ( .I(n8114), .Z(n8169) );
  CKBD0 U8086 ( .CLK(n8145), .C(n8170) );
  CKBD0 U8087 ( .CLK(n8117), .C(n8171) );
  BUFFD0 U8088 ( .I(n8419), .Z(n8172) );
  CKBD0 U8089 ( .CLK(n8126), .C(n8173) );
  CKBD0 U8090 ( .CLK(n8146), .C(n8174) );
  CKBD0 U8091 ( .CLK(n8129), .C(n8175) );
  BUFFD0 U8092 ( .I(n8147), .Z(n8176) );
  CKBD0 U8093 ( .CLK(n8148), .C(n8177) );
  BUFFD0 U8094 ( .I(n8138), .Z(n8178) );
  BUFFD0 U8095 ( .I(n8149), .Z(n8179) );
  BUFFD0 U8096 ( .I(n8029), .Z(n8180) );
  CKBD0 U8097 ( .CLK(n8141), .C(n8181) );
  BUFFD0 U8098 ( .I(n8446), .Z(n8182) );
  BUFFD0 U8099 ( .I(n8150), .Z(n8183) );
  CKBD0 U8100 ( .CLK(n8155), .C(n8184) );
  CKBD0 U8101 ( .CLK(n8156), .C(n8185) );
  CKBD0 U8102 ( .CLK(n8163), .C(n8186) );
  CKBD0 U8103 ( .CLK(n8170), .C(n8187) );
  CKBD0 U8104 ( .CLK(n8174), .C(n8188) );
  CKBD0 U8105 ( .CLK(n8176), .C(n8189) );
  CKBD0 U8106 ( .CLK(n8177), .C(n8190) );
  CKBD0 U8107 ( .CLK(n8179), .C(n8191) );
  BUFFD0 U8108 ( .I(n8078), .Z(n8192) );
  BUFFD0 U8109 ( .I(n8153), .Z(n8193) );
  BUFFD0 U8110 ( .I(n8154), .Z(n8194) );
  BUFFD0 U8111 ( .I(n8184), .Z(n8195) );
  BUFFD0 U8112 ( .I(n8185), .Z(n8196) );
  BUFFD0 U8113 ( .I(n8806), .Z(n8197) );
  BUFFD0 U8114 ( .I(n8157), .Z(n8198) );
  CKBD0 U8115 ( .CLK(n8158), .C(n8199) );
  CKBD0 U8116 ( .CLK(n8186), .C(n8200) );
  BUFFD0 U8117 ( .I(n8187), .Z(n8201) );
  CKBD0 U8118 ( .CLK(n8188), .C(n8202) );
  CKBD0 U8119 ( .CLK(n8189), .C(n8203) );
  CKBD0 U8120 ( .CLK(n8190), .C(n8204) );
  CKBD0 U8121 ( .CLK(n8191), .C(n8205) );
  CKBD0 U8122 ( .CLK(n8160), .C(n8206) );
  BUFFD0 U8123 ( .I(n8962), .Z(n8207) );
  BUFFD0 U8124 ( .I(n8161), .Z(n8208) );
  CKBD0 U8125 ( .CLK(n8195), .C(n8209) );
  CKBD0 U8126 ( .CLK(n8196), .C(n8210) );
  BUFFD0 U8127 ( .I(n8295), .Z(n8211) );
  BUFFD0 U8128 ( .I(n8164), .Z(n8212) );
  CKBD0 U8129 ( .CLK(n8200), .C(n8213) );
  CKBD0 U8130 ( .CLK(n8201), .C(n8214) );
  CKBD0 U8131 ( .CLK(n8202), .C(n8215) );
  CKBD0 U8132 ( .CLK(n8203), .C(n8216) );
  CKBD0 U8133 ( .CLK(n8204), .C(n8217) );
  CKBD0 U8134 ( .CLK(n8205), .C(n8218) );
  CKBD0 U8135 ( .CLK(n8166), .C(n8219) );
  BUFFD0 U8136 ( .I(n8165), .Z(n8220) );
  CKBD0 U8137 ( .CLK(n8169), .C(n8221) );
  BUFFD0 U8138 ( .I(n8168), .Z(n8222) );
  BUFFD0 U8139 ( .I(n8301), .Z(n8223) );
  BUFFD0 U8140 ( .I(n8511), .Z(n8224) );
  CKBD0 U8141 ( .CLK(n8209), .C(n8225) );
  CKBD0 U8142 ( .CLK(n8210), .C(n8226) );
  BUFFD0 U8143 ( .I(n8127), .Z(n8227) );
  BUFFD0 U8144 ( .I(n8213), .Z(n8228) );
  CKBD0 U8145 ( .CLK(n8214), .C(n8229) );
  BUFFD0 U8146 ( .I(n8215), .Z(n8230) );
  CKBD0 U8147 ( .CLK(n8216), .C(n8231) );
  BUFFD0 U8148 ( .I(n8217), .Z(n8232) );
  CKBD0 U8149 ( .CLK(n8218), .C(n8233) );
  BUFFD0 U8150 ( .I(n8311), .Z(n8234) );
  CKBD0 U8151 ( .CLK(n8225), .C(n8235) );
  CKBD0 U8152 ( .CLK(n8226), .C(n8236) );
  CKBD0 U8153 ( .CLK(n8228), .C(n8237) );
  CKBD0 U8154 ( .CLK(n8229), .C(n8238) );
  CKBD0 U8155 ( .CLK(n8230), .C(n8239) );
  CKBD0 U8156 ( .CLK(n8231), .C(n8240) );
  CKBD0 U8157 ( .CLK(n8178), .C(n8241) );
  CKBD0 U8158 ( .CLK(n8180), .C(n8242) );
  BUFFD0 U8159 ( .I(n8181), .Z(n8243) );
  CKBD0 U8160 ( .CLK(n8232), .C(n8244) );
  CKBD0 U8161 ( .CLK(n8233), .C(n8245) );
  CKBD0 U8162 ( .CLK(n8235), .C(n8246) );
  CKBD0 U8163 ( .CLK(n8236), .C(n8247) );
  CKBD0 U8164 ( .CLK(n8237), .C(n8248) );
  CKBD0 U8165 ( .CLK(n8238), .C(n8249) );
  CKBD0 U8166 ( .CLK(n8239), .C(n8250) );
  CKBD0 U8167 ( .CLK(n8240), .C(n8251) );
  CKBD0 U8168 ( .CLK(n8183), .C(n8252) );
  BUFFD0 U8169 ( .I(n8151), .Z(n8253) );
  CKBD0 U8170 ( .CLK(n8192), .C(n8254) );
  CKBD0 U8171 ( .CLK(n8193), .C(n8255) );
  CKBD0 U8172 ( .CLK(n8194), .C(n8256) );
  CKBD0 U8173 ( .CLK(n8244), .C(n8257) );
  CKBD0 U8174 ( .CLK(n8245), .C(n8258) );
  CKBD0 U8175 ( .CLK(n8246), .C(n8259) );
  CKBD0 U8176 ( .CLK(n8247), .C(n8260) );
  CKBD0 U8177 ( .CLK(n8248), .C(n8261) );
  CKBD0 U8178 ( .CLK(n8249), .C(n8262) );
  CKBD0 U8179 ( .CLK(n8250), .C(n8263) );
  CKBD0 U8180 ( .CLK(n8251), .C(n8264) );
  CKBD0 U8181 ( .CLK(n8198), .C(n8265) );
  BUFFD0 U8182 ( .I(n8347), .Z(n8266) );
  BUFFD0 U8183 ( .I(n8159), .Z(n8267) );
  BUFFD0 U8184 ( .I(n8199), .Z(n8268) );
  BUFFD0 U8185 ( .I(n8219), .Z(n8269) );
  CKBD0 U8186 ( .CLK(n8257), .C(n8270) );
  CKBD0 U8187 ( .CLK(n8208), .C(n8271) );
  CKBD0 U8188 ( .CLK(n8258), .C(n8272) );
  CKBD0 U8189 ( .CLK(n8259), .C(n8273) );
  CKBD0 U8190 ( .CLK(n8260), .C(n8274) );
  CKBD0 U8191 ( .CLK(n8261), .C(n8275) );
  CKBD0 U8192 ( .CLK(n8262), .C(n8276) );
  CKBD0 U8193 ( .CLK(n8263), .C(n8277) );
  CKBD0 U8194 ( .CLK(n8264), .C(n8278) );
  CKBD0 U8195 ( .CLK(n8270), .C(n8279) );
  CKBD0 U8196 ( .CLK(n8272), .C(n8280) );
  CKBD0 U8197 ( .CLK(n8273), .C(n8281) );
  CKBD0 U8198 ( .CLK(n8274), .C(n8282) );
  CKBD0 U8199 ( .CLK(n8275), .C(n8283) );
  CKBD0 U8200 ( .CLK(n8276), .C(n8284) );
  CKBD0 U8201 ( .CLK(n8277), .C(n8285) );
  CKBD0 U8202 ( .CLK(n8278), .C(n8286) );
  CKBD0 U8203 ( .CLK(n8279), .C(n8287) );
  CKBD0 U8204 ( .CLK(n8280), .C(n8288) );
  CKBD0 U8205 ( .CLK(n8281), .C(n8289) );
  CKBD0 U8206 ( .CLK(n8282), .C(n8290) );
  CKBD0 U8207 ( .CLK(n8283), .C(n8291) );
  CKBD0 U8208 ( .CLK(n8284), .C(n8292) );
  BUFFD0 U8209 ( .I(n8102), .Z(n8293) );
  CKBD0 U8210 ( .CLK(n8285), .C(n8294) );
  BUFFD0 U8211 ( .I(n8723), .Z(n8295) );
  CKBD0 U8212 ( .CLK(n8212), .C(n8296) );
  CKBD0 U8213 ( .CLK(n8220), .C(n8297) );
  BUFFD0 U8214 ( .I(n8173), .Z(n8298) );
  BUFFD0 U8215 ( .I(n8421), .Z(n8299) );
  BUFFD0 U8216 ( .I(n8286), .Z(n8300) );
  BUFFD0 U8217 ( .I(n8582), .Z(n8301) );
  CKBD0 U8218 ( .CLK(n8287), .C(n8302) );
  BUFFD0 U8219 ( .I(n8288), .Z(n8303) );
  CKBD0 U8220 ( .CLK(n8289), .C(n8304) );
  CKBD0 U8221 ( .CLK(n8290), .C(n8305) );
  CKBD0 U8222 ( .CLK(n8291), .C(n8306) );
  CKBD0 U8223 ( .CLK(n8292), .C(n8307) );
  CKBD0 U8224 ( .CLK(n8294), .C(n8308) );
  CKBD0 U8225 ( .CLK(n8222), .C(n8309) );
  CKBD0 U8226 ( .CLK(n8300), .C(n8310) );
  BUFFD0 U8227 ( .I(n8418), .Z(n8311) );
  CKBD0 U8228 ( .CLK(n8302), .C(n8312) );
  CKBD0 U8229 ( .CLK(n8303), .C(n8313) );
  BUFFD0 U8230 ( .I(n8304), .Z(n8314) );
  CKBD0 U8231 ( .CLK(n8305), .C(n8315) );
  CKBD0 U8232 ( .CLK(n8306), .C(n8316) );
  BUFFD0 U8233 ( .I(n8307), .Z(n8317) );
  CKBD0 U8234 ( .CLK(n8308), .C(n8318) );
  CKBD0 U8235 ( .CLK(n8227), .C(n8319) );
  CKBD0 U8236 ( .CLK(n8310), .C(n8320) );
  CKBD0 U8237 ( .CLK(n8312), .C(n8321) );
  CKBD0 U8238 ( .CLK(n8313), .C(n8322) );
  CKBD0 U8239 ( .CLK(n8314), .C(n8323) );
  BUFFD0 U8240 ( .I(n8315), .Z(n8324) );
  CKBD0 U8241 ( .CLK(n8316), .C(n8325) );
  CKBD0 U8242 ( .CLK(n8317), .C(n8326) );
  CKBD0 U8243 ( .CLK(n8318), .C(n8327) );
  CKBD0 U8244 ( .CLK(n8320), .C(n8328) );
  CKBD0 U8245 ( .CLK(n8321), .C(n8329) );
  BUFFD0 U8246 ( .I(n8730), .Z(n8330) );
  CKBD0 U8247 ( .CLK(n8322), .C(n8331) );
  BUFFD0 U8248 ( .I(n8242), .Z(n8332) );
  CKBD0 U8249 ( .CLK(n8243), .C(n8333) );
  CKBD0 U8250 ( .CLK(n8253), .C(n8334) );
  BUFFD0 U8251 ( .I(n8449), .Z(n8335) );
  BUFFD0 U8252 ( .I(n8252), .Z(n8336) );
  CKBD0 U8253 ( .CLK(n8323), .C(n8337) );
  CKBD0 U8254 ( .CLK(n8324), .C(n8338) );
  BUFFD0 U8255 ( .I(n8254), .Z(n8339) );
  BUFFD0 U8256 ( .I(n8325), .Z(n8340) );
  CKBD0 U8257 ( .CLK(n8326), .C(n8341) );
  CKBD0 U8258 ( .CLK(n8327), .C(n8342) );
  CKBD0 U8259 ( .CLK(n8328), .C(n8343) );
  BUFFD0 U8260 ( .I(n8329), .Z(n8344) );
  CKBD0 U8261 ( .CLK(n8331), .C(n8345) );
  BUFFD0 U8262 ( .I(n8256), .Z(n8346) );
  BUFFD0 U8263 ( .I(n8805), .Z(n8347) );
  CKBD0 U8264 ( .CLK(n8267), .C(n8348) );
  BUFFD0 U8265 ( .I(n8265), .Z(n8349) );
  CKBD0 U8266 ( .CLK(n8337), .C(n8350) );
  CKBD0 U8267 ( .CLK(n8268), .C(n8351) );
  CKBD0 U8268 ( .CLK(n8338), .C(n8352) );
  CKBD0 U8269 ( .CLK(n8340), .C(n8353) );
  CKBD0 U8270 ( .CLK(n8341), .C(n8354) );
  BUFFD0 U8271 ( .I(n8342), .Z(n8355) );
  CKBD0 U8272 ( .CLK(n8343), .C(n8356) );
  CKBD0 U8273 ( .CLK(n8344), .C(n8357) );
  CKBD0 U8274 ( .CLK(n8345), .C(n8358) );
  BUFFD0 U8275 ( .I(n8618), .Z(n8359) );
  CKBD0 U8276 ( .CLK(n8269), .C(n8360) );
  CKBD0 U8277 ( .CLK(n8350), .C(n8361) );
  CKBD0 U8278 ( .CLK(n8352), .C(n8362) );
  CKBD0 U8279 ( .CLK(n8353), .C(n8363) );
  CKBD0 U8280 ( .CLK(n8354), .C(n8364) );
  CKBD0 U8281 ( .CLK(n8355), .C(n8365) );
  CKBD0 U8282 ( .CLK(n8356), .C(n8366) );
  CKBD0 U8283 ( .CLK(n8357), .C(n8367) );
  CKBD0 U8284 ( .CLK(n8358), .C(n8368) );
  CKBD0 U8285 ( .CLK(n8361), .C(n8369) );
  CKBD0 U8286 ( .CLK(n8362), .C(n8370) );
  CKBD0 U8287 ( .CLK(n8363), .C(n8371) );
  CKBD0 U8288 ( .CLK(n8364), .C(n8372) );
  CKBD0 U8289 ( .CLK(n8365), .C(n8373) );
  CKBD0 U8290 ( .CLK(n8366), .C(n8374) );
  CKBD0 U8291 ( .CLK(n8367), .C(n8375) );
  CKBD0 U8292 ( .CLK(n8368), .C(n8376) );
  CKBD0 U8293 ( .CLK(n8369), .C(n8377) );
  CKBD0 U8294 ( .CLK(n8370), .C(n8378) );
  CKBD0 U8295 ( .CLK(n8371), .C(n8379) );
  CKBD0 U8296 ( .CLK(n8372), .C(n8380) );
  CKBD0 U8297 ( .CLK(n8373), .C(n8381) );
  CKBD0 U8298 ( .CLK(n8374), .C(n8382) );
  CKBD0 U8299 ( .CLK(n8375), .C(n8383) );
  CKBD0 U8300 ( .CLK(n8376), .C(n8384) );
  CKBD0 U8301 ( .CLK(n8377), .C(n8385) );
  CKBD0 U8302 ( .CLK(n8378), .C(n8386) );
  CKBD0 U8303 ( .CLK(n8379), .C(n8387) );
  CKBD0 U8304 ( .CLK(n8380), .C(n8388) );
  CKBD0 U8305 ( .CLK(n8381), .C(n8389) );
  CKBD0 U8306 ( .CLK(n8382), .C(n8390) );
  CKBD0 U8307 ( .CLK(n8383), .C(n8391) );
  CKBD0 U8308 ( .CLK(n8293), .C(n8392) );
  CKBD0 U8309 ( .CLK(n8384), .C(n8393) );
  CKBD0 U8310 ( .CLK(n8385), .C(n8394) );
  CKBD0 U8311 ( .CLK(n8386), .C(n8395) );
  CKBD0 U8312 ( .CLK(n8387), .C(n8396) );
  CKBD0 U8313 ( .CLK(n8388), .C(n8397) );
  CKBD0 U8314 ( .CLK(n8389), .C(n8398) );
  CKBD0 U8315 ( .CLK(n8390), .C(n8399) );
  CKBD0 U8316 ( .CLK(n8391), .C(n8400) );
  CKBD0 U8317 ( .CLK(n8393), .C(n8401) );
  CKBD0 U8318 ( .CLK(n8394), .C(n8402) );
  CKBD0 U8319 ( .CLK(n8395), .C(n8403) );
  CKBD0 U8320 ( .CLK(n8396), .C(n8404) );
  CKBD0 U8321 ( .CLK(n8397), .C(n8405) );
  CKBD0 U8322 ( .CLK(n8398), .C(n8406) );
  CKBD0 U8323 ( .CLK(n8399), .C(n8407) );
  CKBD0 U8324 ( .CLK(n8400), .C(n8408) );
  BUFFD0 U8325 ( .I(n8401), .Z(n8409) );
  CKBD0 U8326 ( .CLK(n8402), .C(n8410) );
  CKBD0 U8327 ( .CLK(n8403), .C(n8411) );
  CKBD0 U8328 ( .CLK(n8404), .C(n8412) );
  CKBD0 U8329 ( .CLK(n8405), .C(n8413) );
  CKBD0 U8330 ( .CLK(n8406), .C(n8414) );
  BUFFD0 U8331 ( .I(n8514), .Z(n8415) );
  BUFFD0 U8332 ( .I(n8167), .Z(n8416) );
  BUFFD0 U8333 ( .I(n8516), .Z(n8417) );
  BUFFD0 U8334 ( .I(n8503), .Z(n8418) );
  BUFFD0 U8335 ( .I(n8601), .Z(n8419) );
  CKBD0 U8336 ( .CLK(n8298), .C(n8420) );
  BUFFD0 U8337 ( .I(n8632), .Z(n8421) );
  BUFFD0 U8338 ( .I(n8407), .Z(n8422) );
  CKBD0 U8339 ( .CLK(n8408), .C(n8423) );
  CKBD0 U8340 ( .CLK(n8409), .C(n8424) );
  BUFFD0 U8341 ( .I(n8410), .Z(n8425) );
  CKBD0 U8342 ( .CLK(n8411), .C(n8426) );
  CKBD0 U8343 ( .CLK(n8412), .C(n8427) );
  BUFFD0 U8344 ( .I(n8413), .Z(n8428) );
  CKBD0 U8345 ( .CLK(n8414), .C(n8429) );
  BUFFD0 U8346 ( .I(n8171), .Z(n8430) );
  BUFFD0 U8347 ( .I(n8309), .Z(n8431) );
  CKBD0 U8348 ( .CLK(n8422), .C(n8432) );
  CKBD0 U8349 ( .CLK(n8423), .C(n8433) );
  CKBD0 U8350 ( .CLK(n8424), .C(n8434) );
  CKBD0 U8351 ( .CLK(n8425), .C(n8435) );
  BUFFD0 U8352 ( .I(n8426), .Z(n8436) );
  CKBD0 U8353 ( .CLK(n8427), .C(n8437) );
  CKBD0 U8354 ( .CLK(n8428), .C(n8438) );
  CKBD0 U8355 ( .CLK(n8429), .C(n8439) );
  CKBD0 U8356 ( .CLK(n8432), .C(n8440) );
  CKBD0 U8357 ( .CLK(n8433), .C(n8441) );
  BUFFD0 U8358 ( .I(n8241), .Z(n8442) );
  CKBD0 U8359 ( .CLK(n8434), .C(n8443) );
  BUFFD0 U8360 ( .I(n8989), .Z(n8444) );
  CKBD0 U8361 ( .CLK(n8332), .C(n8445) );
  BUFFD0 U8362 ( .I(n8988), .Z(n8446) );
  CKBD0 U8363 ( .CLK(n8435), .C(n8447) );
  CKBD0 U8364 ( .CLK(n8436), .C(n8448) );
  BUFFD0 U8365 ( .I(n8993), .Z(n8449) );
  CKBD0 U8366 ( .CLK(n8437), .C(n8450) );
  CKBD0 U8367 ( .CLK(n8438), .C(n8451) );
  BUFFD0 U8368 ( .I(n8439), .Z(n8452) );
  CKBD0 U8369 ( .CLK(n8440), .C(n8453) );
  BUFFD0 U8370 ( .I(n8441), .Z(n8454) );
  CKBD0 U8371 ( .CLK(n8443), .C(n8455) );
  CKBD0 U8372 ( .CLK(n8336), .C(n8456) );
  CKBD0 U8373 ( .CLK(n8339), .C(n8457) );
  CKBD0 U8374 ( .CLK(n8346), .C(n8458) );
  CKBD0 U8375 ( .CLK(n8447), .C(n8459) );
  BUFFD0 U8376 ( .I(n8360), .Z(n8460) );
  CKBD0 U8377 ( .CLK(n8448), .C(n8461) );
  BUFFD0 U8378 ( .I(n8450), .Z(n8462) );
  CKBD0 U8379 ( .CLK(n8451), .C(n8463) );
  CKBD0 U8380 ( .CLK(n8452), .C(n8464) );
  CKBD0 U8381 ( .CLK(n8453), .C(n8465) );
  CKBD0 U8382 ( .CLK(n8454), .C(n8466) );
  CKBD0 U8383 ( .CLK(n8455), .C(n8467) );
  BUFFD0 U8384 ( .I(n8206), .Z(n8468) );
  CKBD0 U8385 ( .CLK(n8349), .C(n8469) );
  CKBD0 U8386 ( .CLK(n8459), .C(n8470) );
  CKBD0 U8387 ( .CLK(n8461), .C(n8471) );
  CKBD0 U8388 ( .CLK(n8462), .C(n8472) );
  CKBD0 U8389 ( .CLK(n8463), .C(n8473) );
  CKBD0 U8390 ( .CLK(n8464), .C(n8474) );
  CKBD0 U8391 ( .CLK(n8465), .C(n8475) );
  CKBD0 U8392 ( .CLK(n8466), .C(n8476) );
  CKBD0 U8393 ( .CLK(n8467), .C(n8477) );
  CKBD0 U8394 ( .CLK(n8470), .C(n8478) );
  CKBD0 U8395 ( .CLK(n8471), .C(n8479) );
  CKBD0 U8396 ( .CLK(n8472), .C(n8480) );
  CKBD0 U8397 ( .CLK(n8473), .C(n8481) );
  CKBD0 U8398 ( .CLK(n8474), .C(n8482) );
  CKBD0 U8399 ( .CLK(n8475), .C(n8483) );
  CKBD0 U8400 ( .CLK(n8476), .C(n8484) );
  CKBD0 U8401 ( .CLK(n8477), .C(n8485) );
  CKBD0 U8402 ( .CLK(n8478), .C(n8486) );
  CKBD0 U8403 ( .CLK(n8479), .C(n8487) );
  CKBD0 U8404 ( .CLK(n8480), .C(n8488) );
  CKBD0 U8405 ( .CLK(n8481), .C(n8489) );
  CKBD0 U8406 ( .CLK(n8482), .C(n8490) );
  CKBD0 U8407 ( .CLK(n8483), .C(n8491) );
  CKBD0 U8408 ( .CLK(n8484), .C(n8492) );
  CKBD0 U8409 ( .CLK(n8485), .C(n8493) );
  CKBD0 U8410 ( .CLK(n8486), .C(n8494) );
  CKBD0 U8411 ( .CLK(n8487), .C(n8495) );
  CKBD0 U8412 ( .CLK(n8488), .C(n8496) );
  CKBD0 U8413 ( .CLK(n8489), .C(n8497) );
  CKBD0 U8414 ( .CLK(n8490), .C(n8498) );
  CKBD0 U8415 ( .CLK(n8491), .C(n8499) );
  BUFFD0 U8416 ( .I(n8348), .Z(n8500) );
  CKBD0 U8417 ( .CLK(n8492), .C(n8501) );
  BUFFD0 U8418 ( .I(n8351), .Z(n8502) );
  BUFFD0 U8419 ( .I(n8980), .Z(n8503) );
  CKBD0 U8420 ( .CLK(n8493), .C(n8504) );
  CKBD0 U8421 ( .CLK(n8494), .C(n8505) );
  CKBD0 U8422 ( .CLK(n8495), .C(n8506) );
  CKBD0 U8423 ( .CLK(n8496), .C(n8507) );
  CKBD0 U8424 ( .CLK(n8497), .C(n8508) );
  CKBD0 U8425 ( .CLK(n8498), .C(n8509) );
  CKBD0 U8426 ( .CLK(n8499), .C(n8510) );
  BUFFD0 U8427 ( .I(n8559), .Z(n8511) );
  BUFFD0 U8428 ( .I(n8319), .Z(n8512) );
  BUFFD0 U8429 ( .I(n8271), .Z(n8513) );
  BUFFD0 U8430 ( .I(n8720), .Z(n8514) );
  BUFFD0 U8431 ( .I(n8392), .Z(n8515) );
  BUFFD0 U8432 ( .I(n8577), .Z(n8516) );
  CKBD0 U8433 ( .CLK(n8416), .C(n8517) );
  CKBD0 U8434 ( .CLK(n8501), .C(n8518) );
  CKBD0 U8435 ( .CLK(n8504), .C(n8519) );
  CKBD0 U8436 ( .CLK(n8506), .C(n8520) );
  CKBD0 U8437 ( .CLK(n8505), .C(n8521) );
  CKBD0 U8438 ( .CLK(n8507), .C(n8522) );
  CKBD0 U8439 ( .CLK(n8508), .C(n8523) );
  CKBD0 U8440 ( .CLK(n8509), .C(n8524) );
  CKBD0 U8441 ( .CLK(n8510), .C(n8525) );
  BUFFD0 U8442 ( .I(n8221), .Z(n8526) );
  CKBD0 U8443 ( .CLK(n8430), .C(n8527) );
  CKBD0 U8444 ( .CLK(n8431), .C(n8528) );
  CKBD0 U8445 ( .CLK(n8518), .C(n8529) );
  CKBD0 U8446 ( .CLK(n8519), .C(n8530) );
  BUFFD0 U8447 ( .I(n8520), .Z(n8531) );
  CKBD0 U8448 ( .CLK(n8521), .C(n8532) );
  CKBD0 U8449 ( .CLK(n8522), .C(n8533) );
  CKBD0 U8450 ( .CLK(n8442), .C(n8534) );
  BUFFD0 U8451 ( .I(n8333), .Z(n8535) );
  BUFFD0 U8452 ( .I(n8445), .Z(n8536) );
  CKBD0 U8453 ( .CLK(n8523), .C(n8537) );
  CKBD0 U8454 ( .CLK(n8524), .C(n8538) );
  CKBD0 U8455 ( .CLK(n8525), .C(n8539) );
  CKBD0 U8456 ( .CLK(n8529), .C(n8540) );
  BUFFD0 U8457 ( .I(n8530), .Z(n8541) );
  BUFFD0 U8458 ( .I(n8532), .Z(n8542) );
  CKBD0 U8459 ( .CLK(n8531), .C(n8543) );
  CKBD0 U8460 ( .CLK(n8533), .C(n8544) );
  BUFFD0 U8461 ( .I(n8537), .Z(n8545) );
  BUFFD0 U8462 ( .I(n8334), .Z(n8546) );
  BUFFD0 U8463 ( .I(n8594), .Z(n8547) );
  BUFFD0 U8464 ( .I(n8255), .Z(n8548) );
  BUFFD0 U8465 ( .I(n8456), .Z(n8549) );
  BUFFD0 U8466 ( .I(n8959), .Z(n8550) );
  CKBD0 U8467 ( .CLK(n8538), .C(n8551) );
  BUFFD0 U8468 ( .I(n8539), .Z(n8552) );
  BUFFD0 U8469 ( .I(n8540), .Z(n8553) );
  CKBD0 U8470 ( .CLK(n8541), .C(n8554) );
  CKBD0 U8471 ( .CLK(n8542), .C(n8555) );
  CKBD0 U8472 ( .CLK(n8543), .C(n8556) );
  CKBD0 U8473 ( .CLK(n8544), .C(n8557) );
  CKBD0 U8474 ( .CLK(n8545), .C(n8558) );
  BUFFD0 U8475 ( .I(n8592), .Z(n8559) );
  BUFFD0 U8476 ( .I(n8175), .Z(n8560) );
  BUFFD0 U8477 ( .I(n8804), .Z(n8561) );
  CKBD0 U8478 ( .CLK(n8460), .C(n8562) );
  CKBD0 U8479 ( .CLK(n8468), .C(n8563) );
  CKBD0 U8480 ( .CLK(n8500), .C(n8564) );
  CKBD0 U8481 ( .CLK(n8502), .C(n8565) );
  BUFFD0 U8482 ( .I(n8551), .Z(n8566) );
  CKBD0 U8483 ( .CLK(n8552), .C(n8567) );
  CKBD0 U8484 ( .CLK(n8553), .C(n8568) );
  CKBD0 U8485 ( .CLK(n8554), .C(n8569) );
  CKBD0 U8486 ( .CLK(n8555), .C(n8570) );
  CKBD0 U8487 ( .CLK(n8556), .C(n8571) );
  CKBD0 U8488 ( .CLK(n8557), .C(n8572) );
  CKBD0 U8489 ( .CLK(n8513), .C(n8573) );
  CKBD0 U8490 ( .CLK(n8512), .C(n8574) );
  CKBD0 U8491 ( .CLK(n8558), .C(n8575) );
  CKBD0 U8492 ( .CLK(n8515), .C(n8576) );
  BUFFD0 U8493 ( .I(n8955), .Z(n8577) );
  BUFFD0 U8494 ( .I(n8296), .Z(n8578) );
  BUFFD0 U8495 ( .I(n8517), .Z(n8579) );
  CKBD0 U8496 ( .CLK(n8526), .C(n8580) );
  CKBD0 U8497 ( .CLK(n8566), .C(n8581) );
  BUFFD0 U8498 ( .I(n8977), .Z(n8582) );
  BUFFD0 U8499 ( .I(n8528), .Z(n8583) );
  CKBD0 U8500 ( .CLK(n8567), .C(n8584) );
  CKBD0 U8501 ( .CLK(n8568), .C(n8585) );
  CKBD0 U8502 ( .CLK(n8569), .C(n8586) );
  BUFFD0 U8503 ( .I(n8534), .Z(n8587) );
  CKBD0 U8504 ( .CLK(n8535), .C(n8588) );
  CKBD0 U8505 ( .CLK(n8536), .C(n8589) );
  CKBD0 U8506 ( .CLK(n8570), .C(n8590) );
  CKBD0 U8507 ( .CLK(n8571), .C(n8591) );
  BUFFD0 U8508 ( .I(n8978), .Z(n8592) );
  CKBD0 U8509 ( .CLK(n8546), .C(n8593) );
  BUFFD0 U8510 ( .I(n8838), .Z(n8594) );
  CKBD0 U8511 ( .CLK(n8548), .C(n8595) );
  CKBD0 U8512 ( .CLK(n8549), .C(n8596) );
  BUFFD0 U8513 ( .I(n8562), .Z(n8597) );
  BUFFD0 U8514 ( .I(n8458), .Z(n8598) );
  BUFFD0 U8515 ( .I(n8572), .Z(n8599) );
  CKBD0 U8516 ( .CLK(n8560), .C(n8600) );
  BUFFD0 U8517 ( .I(n8982), .Z(n8601) );
  CKBD0 U8518 ( .CLK(n8575), .C(n8602) );
  CKBD0 U8519 ( .CLK(n8581), .C(n8603) );
  CKBD0 U8520 ( .CLK(n8584), .C(n8604) );
  CKBD0 U8521 ( .CLK(n8585), .C(n8605) );
  CKBD0 U8522 ( .CLK(n8586), .C(n8606) );
  CKBD0 U8523 ( .CLK(n8590), .C(n8607) );
  CKBD0 U8524 ( .CLK(n8591), .C(n8608) );
  CKBD0 U8525 ( .CLK(n8599), .C(n8609) );
  CKBD0 U8526 ( .CLK(n8602), .C(n8610) );
  CKBD0 U8527 ( .CLK(n8603), .C(n8611) );
  CKBD0 U8528 ( .CLK(n8604), .C(n8612) );
  CKBD0 U8529 ( .CLK(n8605), .C(n8613) );
  CKBD0 U8530 ( .CLK(n8606), .C(n8614) );
  BUFFD0 U8531 ( .I(n8469), .Z(n8615) );
  BUFFD0 U8532 ( .I(n8563), .Z(n8616) );
  BUFFD0 U8533 ( .I(n8564), .Z(n8617) );
  BUFFD0 U8534 ( .I(n8679), .Z(n8618) );
  BUFFD0 U8535 ( .I(n8565), .Z(n8619) );
  CKBD0 U8536 ( .CLK(n8607), .C(n8620) );
  CKBD0 U8537 ( .CLK(n8578), .C(n8621) );
  CKBD0 U8538 ( .CLK(n8608), .C(n8622) );
  BUFFD0 U8539 ( .I(n8576), .Z(n8623) );
  BUFFD0 U8540 ( .I(n8297), .Z(n8624) );
  CKBD0 U8541 ( .CLK(n8609), .C(n8625) );
  CKBD0 U8542 ( .CLK(n8610), .C(n8626) );
  CKBD0 U8543 ( .CLK(n8611), .C(n8627) );
  CKBD0 U8544 ( .CLK(n8612), .C(n8628) );
  CKBD0 U8545 ( .CLK(n8613), .C(n8629) );
  CKBD0 U8546 ( .CLK(n8614), .C(n8630) );
  CKBD0 U8547 ( .CLK(n8579), .C(n8631) );
  BUFFD0 U8548 ( .I(n8883), .Z(n8632) );
  BUFFD0 U8549 ( .I(n8527), .Z(n8633) );
  CKBD0 U8550 ( .CLK(n8620), .C(n8634) );
  CKBD0 U8551 ( .CLK(n8622), .C(n8635) );
  CKBD0 U8552 ( .CLK(n8583), .C(n8636) );
  CKBD0 U8553 ( .CLK(n8625), .C(n8637) );
  CKBD0 U8554 ( .CLK(n8626), .C(n8638) );
  CKBD0 U8555 ( .CLK(n8627), .C(n8639) );
  CKBD0 U8556 ( .CLK(n8628), .C(n8640) );
  CKBD0 U8557 ( .CLK(n8629), .C(n8641) );
  CKBD0 U8558 ( .CLK(n8630), .C(n8642) );
  CKBD0 U8559 ( .CLK(n8634), .C(n8643) );
  CKBD0 U8560 ( .CLK(n8635), .C(n8644) );
  CKBD0 U8561 ( .CLK(n8637), .C(n8645) );
  CKBD0 U8562 ( .CLK(n8638), .C(n8646) );
  CKBD0 U8563 ( .CLK(n8639), .C(n8647) );
  CKBD0 U8564 ( .CLK(n8640), .C(n8648) );
  CKBD0 U8565 ( .CLK(n8587), .C(n8649) );
  BUFFD0 U8566 ( .I(n8420), .Z(n8650) );
  CKBD0 U8567 ( .CLK(n8641), .C(n8651) );
  CKBD0 U8568 ( .CLK(n8642), .C(n8652) );
  CKBD0 U8569 ( .CLK(n8643), .C(n8653) );
  CKBD0 U8570 ( .CLK(n8644), .C(n8654) );
  CKBD0 U8571 ( .CLK(n8645), .C(n8655) );
  CKBD0 U8572 ( .CLK(n8646), .C(n8656) );
  CKBD0 U8573 ( .CLK(n8647), .C(n8657) );
  CKBD0 U8574 ( .CLK(n8648), .C(n8658) );
  BUFFD0 U8575 ( .I(n8588), .Z(n8659) );
  BUFFD0 U8576 ( .I(n8589), .Z(n8660) );
  BUFFD0 U8577 ( .I(n8600), .Z(n8661) );
  BUFFD0 U8578 ( .I(n8593), .Z(n8662) );
  BUFFD0 U8579 ( .I(n8457), .Z(n8663) );
  BUFFD0 U8580 ( .I(n8574), .Z(n8664) );
  BUFFD0 U8581 ( .I(n8595), .Z(n8665) );
  CKBD0 U8582 ( .CLK(n8597), .C(n8666) );
  BUFFD0 U8583 ( .I(n8596), .Z(n8667) );
  CKBD0 U8584 ( .CLK(n8651), .C(n8668) );
  CKBD0 U8585 ( .CLK(n8598), .C(n8669) );
  BUFFD0 U8586 ( .I(n8653), .Z(n8670) );
  CKBD0 U8587 ( .CLK(n8652), .C(n8671) );
  CKBD0 U8588 ( .CLK(n8654), .C(n8672) );
  CKBD0 U8589 ( .CLK(n8655), .C(n8673) );
  CKBD0 U8590 ( .CLK(n8656), .C(n8674) );
  CKBD0 U8591 ( .CLK(n8657), .C(n8675) );
  CKBD0 U8592 ( .CLK(n8658), .C(n8676) );
  CKBD0 U8593 ( .CLK(n8615), .C(n8677) );
  CKBD0 U8594 ( .CLK(n8616), .C(n8678) );
  BUFFD0 U8595 ( .I(n8961), .Z(n8679) );
  CKBD0 U8596 ( .CLK(n8617), .C(n8680) );
  CKBD0 U8597 ( .CLK(n8668), .C(n8681) );
  CKBD0 U8598 ( .CLK(n8671), .C(n8682) );
  CKBD0 U8599 ( .CLK(n8670), .C(n8683) );
  BUFFD0 U8600 ( .I(n8672), .Z(n8684) );
  CKBD0 U8601 ( .CLK(n8673), .C(n8685) );
  BUFFD0 U8602 ( .I(n8674), .Z(n8686) );
  CKBD0 U8603 ( .CLK(n8675), .C(n8687) );
  CKBD0 U8604 ( .CLK(n8676), .C(n8688) );
  CKBD0 U8605 ( .CLK(n8619), .C(n8689) );
  CKBD0 U8606 ( .CLK(n8681), .C(n8690) );
  BUFFD0 U8607 ( .I(n8682), .Z(n8691) );
  CKBD0 U8608 ( .CLK(n8683), .C(n8692) );
  CKBD0 U8609 ( .CLK(n8684), .C(n8693) );
  CKBD0 U8610 ( .CLK(n8685), .C(n8694) );
  CKBD0 U8611 ( .CLK(n8686), .C(n8695) );
  CKBD0 U8612 ( .CLK(n8687), .C(n8696) );
  BUFFD0 U8613 ( .I(n8688), .Z(n8697) );
  CKBD0 U8614 ( .CLK(n8690), .C(n8698) );
  CKBD0 U8615 ( .CLK(n8691), .C(n8699) );
  CKBD0 U8616 ( .CLK(n8692), .C(n8700) );
  CKBD0 U8617 ( .CLK(n8693), .C(n8701) );
  CKBD0 U8618 ( .CLK(n8694), .C(n8702) );
  CKBD0 U8619 ( .CLK(n8695), .C(n8703) );
  CKBD0 U8620 ( .CLK(n8696), .C(n8704) );
  CKBD0 U8621 ( .CLK(n8697), .C(n8705) );
  CKBD0 U8622 ( .CLK(n8698), .C(n8706) );
  CKBD0 U8623 ( .CLK(n8699), .C(n8707) );
  CKBD0 U8624 ( .CLK(n8700), .C(n8708) );
  CKBD0 U8625 ( .CLK(n8701), .C(n8709) );
  BUFFD0 U8626 ( .I(n8702), .Z(n8710) );
  CKBD0 U8627 ( .CLK(n8703), .C(n8711) );
  CKBD0 U8628 ( .CLK(n8704), .C(n8712) );
  CKBD0 U8629 ( .CLK(n8705), .C(n8713) );
  BUFFD0 U8630 ( .I(n8706), .Z(n8714) );
  CKBD0 U8631 ( .CLK(n8707), .C(n8715) );
  CKBD0 U8632 ( .CLK(n8708), .C(n8716) );
  CKBD0 U8633 ( .CLK(n8709), .C(n8717) );
  CKBD0 U8634 ( .CLK(n8710), .C(n8718) );
  CKBD0 U8635 ( .CLK(n8711), .C(n8719) );
  BUFFD0 U8636 ( .I(n8956), .Z(n8720) );
  CKBD0 U8637 ( .CLK(n8623), .C(n8721) );
  CKBD0 U8638 ( .CLK(n8624), .C(n8722) );
  BUFFD0 U8639 ( .I(n8810), .Z(n8723) );
  BUFFD0 U8640 ( .I(n8712), .Z(n8724) );
  BUFFD0 U8641 ( .I(n8580), .Z(n8725) );
  CKBD0 U8642 ( .CLK(n8633), .C(n8726) );
  BUFFD0 U8643 ( .I(n8636), .Z(n8727) );
  CKBD0 U8644 ( .CLK(n8713), .C(n8728) );
  CKBD0 U8645 ( .CLK(n8714), .C(n8729) );
  BUFFD0 U8646 ( .I(n8987), .Z(n8730) );
  CKBD0 U8647 ( .CLK(n8715), .C(n8731) );
  CKBD0 U8648 ( .CLK(n8650), .C(n8732) );
  CKBD0 U8649 ( .CLK(n8659), .C(n8733) );
  CKBD0 U8650 ( .CLK(n8660), .C(n8734) );
  BUFFD0 U8651 ( .I(n8666), .Z(n8735) );
  CKBD0 U8652 ( .CLK(n8716), .C(n8736) );
  CKBD0 U8653 ( .CLK(n8717), .C(n8737) );
  CKBD0 U8654 ( .CLK(n8718), .C(n8738) );
  CKBD0 U8655 ( .CLK(n8719), .C(n8739) );
  CKBD0 U8656 ( .CLK(n8724), .C(n8740) );
  CKBD0 U8657 ( .CLK(n8728), .C(n8741) );
  CKBD0 U8658 ( .CLK(n8729), .C(n8742) );
  CKBD0 U8659 ( .CLK(n8731), .C(n8743) );
  CKBD0 U8660 ( .CLK(n8662), .C(n8744) );
  CKBD0 U8661 ( .CLK(n8663), .C(n8745) );
  CKBD0 U8662 ( .CLK(n8736), .C(n8746) );
  CKBD0 U8663 ( .CLK(n8737), .C(n8747) );
  CKBD0 U8664 ( .CLK(n8738), .C(n8748) );
  CKBD0 U8665 ( .CLK(n8739), .C(n8749) );
  CKBD0 U8666 ( .CLK(n8740), .C(n8750) );
  CKBD0 U8667 ( .CLK(n8741), .C(n8751) );
  CKBD0 U8668 ( .CLK(n8742), .C(n8752) );
  CKBD0 U8669 ( .CLK(n8743), .C(n8753) );
  CKBD0 U8670 ( .CLK(n8746), .C(n8754) );
  CKBD0 U8671 ( .CLK(n8747), .C(n8755) );
  CKBD0 U8672 ( .CLK(n8748), .C(n8756) );
  CKBD0 U8673 ( .CLK(n8749), .C(n8757) );
  CKBD0 U8674 ( .CLK(n8750), .C(n8758) );
  CKBD0 U8675 ( .CLK(n8751), .C(n8759) );
  CKBD0 U8676 ( .CLK(n8752), .C(n8760) );
  CKBD0 U8677 ( .CLK(n8753), .C(n8761) );
  CKBD0 U8678 ( .CLK(n8754), .C(n8762) );
  CKBD0 U8679 ( .CLK(n8755), .C(n8763) );
  CKBD0 U8680 ( .CLK(n8756), .C(n8764) );
  CKBD0 U8681 ( .CLK(n8757), .C(n8765) );
  CKBD0 U8682 ( .CLK(n8758), .C(n8766) );
  CKBD0 U8683 ( .CLK(n8759), .C(n8767) );
  CKBD0 U8684 ( .CLK(n8760), .C(n8768) );
  CKBD0 U8685 ( .CLK(n8761), .C(n8769) );
  CKBD0 U8686 ( .CLK(n8762), .C(n8770) );
  CKBD0 U8687 ( .CLK(n8763), .C(n8771) );
  CKBD0 U8688 ( .CLK(n8764), .C(n8772) );
  CKBD0 U8689 ( .CLK(n8765), .C(n8773) );
  CKBD0 U8690 ( .CLK(n8766), .C(n8774) );
  CKBD0 U8691 ( .CLK(n8767), .C(n8775) );
  CKBD0 U8692 ( .CLK(n8768), .C(n8776) );
  CKBD0 U8693 ( .CLK(n8661), .C(n8777) );
  CKBD0 U8694 ( .CLK(n8664), .C(n8778) );
  CKBD0 U8695 ( .CLK(n8665), .C(n8779) );
  BUFFD0 U8696 ( .I(n8770), .Z(n8780) );
  CKBD0 U8697 ( .CLK(n8769), .C(n8781) );
  CKBD0 U8698 ( .CLK(n8771), .C(n8782) );
  CKBD0 U8699 ( .CLK(n8772), .C(n8783) );
  BUFFD0 U8700 ( .I(n8773), .Z(n8784) );
  CKBD0 U8701 ( .CLK(n8774), .C(n8785) );
  CKBD0 U8702 ( .CLK(n8775), .C(n8786) );
  CKBD0 U8703 ( .CLK(n8776), .C(n8787) );
  CKBD0 U8704 ( .CLK(n8781), .C(n8788) );
  CKBD0 U8705 ( .CLK(n8780), .C(n8789) );
  BUFFD0 U8706 ( .I(n8782), .Z(n8790) );
  CKBD0 U8707 ( .CLK(n8783), .C(n8791) );
  CKBD0 U8708 ( .CLK(n8784), .C(n8792) );
  CKBD0 U8709 ( .CLK(n8785), .C(n8793) );
  CKBD0 U8710 ( .CLK(n8786), .C(n8794) );
  CKBD0 U8711 ( .CLK(n8787), .C(n8795) );
  BUFFD0 U8712 ( .I(n8788), .Z(n8796) );
  CKBD0 U8713 ( .CLK(n8789), .C(n8797) );
  CKBD0 U8714 ( .CLK(n8790), .C(n8798) );
  CKBD0 U8715 ( .CLK(n8791), .C(n8799) );
  CKBD0 U8716 ( .CLK(n8792), .C(n8800) );
  CKBD0 U8717 ( .CLK(n8793), .C(n8801) );
  CKBD0 U8718 ( .CLK(n8667), .C(n8802) );
  BUFFD0 U8719 ( .I(n8669), .Z(n8803) );
  BUFFD0 U8720 ( .I(n8851), .Z(n8804) );
  BUFFD0 U8721 ( .I(n8997), .Z(n8805) );
  BUFFD0 U8722 ( .I(n8852), .Z(n8806) );
  BUFFD0 U8723 ( .I(n8794), .Z(n8807) );
  BUFFD0 U8724 ( .I(n8853), .Z(n8808) );
  BUFFD0 U8725 ( .I(n8573), .Z(n8809) );
  BUFFD0 U8726 ( .I(n8864), .Z(n8810) );
  BUFFD0 U8727 ( .I(n8621), .Z(n8811) );
  BUFFD0 U8728 ( .I(n8721), .Z(n8812) );
  BUFFD0 U8729 ( .I(n8722), .Z(n8813) );
  CKBD0 U8730 ( .CLK(n8795), .C(n8814) );
  CKBD0 U8731 ( .CLK(n8796), .C(n8815) );
  CKBD0 U8732 ( .CLK(n8797), .C(n8816) );
  CKBD0 U8733 ( .CLK(n8798), .C(n8817) );
  CKBD0 U8734 ( .CLK(n8799), .C(n8818) );
  CKBD0 U8735 ( .CLK(n8800), .C(n8819) );
  CKBD0 U8736 ( .CLK(n8801), .C(n8820) );
  CKBD0 U8737 ( .CLK(n8807), .C(n8821) );
  CKBD0 U8738 ( .CLK(n8725), .C(n8822) );
  BUFFD0 U8739 ( .I(n8726), .Z(n8823) );
  CKBD0 U8740 ( .CLK(n8727), .C(n8824) );
  BUFFD0 U8741 ( .I(n8814), .Z(n8825) );
  CKBD0 U8742 ( .CLK(n8815), .C(n8826) );
  CKBD0 U8743 ( .CLK(n8816), .C(n8827) );
  CKBD0 U8744 ( .CLK(n8817), .C(n8828) );
  BUFFD0 U8745 ( .I(n8818), .Z(n8829) );
  BUFFD0 U8746 ( .I(n8732), .Z(n8830) );
  BUFFD0 U8747 ( .I(n8649), .Z(n8831) );
  BUFFD0 U8748 ( .I(n8777), .Z(n8832) );
  CKBD0 U8749 ( .CLK(n8819), .C(n8833) );
  BUFFD0 U8750 ( .I(n8778), .Z(n8834) );
  BUFFD0 U8751 ( .I(n8733), .Z(n8835) );
  CKBD0 U8752 ( .CLK(n8735), .C(n8836) );
  BUFFD0 U8753 ( .I(n8734), .Z(n8837) );
  BUFFD0 U8754 ( .I(n8954), .Z(n8838) );
  BUFFD0 U8755 ( .I(n8744), .Z(n8839) );
  BUFFD0 U8756 ( .I(n8779), .Z(n8840) );
  BUFFD0 U8757 ( .I(n8820), .Z(n8841) );
  BUFFD0 U8758 ( .I(n8802), .Z(n8842) );
  CKBD0 U8759 ( .CLK(n8821), .C(n8843) );
  CKBD0 U8760 ( .CLK(n8825), .C(n8844) );
  CKBD0 U8761 ( .CLK(n8826), .C(n8845) );
  CKBD0 U8762 ( .CLK(n8827), .C(n8846) );
  CKBD0 U8763 ( .CLK(n8828), .C(n8847) );
  CKBD0 U8764 ( .CLK(n8829), .C(n8848) );
  CKBD0 U8765 ( .CLK(n8833), .C(n8849) );
  CKBD0 U8766 ( .CLK(n8803), .C(n8850) );
  BUFFD0 U8767 ( .I(n8958), .Z(n8851) );
  BUFFD0 U8768 ( .I(n8950), .Z(n8852) );
  BUFFD0 U8769 ( .I(n8960), .Z(n8853) );
  CKBD0 U8770 ( .CLK(n8841), .C(n8854) );
  CKBD0 U8771 ( .CLK(n8843), .C(n8855) );
  CKBD0 U8772 ( .CLK(n8844), .C(n8856) );
  CKBD0 U8773 ( .CLK(n8845), .C(n8857) );
  CKBD0 U8774 ( .CLK(n8846), .C(n8858) );
  CKBD0 U8775 ( .CLK(n8847), .C(n8859) );
  CKBD0 U8776 ( .CLK(n8848), .C(n8860) );
  BUFFD0 U8777 ( .I(n8678), .Z(n8861) );
  CKBD0 U8778 ( .CLK(n8809), .C(n8862) );
  CKBD0 U8779 ( .CLK(n8849), .C(n8863) );
  BUFFD0 U8780 ( .I(n8972), .Z(n8864) );
  CKBD0 U8781 ( .CLK(n8811), .C(n8865) );
  CKBD0 U8782 ( .CLK(n8812), .C(n8866) );
  CKBD0 U8783 ( .CLK(n8813), .C(n8867) );
  CKBD0 U8784 ( .CLK(n8854), .C(n8868) );
  CKBD0 U8785 ( .CLK(n8855), .C(n8869) );
  CKBD0 U8786 ( .CLK(n8856), .C(n8870) );
  CKBD0 U8787 ( .CLK(n8857), .C(n8871) );
  CKBD0 U8788 ( .CLK(n8858), .C(n8872) );
  CKBD0 U8789 ( .CLK(n8859), .C(n8873) );
  CKBD0 U8790 ( .CLK(n8860), .C(n8874) );
  CKBD0 U8791 ( .CLK(n8863), .C(n8875) );
  CKBD0 U8792 ( .CLK(n8868), .C(n8876) );
  BUFFD0 U8793 ( .I(n8908), .Z(n8877) );
  CKBD0 U8794 ( .CLK(n8869), .C(n8878) );
  BUFFD0 U8795 ( .I(n8926), .Z(n8879) );
  BUFFD0 U8796 ( .I(n8893), .Z(n8880) );
  BUFFD0 U8797 ( .I(n8872), .Z(n8881) );
  BUFFD0 U8798 ( .I(n8929), .Z(n8882) );
  BUFFD0 U8799 ( .I(n8974), .Z(n8883) );
  BUFFD0 U8800 ( .I(n8875), .Z(n8884) );
  BUFFD0 U8801 ( .I(n8973), .Z(n8885) );
  BUFFD0 U8802 ( .I(n8876), .Z(n8886) );
  CKBD0 U8803 ( .CLK(n8823), .C(n8887) );
  BUFFD0 U8804 ( .I(n8917), .Z(n8888) );
  BUFFD0 U8805 ( .I(n8870), .Z(n8889) );
  CKBD0 U8806 ( .CLK(n8830), .C(n8890) );
  BUFFD0 U8807 ( .I(n8871), .Z(n8891) );
  BUFFD0 U8808 ( .I(n8979), .Z(n8892) );
  BUFFD0 U8809 ( .I(n8918), .Z(n8893) );
  CKBD0 U8810 ( .CLK(n8832), .C(n8894) );
  CKBD0 U8811 ( .CLK(n8834), .C(n8895) );
  CKBD0 U8812 ( .CLK(n8881), .C(n8896) );
  BUFFD0 U8813 ( .I(n8874), .Z(n8897) );
  CKBD0 U8814 ( .CLK(n8884), .C(n8898) );
  CKBD0 U8815 ( .CLK(n8886), .C(n8899) );
  BUFFD0 U8816 ( .I(n8878), .Z(n8900) );
  CKBD0 U8817 ( .CLK(n8889), .C(n8901) );
  CKBD0 U8818 ( .CLK(n8891), .C(n8902) );
  BUFFD0 U8819 ( .I(n8873), .Z(n8903) );
  BUFFD0 U8820 ( .I(n8928), .Z(n8904) );
  CKBD0 U8821 ( .CLK(n8897), .C(n8905) );
  BUFFD0 U8822 ( .I(n8898), .Z(n8906) );
  BUFFD0 U8823 ( .I(n8899), .Z(n8907) );
  BUFFD0 U8824 ( .I(n8916), .Z(n8908) );
  CKBD0 U8825 ( .CLK(n8900), .C(n8909) );
  BUFFD0 U8826 ( .I(n8902), .Z(n8910) );
  CKBD0 U8827 ( .CLK(n8903), .C(n8911) );
  BUFFD0 U8828 ( .I(n8896), .Z(n8912) );
  BUFFD0 U8829 ( .I(n8905), .Z(n8913) );
  CKBD0 U8830 ( .CLK(n8906), .C(n8914) );
  CKBD0 U8831 ( .CLK(n8907), .C(n8915) );
  BUFFD0 U8832 ( .I(n9016), .Z(n8916) );
  BUFFD0 U8833 ( .I(n8924), .Z(n8917) );
  BUFFD0 U8834 ( .I(n9010), .Z(n8918) );
  CKBD0 U8835 ( .CLK(n8910), .C(n8919) );
  CKBD0 U8836 ( .CLK(n8912), .C(n8920) );
  CKBD0 U8837 ( .CLK(n8913), .C(n8921) );
  BUFFD0 U8838 ( .I(n8930), .Z(n8922) );
  BUFFD0 U8839 ( .I(n8915), .Z(n8923) );
  BUFFD0 U8840 ( .I(n9015), .Z(n8924) );
  BUFFD0 U8841 ( .I(n8901), .Z(n8925) );
  BUFFD0 U8842 ( .I(n8966), .Z(n8926) );
  BUFFD0 U8843 ( .I(n8911), .Z(n8927) );
  BUFFD0 U8844 ( .I(n8936), .Z(n8928) );
  BUFFD0 U8845 ( .I(n8938), .Z(n8929) );
  BUFFD0 U8846 ( .I(n9002), .Z(n8930) );
  CKBD0 U8847 ( .CLK(n8923), .C(n8931) );
  BUFFD0 U8848 ( .I(n8909), .Z(n8932) );
  CKBD0 U8849 ( .CLK(n8925), .C(n8933) );
  BUFFD0 U8850 ( .I(n8919), .Z(n8934) );
  CKBD0 U8851 ( .CLK(n8831), .C(n8935) );
  BUFFD0 U8852 ( .I(n9009), .Z(n8936) );
  CKBD0 U8853 ( .CLK(n8927), .C(n8937) );
  BUFFD0 U8854 ( .I(n9011), .Z(n8938) );
  BUFFD0 U8855 ( .I(n8914), .Z(n8939) );
  BUFFD0 U8856 ( .I(n8931), .Z(n8940) );
  CKBD0 U8857 ( .CLK(n8932), .C(n8941) );
  BUFFD0 U8858 ( .I(n8933), .Z(n8942) );
  CKBD0 U8859 ( .CLK(n8934), .C(n8943) );
  BUFFD0 U8860 ( .I(n8920), .Z(n8944) );
  BUFFD0 U8861 ( .I(n8937), .Z(n8945) );
  CKBD0 U8862 ( .CLK(n8839), .C(n8946) );
  CKBD0 U8863 ( .CLK(n8835), .C(n8947) );
  CKBD0 U8864 ( .CLK(n8837), .C(n8948) );
  BUFFD0 U8865 ( .I(n8921), .Z(n8949) );
  BUFFD0 U8866 ( .I(n8992), .Z(n8950) );
  CKBD0 U8867 ( .CLK(n8840), .C(n8951) );
  CKBD0 U8868 ( .CLK(n8842), .C(n8952) );
  CKBD0 U8869 ( .CLK(n8939), .C(n8953) );
  BUFFD0 U8870 ( .I(n8745), .Z(n8954) );
  BUFFD0 U8871 ( .I(n9008), .Z(n8955) );
  BUFFD0 U8872 ( .I(n9007), .Z(n8956) );
  CKBD0 U8873 ( .CLK(n8861), .C(n8957) );
  BUFFD0 U8874 ( .I(n8677), .Z(n8958) );
  BUFFD0 U8875 ( .I(n8850), .Z(n8959) );
  BUFFD0 U8876 ( .I(n8689), .Z(n8960) );
  BUFFD0 U8877 ( .I(n8862), .Z(n8961) );
  BUFFD0 U8878 ( .I(n8866), .Z(n8962) );
  CKBD0 U8879 ( .CLK(n8940), .C(n8963) );
  BUFFD0 U8880 ( .I(n8941), .Z(n8964) );
  CKBD0 U8881 ( .CLK(n8942), .C(n8965) );
  BUFFD0 U8882 ( .I(n9006), .Z(n8966) );
  CKBD0 U8883 ( .CLK(n8944), .C(n8967) );
  CKBD0 U8884 ( .CLK(n8945), .C(n8968) );
  CKBD0 U8885 ( .CLK(n8949), .C(n8969) );
  BUFFD0 U8886 ( .I(n8953), .Z(n8970) );
  BUFFD0 U8887 ( .I(n8990), .Z(n8971) );
  BUFFD0 U8888 ( .I(n8631), .Z(n8972) );
  BUFFD0 U8889 ( .I(n8824), .Z(n8973) );
  BUFFD0 U8890 ( .I(n8822), .Z(n8974) );
  CKBD0 U8891 ( .CLK(n8964), .C(n8975) );
  CKBD0 U8892 ( .CLK(n8965), .C(n8976) );
  BUFFD0 U8893 ( .I(n9012), .Z(n8977) );
  BUFFD0 U8894 ( .I(n8890), .Z(n8978) );
  BUFFD0 U8895 ( .I(n8836), .Z(n8979) );
  BUFFD0 U8896 ( .I(n8894), .Z(n8980) );
  BUFFD0 U8897 ( .I(n8943), .Z(n8981) );
  BUFFD0 U8898 ( .I(n8895), .Z(n8982) );
  BUFFD0 U8899 ( .I(n8967), .Z(n8983) );
  BUFFD0 U8900 ( .I(n8968), .Z(n8984) );
  BUFFD0 U8901 ( .I(n8969), .Z(n8985) );
  CKBD0 U8902 ( .CLK(n8970), .C(n8986) );
  BUFFD0 U8903 ( .I(n8935), .Z(n8987) );
  BUFFD0 U8904 ( .I(n8946), .Z(n8988) );
  BUFFD0 U8905 ( .I(n8947), .Z(n8989) );
  BUFFD0 U8906 ( .I(n9003), .Z(n8990) );
  BUFFD0 U8907 ( .I(n8948), .Z(n8991) );
  BUFFD0 U8908 ( .I(n8680), .Z(n8992) );
  BUFFD0 U8909 ( .I(n8951), .Z(n8993) );
  BUFFD0 U8910 ( .I(n8975), .Z(n8994) );
  BUFFD0 U8911 ( .I(n8976), .Z(n8995) );
  BUFFD0 U8912 ( .I(n8952), .Z(n8996) );
  BUFFD0 U8913 ( .I(n8957), .Z(n8997) );
  CKBD0 U8914 ( .CLK(n8981), .C(n8998) );
  CKBD0 U8915 ( .CLK(n8983), .C(n8999) );
  CKBD0 U8916 ( .CLK(n8984), .C(n9000) );
  CKBD0 U8917 ( .CLK(n8985), .C(n9001) );
  BUFFD0 U8918 ( .I(n9013), .Z(n9002) );
  BUFFD0 U8919 ( .I(n9014), .Z(n9003) );
  CKBD0 U8920 ( .CLK(n8994), .C(n9004) );
  CKBD0 U8921 ( .CLK(n8995), .C(n9005) );
  BUFFD0 U8922 ( .I(n8998), .Z(n9006) );
  BUFFD0 U8923 ( .I(n8865), .Z(n9007) );
  BUFFD0 U8924 ( .I(n8867), .Z(n9008) );
  BUFFD0 U8925 ( .I(n8999), .Z(n9009) );
  BUFFD0 U8926 ( .I(n9000), .Z(n9010) );
  BUFFD0 U8927 ( .I(n9001), .Z(n9011) );
  BUFFD0 U8928 ( .I(n8887), .Z(n9012) );
  BUFFD0 U8929 ( .I(n8986), .Z(n9013) );
  BUFFD0 U8930 ( .I(n8963), .Z(n9014) );
  BUFFD0 U8931 ( .I(n9004), .Z(n9015) );
  BUFFD0 U8932 ( .I(n9005), .Z(n9016) );
  BUFFD0 U8933 ( .I(n9125), .Z(n9017) );
  INR2XD0 U8934 ( .A1(n9026), .B1(n9127), .ZN(n9235) );
  BUFFD0 U8935 ( .I(n9019), .Z(n9018) );
  BUFFD0 U8936 ( .I(n9235), .Z(n9019) );
  CKBD0 U8937 ( .CLK(ParValidTimer[1]), .C(n9020) );
  BUFFD0 U8938 ( .I(n9234), .Z(n9021) );
  BUFFD0 U8939 ( .I(n9023), .Z(n9022) );
  BUFFD0 U8940 ( .I(n9290), .Z(n9023) );
  BUFFD1 U8941 ( .I(n9161), .Z(n9160) );
  BUFFD1 U8942 ( .I(n9161), .Z(n9159) );
  BUFFD1 U8943 ( .I(n9162), .Z(n9158) );
  BUFFD1 U8944 ( .I(n9162), .Z(n9157) );
  BUFFD1 U8945 ( .I(n9163), .Z(n9161) );
  BUFFD1 U8946 ( .I(n9163), .Z(n9162) );
  BUFFD1 U8947 ( .I(n9164), .Z(n9163) );
  INVD1 U8948 ( .I(Reset), .ZN(n9164) );
  INVD1 U8949 ( .I(n9285), .ZN(n9125) );
  BUFFD1 U8950 ( .I(n9130), .Z(n9141) );
  BUFFD1 U8951 ( .I(n9130), .Z(n9142) );
  BUFFD1 U8952 ( .I(n9131), .Z(n9143) );
  BUFFD1 U8953 ( .I(n9131), .Z(n9144) );
  BUFFD1 U8954 ( .I(n9132), .Z(n9145) );
  BUFFD1 U8955 ( .I(n9132), .Z(n9146) );
  BUFFD1 U8956 ( .I(n9133), .Z(n9147) );
  BUFFD1 U8957 ( .I(n9133), .Z(n9148) );
  BUFFD1 U8958 ( .I(n9134), .Z(n9149) );
  BUFFD1 U8959 ( .I(n9134), .Z(n9150) );
  BUFFD1 U8960 ( .I(n9135), .Z(n9151) );
  BUFFD1 U8961 ( .I(n9135), .Z(n9152) );
  BUFFD1 U8962 ( .I(n9136), .Z(n9153) );
  BUFFD1 U8963 ( .I(n9136), .Z(n9154) );
  BUFFD1 U8964 ( .I(n9137), .Z(n9155) );
  BUFFD1 U8965 ( .I(n9137), .Z(n9156) );
  INVD1 U8966 ( .I(n9166), .ZN(n9127) );
  INVD1 U8967 ( .I(n9166), .ZN(n9128) );
  INVD1 U8968 ( .I(n9166), .ZN(n9129) );
  BUFFD1 U8969 ( .I(n9285), .Z(n9126) );
  BUFFD1 U8970 ( .I(n9139), .Z(n9132) );
  BUFFD1 U8971 ( .I(n9139), .Z(n9133) );
  BUFFD1 U8972 ( .I(n9139), .Z(n9134) );
  BUFFD1 U8973 ( .I(n9138), .Z(n9135) );
  BUFFD1 U8974 ( .I(n9138), .Z(n9136) );
  BUFFD1 U8975 ( .I(n9138), .Z(n9137) );
  BUFFD1 U8976 ( .I(n9140), .Z(n9130) );
  BUFFD1 U8977 ( .I(n9140), .Z(n9131) );
  IND2D1 U8978 ( .A1(n9284), .B1(n9283), .ZN(n9285) );
  BUFFD1 U8979 ( .I(SerClock), .Z(n9139) );
  BUFFD1 U8980 ( .I(SerClock), .Z(n9138) );
  BUFFD1 U8981 ( .I(SerClock), .Z(n9140) );
  NR2D1 U8982 ( .A1(ParClk), .A2(n9165), .ZN(n9293) );
  NR2D1 U8983 ( .A1(ParClk), .A2(n9271), .ZN(N37) );
  NR4D0 U8984 ( .A1(n9270), .A2(Count32[2]), .A3(Count32[4]), .A4(Count32[3]), 
        .ZN(n9272) );
  AN2D1 U8985 ( .A1(N34), .A2(n9294), .Z(N42) );
  AN2D1 U8986 ( .A1(N33), .A2(n9294), .Z(N41) );
  AN2D1 U8987 ( .A1(N32), .A2(n9294), .Z(N40) );
  AN2D1 U8988 ( .A1(N31), .A2(n9294), .Z(N39) );
  INVD1 U8989 ( .I(n9020), .ZN(n9291) );
  AO22D0 U8990 ( .A1(n6965), .A2(n9017), .B1(n6830), .B2(n9285), .Z(n9199) );
  AO22D0 U8991 ( .A1(n6828), .A2(n9017), .B1(n6693), .B2(n9285), .Z(n9198) );
  AO22D0 U8992 ( .A1(n6691), .A2(n9017), .B1(n6556), .B2(n9285), .Z(n9197) );
  AO22D0 U8993 ( .A1(n6554), .A2(n9017), .B1(n6419), .B2(n9285), .Z(n9196) );
  AO22D0 U8994 ( .A1(n6417), .A2(n9017), .B1(n6282), .B2(n9285), .Z(n9195) );
  AO22D0 U8995 ( .A1(n6280), .A2(n9017), .B1(n6145), .B2(n9285), .Z(n9194) );
  AO22D0 U8996 ( .A1(n6006), .A2(n9017), .B1(Decoder[7]), .B2(n9285), .Z(n9192) );
  AO22D0 U8997 ( .A1(n5870), .A2(n9125), .B1(Decoder[8]), .B2(n9126), .Z(n9191) );
  AO22D0 U8998 ( .A1(n5734), .A2(n9125), .B1(Decoder[9]), .B2(n9126), .Z(n9190) );
  AO22D0 U8999 ( .A1(n5598), .A2(n9125), .B1(Decoder[10]), .B2(n9126), .Z(
        n9189) );
  AO22D0 U9000 ( .A1(n5462), .A2(n9017), .B1(Decoder[11]), .B2(n9126), .Z(
        n9188) );
  AO22D0 U9001 ( .A1(n5326), .A2(n9125), .B1(n5190), .B2(n9126), .Z(n9187) );
  AO22D0 U9002 ( .A1(n5189), .A2(n9125), .B1(Decoder[13]), .B2(n9126), .Z(
        n9186) );
  AO22D0 U9003 ( .A1(n5053), .A2(n9125), .B1(Decoder[14]), .B2(n9126), .Z(
        n9185) );
  AO22D0 U9004 ( .A1(n4917), .A2(n9125), .B1(Decoder[15]), .B2(n9126), .Z(
        n9184) );
  AO22D0 U9005 ( .A1(n4781), .A2(n9125), .B1(Decoder[16]), .B2(n9126), .Z(
        n9183) );
  AO22D0 U9006 ( .A1(n4645), .A2(n9125), .B1(Decoder[17]), .B2(n9126), .Z(
        n9182) );
  AO22D0 U9007 ( .A1(n4509), .A2(n9125), .B1(Decoder[18]), .B2(n9126), .Z(
        n9181) );
  AO22D0 U9008 ( .A1(n4373), .A2(n9125), .B1(Decoder[19]), .B2(n9126), .Z(
        n9180) );
  AO22D0 U9009 ( .A1(n4236), .A2(n9125), .B1(Decoder[20]), .B2(n9126), .Z(
        n9179) );
  AO22D0 U9010 ( .A1(n4100), .A2(n9125), .B1(Decoder[21]), .B2(n9126), .Z(
        n9178) );
  AO22D0 U9011 ( .A1(n3964), .A2(n9017), .B1(Decoder[22]), .B2(n9126), .Z(
        n9177) );
  AO22D0 U9012 ( .A1(n3828), .A2(n9017), .B1(Decoder[23]), .B2(n9126), .Z(
        n9176) );
  AO22D0 U9013 ( .A1(n3692), .A2(n9017), .B1(Decoder[24]), .B2(n9285), .Z(
        n9175) );
  AO22D0 U9014 ( .A1(n3556), .A2(n9017), .B1(Decoder[25]), .B2(n9285), .Z(
        n9174) );
  AO22D0 U9015 ( .A1(n3420), .A2(n9125), .B1(Decoder[26]), .B2(n9126), .Z(
        n9173) );
  AO22D0 U9016 ( .A1(n3284), .A2(n9125), .B1(Decoder[27]), .B2(n9285), .Z(
        n9172) );
  AO22D0 U9017 ( .A1(n3148), .A2(n9125), .B1(Decoder[28]), .B2(n9126), .Z(
        n9171) );
  AO22D0 U9018 ( .A1(n3012), .A2(n9125), .B1(Decoder[29]), .B2(n9285), .Z(
        n9170) );
  AO22D0 U9019 ( .A1(n2876), .A2(n9125), .B1(Decoder[30]), .B2(n9285), .Z(
        n9169) );
  AO22D0 U9020 ( .A1(n2737), .A2(n9125), .B1(Decoder[31]), .B2(n9126), .Z(
        n9168) );
  OAI31D0 U9021 ( .A1(n9292), .A2(n9167), .A3(n9291), .B(n9165), .ZN(n9026) );
  NR2D1 U9022 ( .A1(n9287), .A2(n9127), .ZN(n9233) );
  NR2D1 U9023 ( .A1(n6971), .A2(n9127), .ZN(n9232) );
  NR2D1 U9024 ( .A1(n9127), .A2(n9022), .ZN(n9234) );
  XOR2D1 U9025 ( .A1(n9167), .A2(n9289), .Z(n9290) );
  NR2D1 U9026 ( .A1(n9291), .A2(n9288), .ZN(n9289) );
  NR4D0 U9027 ( .A1(n9276), .A2(n8996), .A3(n8140), .A4(n8330), .ZN(n9277) );
  ND2D1 U9028 ( .A1(n9282), .A2(n9281), .ZN(n9284) );
  NR4D0 U9029 ( .A1(n8888), .A2(n8922), .A3(n8904), .A4(n8879), .ZN(n9282) );
  NR4D0 U9030 ( .A1(n8877), .A2(n8971), .A3(n8882), .A4(n8880), .ZN(n9281) );
  AN4D1 U9031 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .Z(n9283) );
  INR4D0 U9032 ( .A1(n8172), .B1(n9273), .B2(n8417), .B3(n8223), .ZN(n9280) );
  NR4D0 U9033 ( .A1(n9274), .A2(n8415), .A3(n8197), .A4(n8182), .ZN(n9279) );
  NR4D0 U9034 ( .A1(n9275), .A2(n8266), .A3(n8335), .A4(n8444), .ZN(n9278) );
  ND3D1 U9035 ( .A1(n8234), .A2(n8892), .A3(n8224), .ZN(n9273) );
  AN2D1 U9036 ( .A1(SerClk), .A2(SerValid), .Z(SerClock) );
endmodule


module SerialRx_1 ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;
  wire   n2;

  PLLTop_1 PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid3_1 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [2:0] ReadAddr;
  output [2:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n927, n928, n929, StateClockRaw, StateClock, N46, N47, N48, N49, N63,
         N64, N65, N66, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n53, n70, n71, n91, n114, n116,
         n117, n118, n119, n120, n123, n125, n126, n139, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [2:0] OldReadAr;
  wire   [2:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n13), .CPN(StateClock), .Q(FullFIFO), .QN(n851) );
  DFND1 EmptyFIFOr_reg ( .D(n847), .CPN(StateClock), .Q(n927) );
  IAO21D1 U6 ( .A1(n922), .A2(n921), .B(Reset), .ZN(n923) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n120), .CPN(StateClock), .CDN(n829), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n171), .CPN(StateClock), .CDN(n829), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n174), .CPN(StateClock), .CDN(n829), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n176), .CPN(StateClock), .CDN(n829), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n178), .CPN(StateClock), .CDN(n829), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n209), .CPN(StateClock), .CDN(n829), .Q(
        OldReadAr[1]) );
  DFNCND1 ReadCmdr_reg ( .D(n239), .CPN(StateClock), .CDN(n829), .Q(n928), 
        .QN(n6) );
  DFNCND1 WriteCmdr_reg ( .D(n288), .CPN(StateClock), .CDN(n829), .Q(n929) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n830), 
        .Q(CurState[2]), .QN(n894) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n830), 
        .Q(CurState[1]), .QN(n910) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n830), 
        .Q(CurState[0]), .QN(n885) );
  EDFCND1 \WriteAr_reg[2]  ( .D(n468), .E(n3), .CP(StateClock), .CDN(n830), 
        .Q(WriteAddr[2]), .QN(n917) );
  EDFCND1 \WriteAr_reg[1]  ( .D(n500), .E(n3), .CP(StateClock), .CDN(n830), 
        .Q(WriteAddr[1]), .QN(n918) );
  EDFCND1 \ReadAr_reg[2]  ( .D(n533), .E(n627), .CP(StateClock), .CDN(n830), 
        .Q(ReadAddr[2]), .QN(n834) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n567), .E(n627), .CP(StateClock), .CDN(n830), 
        .Q(ReadAddr[1]), .QN(n833) );
  EDFCND1 \ReadAr_reg[0]  ( .D(n597), .E(n627), .CP(StateClock), .CDN(n830), 
        .Q(ReadAddr[0]), .QN(n832) );
  EDFCND1 \WriteAr_reg[0]  ( .D(n650), .E(n3), .CP(StateClock), .CDN(n830), 
        .Q(WriteAddr[0]), .QN(n831) );
  DFNCND1 \NextState_reg[1]  ( .D(n713), .CPN(StateClock), .CDN(n830), .Q(
        NextState[1]), .QN(n849) );
  DFNCND1 \NextState_reg[0]  ( .D(n749), .CPN(StateClock), .CDN(n830), .Q(
        NextState[0]), .QN(n848) );
  DFNCND1 \NextState_reg[2]  ( .D(n785), .CPN(StateClock), .CDN(n830), .Q(
        NextState[2]), .QN(n850) );
  CKBD0 U3 ( .CLK(n465), .C(n466) );
  INVD0 U4 ( .I(n921), .ZN(n926) );
  BUFFD0 U5 ( .I(n710), .Z(n1) );
  BUFFD0 U7 ( .I(n628), .Z(n2) );
  BUFFD0 U8 ( .I(n685), .Z(n3) );
  AN3D1 U9 ( .A1(n699), .A2(n710), .A3(n853), .Z(n4) );
  INVD1 U10 ( .I(n4), .ZN(N66) );
  AN2D1 U11 ( .A1(n6), .A2(n2), .Z(n5) );
  INVD1 U12 ( .I(n5), .ZN(N48) );
  CKBD0 U13 ( .CLK(n927), .C(n463) );
  BUFFD0 U14 ( .I(n8), .Z(n7) );
  BUFFD0 U15 ( .I(n9), .Z(n8) );
  BUFFD0 U16 ( .I(n10), .Z(n9) );
  BUFFD0 U17 ( .I(n11), .Z(n10) );
  BUFFD0 U18 ( .I(n12), .Z(n11) );
  BUFFD0 U19 ( .I(n851), .Z(n12) );
  BUFFD0 U20 ( .I(n14), .Z(n13) );
  BUFFD0 U21 ( .I(n15), .Z(n14) );
  BUFFD0 U22 ( .I(n16), .Z(n15) );
  BUFFD0 U23 ( .I(n17), .Z(n16) );
  BUFFD0 U24 ( .I(n18), .Z(n17) );
  BUFFD0 U25 ( .I(n19), .Z(n18) );
  BUFFD0 U26 ( .I(n20), .Z(n19) );
  BUFFD0 U27 ( .I(n21), .Z(n20) );
  BUFFD0 U28 ( .I(n22), .Z(n21) );
  BUFFD0 U29 ( .I(n23), .Z(n22) );
  BUFFD0 U30 ( .I(n24), .Z(n23) );
  BUFFD0 U31 ( .I(n25), .Z(n24) );
  BUFFD0 U32 ( .I(n26), .Z(n25) );
  BUFFD0 U33 ( .I(n27), .Z(n26) );
  BUFFD0 U34 ( .I(n28), .Z(n27) );
  BUFFD0 U35 ( .I(n29), .Z(n28) );
  BUFFD0 U36 ( .I(n30), .Z(n29) );
  BUFFD0 U37 ( .I(n31), .Z(n30) );
  BUFFD0 U38 ( .I(n32), .Z(n31) );
  BUFFD0 U39 ( .I(n33), .Z(n32) );
  BUFFD0 U40 ( .I(n34), .Z(n33) );
  BUFFD0 U41 ( .I(n53), .Z(n34) );
  BUFFD0 U42 ( .I(n70), .Z(n53) );
  BUFFD0 U43 ( .I(n71), .Z(n70) );
  BUFFD0 U44 ( .I(n91), .Z(n71) );
  BUFFD0 U45 ( .I(n114), .Z(n91) );
  BUFFD0 U46 ( .I(n116), .Z(n114) );
  BUFFD0 U47 ( .I(n117), .Z(n116) );
  BUFFD0 U48 ( .I(n118), .Z(n117) );
  BUFFD0 U49 ( .I(n119), .Z(n118) );
  BUFFD0 U50 ( .I(n846), .Z(n119) );
  MOAI22D0 U51 ( .A1(n832), .A2(n920), .B1(n920), .B2(n165), .ZN(n835) );
  BUFFD0 U52 ( .I(n123), .Z(n120) );
  BUFFD0 U53 ( .I(n125), .Z(n123) );
  BUFFD0 U54 ( .I(n126), .Z(n125) );
  BUFFD0 U55 ( .I(n139), .Z(n126) );
  BUFFD0 U56 ( .I(n145), .Z(n139) );
  BUFFD0 U57 ( .I(n146), .Z(n145) );
  BUFFD0 U58 ( .I(n147), .Z(n146) );
  BUFFD0 U59 ( .I(n148), .Z(n147) );
  BUFFD0 U60 ( .I(n149), .Z(n148) );
  BUFFD0 U61 ( .I(n150), .Z(n149) );
  BUFFD0 U62 ( .I(n151), .Z(n150) );
  BUFFD0 U63 ( .I(n152), .Z(n151) );
  BUFFD0 U64 ( .I(n153), .Z(n152) );
  BUFFD0 U65 ( .I(n154), .Z(n153) );
  BUFFD0 U66 ( .I(n155), .Z(n154) );
  BUFFD0 U67 ( .I(n156), .Z(n155) );
  BUFFD0 U68 ( .I(n157), .Z(n156) );
  BUFFD0 U69 ( .I(n158), .Z(n157) );
  BUFFD0 U70 ( .I(n159), .Z(n158) );
  BUFFD0 U71 ( .I(n160), .Z(n159) );
  BUFFD0 U72 ( .I(n161), .Z(n160) );
  BUFFD0 U73 ( .I(n162), .Z(n161) );
  BUFFD0 U74 ( .I(n163), .Z(n162) );
  BUFFD0 U75 ( .I(n164), .Z(n163) );
  BUFFD0 U76 ( .I(n167), .Z(n164) );
  BUFFD0 U77 ( .I(n166), .Z(n165) );
  BUFFD0 U78 ( .I(n168), .Z(n166) );
  BUFFD0 U79 ( .I(n169), .Z(n167) );
  BUFFD0 U80 ( .I(n170), .Z(n168) );
  BUFFD0 U81 ( .I(n835), .Z(n169) );
  BUFFD0 U82 ( .I(n270), .Z(n170) );
  MOAI22D0 U83 ( .A1(n831), .A2(n919), .B1(n919), .B2(n173), .ZN(n841) );
  BUFFD0 U84 ( .I(n172), .Z(n171) );
  BUFFD0 U85 ( .I(n841), .Z(n172) );
  BUFFD0 U86 ( .I(n292), .Z(n173) );
  MOAI22D0 U87 ( .A1(n919), .A2(n917), .B1(n919), .B2(n175), .ZN(n842) );
  BUFFD0 U88 ( .I(n842), .Z(n174) );
  BUFFD0 U89 ( .I(n291), .Z(n175) );
  MOAI22D0 U90 ( .A1(n919), .A2(n918), .B1(n919), .B2(n177), .ZN(n843) );
  BUFFD0 U91 ( .I(n843), .Z(n176) );
  BUFFD0 U92 ( .I(n290), .Z(n177) );
  MOAI22D0 U93 ( .A1(n834), .A2(n920), .B1(n920), .B2(n203), .ZN(n844) );
  BUFFD0 U94 ( .I(n179), .Z(n178) );
  BUFFD0 U95 ( .I(n180), .Z(n179) );
  BUFFD0 U96 ( .I(n181), .Z(n180) );
  BUFFD0 U97 ( .I(n182), .Z(n181) );
  BUFFD0 U98 ( .I(n183), .Z(n182) );
  BUFFD0 U99 ( .I(n184), .Z(n183) );
  BUFFD0 U100 ( .I(n185), .Z(n184) );
  BUFFD0 U101 ( .I(n186), .Z(n185) );
  BUFFD0 U102 ( .I(n187), .Z(n186) );
  BUFFD0 U103 ( .I(n188), .Z(n187) );
  BUFFD0 U104 ( .I(n189), .Z(n188) );
  BUFFD0 U105 ( .I(n190), .Z(n189) );
  BUFFD0 U106 ( .I(n191), .Z(n190) );
  BUFFD0 U107 ( .I(n192), .Z(n191) );
  BUFFD0 U108 ( .I(n193), .Z(n192) );
  BUFFD0 U109 ( .I(n194), .Z(n193) );
  BUFFD0 U110 ( .I(n195), .Z(n194) );
  BUFFD0 U111 ( .I(n196), .Z(n195) );
  BUFFD0 U112 ( .I(n197), .Z(n196) );
  BUFFD0 U113 ( .I(n198), .Z(n197) );
  BUFFD0 U114 ( .I(n199), .Z(n198) );
  BUFFD0 U115 ( .I(n200), .Z(n199) );
  BUFFD0 U116 ( .I(n201), .Z(n200) );
  BUFFD0 U117 ( .I(n202), .Z(n201) );
  BUFFD0 U118 ( .I(n205), .Z(n202) );
  BUFFD0 U119 ( .I(n204), .Z(n203) );
  BUFFD0 U120 ( .I(n206), .Z(n204) );
  BUFFD0 U121 ( .I(n207), .Z(n205) );
  BUFFD0 U122 ( .I(n208), .Z(n206) );
  BUFFD0 U123 ( .I(n844), .Z(n207) );
  BUFFD0 U124 ( .I(n271), .Z(n208) );
  MOAI22D0 U125 ( .A1(n833), .A2(n920), .B1(n920), .B2(n234), .ZN(n845) );
  BUFFD0 U126 ( .I(n210), .Z(n209) );
  BUFFD0 U127 ( .I(n211), .Z(n210) );
  BUFFD0 U128 ( .I(n212), .Z(n211) );
  BUFFD0 U129 ( .I(n213), .Z(n212) );
  BUFFD0 U130 ( .I(n214), .Z(n213) );
  BUFFD0 U131 ( .I(n215), .Z(n214) );
  BUFFD0 U132 ( .I(n216), .Z(n215) );
  BUFFD0 U133 ( .I(n217), .Z(n216) );
  BUFFD0 U134 ( .I(n218), .Z(n217) );
  BUFFD0 U135 ( .I(n219), .Z(n218) );
  BUFFD0 U136 ( .I(n220), .Z(n219) );
  BUFFD0 U137 ( .I(n221), .Z(n220) );
  BUFFD0 U138 ( .I(n222), .Z(n221) );
  BUFFD0 U139 ( .I(n223), .Z(n222) );
  BUFFD0 U140 ( .I(n224), .Z(n223) );
  BUFFD0 U141 ( .I(n225), .Z(n224) );
  BUFFD0 U142 ( .I(n226), .Z(n225) );
  BUFFD0 U143 ( .I(n227), .Z(n226) );
  BUFFD0 U144 ( .I(n228), .Z(n227) );
  BUFFD0 U145 ( .I(n229), .Z(n228) );
  BUFFD0 U146 ( .I(n230), .Z(n229) );
  BUFFD0 U147 ( .I(n231), .Z(n230) );
  BUFFD0 U148 ( .I(n232), .Z(n231) );
  BUFFD0 U149 ( .I(n233), .Z(n232) );
  BUFFD0 U150 ( .I(n235), .Z(n233) );
  BUFFD0 U151 ( .I(n236), .Z(n234) );
  BUFFD0 U152 ( .I(n237), .Z(n235) );
  BUFFD0 U153 ( .I(n238), .Z(n236) );
  BUFFD0 U154 ( .I(n845), .Z(n237) );
  BUFFD0 U155 ( .I(n269), .Z(n238) );
  BUFFD0 U156 ( .I(n240), .Z(n239) );
  BUFFD0 U157 ( .I(n241), .Z(n240) );
  BUFFD0 U158 ( .I(n242), .Z(n241) );
  BUFFD0 U159 ( .I(n243), .Z(n242) );
  BUFFD0 U160 ( .I(n244), .Z(n243) );
  BUFFD0 U161 ( .I(n245), .Z(n244) );
  BUFFD0 U162 ( .I(n246), .Z(n245) );
  BUFFD0 U163 ( .I(n247), .Z(n246) );
  BUFFD0 U164 ( .I(n248), .Z(n247) );
  BUFFD0 U165 ( .I(n249), .Z(n248) );
  BUFFD0 U166 ( .I(n250), .Z(n249) );
  BUFFD0 U167 ( .I(n251), .Z(n250) );
  BUFFD0 U168 ( .I(n252), .Z(n251) );
  BUFFD0 U169 ( .I(n253), .Z(n252) );
  BUFFD0 U170 ( .I(n254), .Z(n253) );
  BUFFD0 U171 ( .I(n255), .Z(n254) );
  BUFFD0 U172 ( .I(n256), .Z(n255) );
  BUFFD0 U173 ( .I(n257), .Z(n256) );
  BUFFD0 U174 ( .I(n258), .Z(n257) );
  BUFFD0 U175 ( .I(n259), .Z(n258) );
  BUFFD0 U176 ( .I(n260), .Z(n259) );
  BUFFD0 U177 ( .I(n261), .Z(n260) );
  BUFFD0 U178 ( .I(n262), .Z(n261) );
  BUFFD0 U179 ( .I(n263), .Z(n262) );
  BUFFD0 U180 ( .I(n264), .Z(n263) );
  BUFFD0 U181 ( .I(n265), .Z(n264) );
  BUFFD0 U182 ( .I(n266), .Z(n265) );
  BUFFD0 U183 ( .I(n267), .Z(n266) );
  BUFFD0 U184 ( .I(n268), .Z(n267) );
  BUFFD0 U185 ( .I(n836), .Z(n268) );
  BUFFD0 U186 ( .I(n272), .Z(n269) );
  BUFFD0 U187 ( .I(n273), .Z(n270) );
  BUFFD0 U188 ( .I(n274), .Z(n271) );
  CKND2D0 U189 ( .A1(ReadCmd), .A2(n2), .ZN(n856) );
  BUFFD0 U190 ( .I(n275), .Z(n272) );
  BUFFD0 U191 ( .I(n276), .Z(n273) );
  BUFFD0 U192 ( .I(n277), .Z(n274) );
  BUFFD0 U193 ( .I(n278), .Z(n275) );
  BUFFD0 U194 ( .I(n279), .Z(n276) );
  BUFFD0 U195 ( .I(n280), .Z(n277) );
  BUFFD0 U196 ( .I(n281), .Z(n278) );
  BUFFD0 U197 ( .I(n282), .Z(n279) );
  BUFFD0 U198 ( .I(n283), .Z(n280) );
  BUFFD0 U199 ( .I(n284), .Z(n281) );
  BUFFD0 U200 ( .I(n285), .Z(n282) );
  BUFFD0 U201 ( .I(n286), .Z(n283) );
  BUFFD0 U202 ( .I(n287), .Z(n284) );
  BUFFD0 U203 ( .I(OldReadAr[0]), .Z(n285) );
  BUFFD0 U204 ( .I(OldReadAr[2]), .Z(n286) );
  BUFFD0 U205 ( .I(OldReadAr[1]), .Z(n287) );
  BUFFD0 U206 ( .I(n289), .Z(n288) );
  BUFFD0 U207 ( .I(n838), .Z(n289) );
  BUFFD0 U208 ( .I(n294), .Z(n290) );
  BUFFD0 U209 ( .I(n295), .Z(n291) );
  BUFFD0 U210 ( .I(n296), .Z(n292) );
  BUFFD0 U211 ( .I(n929), .Z(n293) );
  BUFFD0 U212 ( .I(n298), .Z(n294) );
  BUFFD0 U213 ( .I(n299), .Z(n295) );
  BUFFD0 U214 ( .I(n300), .Z(n296) );
  BUFFD0 U215 ( .I(n293), .Z(n297) );
  BUFFD0 U216 ( .I(n302), .Z(n298) );
  BUFFD0 U217 ( .I(n303), .Z(n299) );
  BUFFD0 U218 ( .I(n304), .Z(n300) );
  BUFFD0 U219 ( .I(n297), .Z(n301) );
  BUFFD0 U220 ( .I(n306), .Z(n302) );
  BUFFD0 U221 ( .I(n307), .Z(n303) );
  BUFFD0 U222 ( .I(n308), .Z(n304) );
  BUFFD0 U223 ( .I(n301), .Z(n305) );
  BUFFD0 U224 ( .I(n310), .Z(n306) );
  BUFFD0 U225 ( .I(n311), .Z(n307) );
  BUFFD0 U226 ( .I(n312), .Z(n308) );
  BUFFD0 U227 ( .I(n305), .Z(n309) );
  BUFFD0 U228 ( .I(n314), .Z(n310) );
  BUFFD0 U229 ( .I(n315), .Z(n311) );
  BUFFD0 U230 ( .I(n316), .Z(n312) );
  BUFFD0 U231 ( .I(n309), .Z(n313) );
  BUFFD0 U232 ( .I(n318), .Z(n314) );
  BUFFD0 U233 ( .I(n319), .Z(n315) );
  BUFFD0 U234 ( .I(n320), .Z(n316) );
  BUFFD0 U235 ( .I(n313), .Z(n317) );
  BUFFD0 U236 ( .I(n322), .Z(n318) );
  BUFFD0 U237 ( .I(n323), .Z(n319) );
  BUFFD0 U238 ( .I(n324), .Z(n320) );
  BUFFD0 U239 ( .I(n317), .Z(n321) );
  BUFFD0 U240 ( .I(n326), .Z(n322) );
  BUFFD0 U241 ( .I(n327), .Z(n323) );
  BUFFD0 U242 ( .I(n328), .Z(n324) );
  BUFFD0 U243 ( .I(n321), .Z(n325) );
  BUFFD0 U244 ( .I(n330), .Z(n326) );
  BUFFD0 U245 ( .I(n331), .Z(n327) );
  BUFFD0 U246 ( .I(n332), .Z(n328) );
  BUFFD0 U247 ( .I(n325), .Z(n329) );
  BUFFD0 U248 ( .I(n334), .Z(n330) );
  BUFFD0 U249 ( .I(n335), .Z(n331) );
  BUFFD0 U250 ( .I(n336), .Z(n332) );
  BUFFD0 U251 ( .I(n329), .Z(n333) );
  BUFFD0 U252 ( .I(n338), .Z(n334) );
  BUFFD0 U253 ( .I(n339), .Z(n335) );
  BUFFD0 U254 ( .I(n340), .Z(n336) );
  BUFFD0 U255 ( .I(n333), .Z(n337) );
  BUFFD0 U256 ( .I(n342), .Z(n338) );
  BUFFD0 U257 ( .I(n343), .Z(n339) );
  BUFFD0 U258 ( .I(n344), .Z(n340) );
  BUFFD0 U259 ( .I(n337), .Z(n341) );
  BUFFD0 U260 ( .I(n346), .Z(n342) );
  BUFFD0 U261 ( .I(n347), .Z(n343) );
  BUFFD0 U262 ( .I(n348), .Z(n344) );
  BUFFD0 U263 ( .I(n341), .Z(n345) );
  BUFFD0 U264 ( .I(n350), .Z(n346) );
  BUFFD0 U265 ( .I(n351), .Z(n347) );
  BUFFD0 U266 ( .I(n352), .Z(n348) );
  BUFFD0 U267 ( .I(n345), .Z(n349) );
  BUFFD0 U268 ( .I(n354), .Z(n350) );
  BUFFD0 U269 ( .I(n355), .Z(n351) );
  BUFFD0 U270 ( .I(n356), .Z(n352) );
  BUFFD0 U271 ( .I(n349), .Z(n353) );
  BUFFD0 U272 ( .I(n358), .Z(n354) );
  BUFFD0 U273 ( .I(n359), .Z(n355) );
  BUFFD0 U274 ( .I(n360), .Z(n356) );
  BUFFD0 U275 ( .I(n353), .Z(n357) );
  BUFFD0 U276 ( .I(n362), .Z(n358) );
  BUFFD0 U277 ( .I(n363), .Z(n359) );
  BUFFD0 U278 ( .I(n364), .Z(n360) );
  BUFFD0 U279 ( .I(n357), .Z(n361) );
  BUFFD0 U280 ( .I(n366), .Z(n362) );
  BUFFD0 U281 ( .I(n367), .Z(n363) );
  BUFFD0 U282 ( .I(n368), .Z(n364) );
  BUFFD0 U283 ( .I(n361), .Z(n365) );
  BUFFD0 U284 ( .I(n370), .Z(n366) );
  BUFFD0 U285 ( .I(n371), .Z(n367) );
  BUFFD0 U286 ( .I(n372), .Z(n368) );
  BUFFD0 U287 ( .I(n365), .Z(n369) );
  BUFFD0 U288 ( .I(n374), .Z(n370) );
  BUFFD0 U289 ( .I(n375), .Z(n371) );
  BUFFD0 U290 ( .I(n376), .Z(n372) );
  BUFFD0 U291 ( .I(n369), .Z(n373) );
  BUFFD0 U292 ( .I(n378), .Z(n374) );
  BUFFD0 U293 ( .I(n379), .Z(n375) );
  BUFFD0 U294 ( .I(n380), .Z(n376) );
  BUFFD0 U295 ( .I(n373), .Z(n377) );
  BUFFD0 U296 ( .I(n382), .Z(n378) );
  BUFFD0 U297 ( .I(n383), .Z(n379) );
  BUFFD0 U298 ( .I(n384), .Z(n380) );
  BUFFD0 U299 ( .I(n377), .Z(n381) );
  BUFFD0 U300 ( .I(n386), .Z(n382) );
  BUFFD0 U301 ( .I(n387), .Z(n383) );
  BUFFD0 U302 ( .I(n388), .Z(n384) );
  BUFFD0 U303 ( .I(n381), .Z(n385) );
  BUFFD0 U304 ( .I(n390), .Z(n386) );
  BUFFD0 U305 ( .I(n391), .Z(n387) );
  BUFFD0 U306 ( .I(n392), .Z(n388) );
  BUFFD0 U307 ( .I(n385), .Z(n389) );
  BUFFD0 U308 ( .I(n394), .Z(n390) );
  BUFFD0 U309 ( .I(n395), .Z(n391) );
  BUFFD0 U310 ( .I(n396), .Z(n392) );
  BUFFD0 U311 ( .I(n389), .Z(n393) );
  BUFFD0 U312 ( .I(n398), .Z(n394) );
  BUFFD0 U313 ( .I(n399), .Z(n395) );
  BUFFD0 U314 ( .I(n400), .Z(n396) );
  BUFFD0 U315 ( .I(n393), .Z(n397) );
  BUFFD0 U316 ( .I(n402), .Z(n398) );
  BUFFD0 U317 ( .I(n403), .Z(n399) );
  BUFFD0 U318 ( .I(n404), .Z(n400) );
  BUFFD0 U319 ( .I(n397), .Z(n401) );
  BUFFD0 U320 ( .I(n406), .Z(n402) );
  BUFFD0 U321 ( .I(n407), .Z(n403) );
  BUFFD0 U322 ( .I(n408), .Z(n404) );
  BUFFD0 U323 ( .I(n401), .Z(n405) );
  BUFFD0 U324 ( .I(n410), .Z(n406) );
  BUFFD0 U325 ( .I(n411), .Z(n407) );
  BUFFD0 U326 ( .I(n412), .Z(n408) );
  BUFFD0 U327 ( .I(n405), .Z(n409) );
  BUFFD0 U328 ( .I(n414), .Z(n410) );
  BUFFD0 U329 ( .I(n415), .Z(n411) );
  BUFFD0 U330 ( .I(n416), .Z(n412) );
  BUFFD0 U331 ( .I(n409), .Z(n413) );
  BUFFD0 U332 ( .I(n418), .Z(n414) );
  BUFFD0 U333 ( .I(n419), .Z(n415) );
  BUFFD0 U334 ( .I(n420), .Z(n416) );
  BUFFD0 U335 ( .I(n413), .Z(n417) );
  BUFFD0 U336 ( .I(n422), .Z(n418) );
  BUFFD0 U337 ( .I(n423), .Z(n419) );
  BUFFD0 U338 ( .I(n424), .Z(n420) );
  BUFFD0 U339 ( .I(n417), .Z(n421) );
  BUFFD0 U340 ( .I(n425), .Z(n422) );
  BUFFD0 U341 ( .I(n426), .Z(n423) );
  BUFFD0 U342 ( .I(OldWriteAr[0]), .Z(n424) );
  BUFFD0 U343 ( .I(OldWriteAr[1]), .Z(n425) );
  BUFFD0 U344 ( .I(OldWriteAr[2]), .Z(n426) );
  CKBD0 U345 ( .CLK(n421), .C(WriteCmd) );
  BUFFD0 U346 ( .I(n429), .Z(EmptyFIFO) );
  BUFFD0 U347 ( .I(n430), .Z(n429) );
  BUFFD0 U348 ( .I(n431), .Z(n430) );
  BUFFD0 U349 ( .I(n432), .Z(n431) );
  BUFFD0 U350 ( .I(n433), .Z(n432) );
  BUFFD0 U351 ( .I(n434), .Z(n433) );
  BUFFD0 U352 ( .I(n435), .Z(n434) );
  BUFFD0 U353 ( .I(n436), .Z(n435) );
  BUFFD0 U354 ( .I(n437), .Z(n436) );
  BUFFD0 U355 ( .I(n438), .Z(n437) );
  BUFFD0 U356 ( .I(n439), .Z(n438) );
  BUFFD0 U357 ( .I(n440), .Z(n439) );
  BUFFD0 U358 ( .I(n441), .Z(n440) );
  BUFFD0 U359 ( .I(n442), .Z(n441) );
  BUFFD0 U360 ( .I(n443), .Z(n442) );
  BUFFD0 U361 ( .I(n444), .Z(n443) );
  BUFFD0 U362 ( .I(n445), .Z(n444) );
  BUFFD0 U363 ( .I(n446), .Z(n445) );
  BUFFD0 U364 ( .I(n447), .Z(n446) );
  BUFFD0 U365 ( .I(n448), .Z(n447) );
  BUFFD0 U366 ( .I(n449), .Z(n448) );
  BUFFD0 U367 ( .I(n450), .Z(n449) );
  BUFFD0 U368 ( .I(n451), .Z(n450) );
  BUFFD0 U369 ( .I(n452), .Z(n451) );
  BUFFD0 U370 ( .I(n453), .Z(n452) );
  BUFFD0 U371 ( .I(n454), .Z(n453) );
  BUFFD0 U372 ( .I(n455), .Z(n454) );
  BUFFD0 U373 ( .I(n456), .Z(n455) );
  BUFFD0 U374 ( .I(n457), .Z(n456) );
  BUFFD0 U375 ( .I(n458), .Z(n457) );
  BUFFD0 U376 ( .I(n459), .Z(n458) );
  BUFFD0 U377 ( .I(n460), .Z(n459) );
  BUFFD0 U378 ( .I(n461), .Z(n460) );
  BUFFD0 U379 ( .I(n462), .Z(n461) );
  BUFFD0 U380 ( .I(n463), .Z(n462) );
  BUFFD0 U381 ( .I(n928), .Z(n464) );
  BUFFD0 U382 ( .I(n464), .Z(n465) );
  CKBD0 U383 ( .CLK(n466), .C(ReadCmd) );
  BUFFD0 U384 ( .I(n471), .Z(n468) );
  BUFFD0 U385 ( .I(N65), .Z(n469) );
  BUFFD0 U386 ( .I(n469), .Z(n470) );
  BUFFD0 U387 ( .I(n472), .Z(n471) );
  BUFFD0 U388 ( .I(n473), .Z(n472) );
  BUFFD0 U389 ( .I(n474), .Z(n473) );
  BUFFD0 U390 ( .I(n475), .Z(n474) );
  BUFFD0 U391 ( .I(n476), .Z(n475) );
  BUFFD0 U392 ( .I(n477), .Z(n476) );
  BUFFD0 U393 ( .I(n478), .Z(n477) );
  BUFFD0 U394 ( .I(n479), .Z(n478) );
  BUFFD0 U395 ( .I(n480), .Z(n479) );
  BUFFD0 U396 ( .I(n481), .Z(n480) );
  BUFFD0 U397 ( .I(n482), .Z(n481) );
  BUFFD0 U398 ( .I(n483), .Z(n482) );
  BUFFD0 U399 ( .I(n484), .Z(n483) );
  BUFFD0 U400 ( .I(n485), .Z(n484) );
  BUFFD0 U401 ( .I(n486), .Z(n485) );
  BUFFD0 U402 ( .I(n487), .Z(n486) );
  BUFFD0 U403 ( .I(n488), .Z(n487) );
  BUFFD0 U404 ( .I(n489), .Z(n488) );
  BUFFD0 U405 ( .I(n490), .Z(n489) );
  BUFFD0 U406 ( .I(n491), .Z(n490) );
  BUFFD0 U407 ( .I(n492), .Z(n491) );
  BUFFD0 U408 ( .I(n493), .Z(n492) );
  BUFFD0 U409 ( .I(n494), .Z(n493) );
  BUFFD0 U410 ( .I(n495), .Z(n494) );
  BUFFD0 U411 ( .I(n496), .Z(n495) );
  BUFFD0 U412 ( .I(n497), .Z(n496) );
  BUFFD0 U413 ( .I(n498), .Z(n497) );
  BUFFD0 U414 ( .I(n499), .Z(n498) );
  BUFFD0 U415 ( .I(n470), .Z(n499) );
  XNR2D0 U416 ( .A1(n917), .A2(n889), .ZN(n887) );
  BUFFD0 U417 ( .I(n503), .Z(n500) );
  BUFFD0 U418 ( .I(N64), .Z(n501) );
  BUFFD0 U419 ( .I(n501), .Z(n502) );
  BUFFD0 U420 ( .I(n504), .Z(n503) );
  BUFFD0 U421 ( .I(n505), .Z(n504) );
  BUFFD0 U422 ( .I(n506), .Z(n505) );
  BUFFD0 U423 ( .I(n507), .Z(n506) );
  BUFFD0 U424 ( .I(n508), .Z(n507) );
  BUFFD0 U425 ( .I(n509), .Z(n508) );
  BUFFD0 U426 ( .I(n510), .Z(n509) );
  BUFFD0 U427 ( .I(n511), .Z(n510) );
  BUFFD0 U428 ( .I(n512), .Z(n511) );
  BUFFD0 U429 ( .I(n513), .Z(n512) );
  BUFFD0 U430 ( .I(n514), .Z(n513) );
  BUFFD0 U431 ( .I(n515), .Z(n514) );
  BUFFD0 U432 ( .I(n516), .Z(n515) );
  BUFFD0 U433 ( .I(n517), .Z(n516) );
  BUFFD0 U434 ( .I(n518), .Z(n517) );
  BUFFD0 U435 ( .I(n519), .Z(n518) );
  BUFFD0 U436 ( .I(n520), .Z(n519) );
  BUFFD0 U437 ( .I(n521), .Z(n520) );
  BUFFD0 U438 ( .I(n522), .Z(n521) );
  BUFFD0 U439 ( .I(n523), .Z(n522) );
  BUFFD0 U440 ( .I(n524), .Z(n523) );
  BUFFD0 U441 ( .I(n525), .Z(n524) );
  BUFFD0 U442 ( .I(n526), .Z(n525) );
  BUFFD0 U443 ( .I(n527), .Z(n526) );
  BUFFD0 U444 ( .I(n528), .Z(n527) );
  BUFFD0 U445 ( .I(n529), .Z(n528) );
  BUFFD0 U446 ( .I(n530), .Z(n529) );
  BUFFD0 U447 ( .I(n531), .Z(n530) );
  BUFFD0 U448 ( .I(n532), .Z(n531) );
  BUFFD0 U449 ( .I(n502), .Z(n532) );
  OAI21D0 U450 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n883), .ZN(n865) );
  BUFFD0 U451 ( .I(n536), .Z(n533) );
  BUFFD0 U452 ( .I(n833), .Z(n534) );
  BUFFD0 U453 ( .I(n566), .Z(n535) );
  BUFFD0 U454 ( .I(n537), .Z(n536) );
  BUFFD0 U455 ( .I(n539), .Z(n537) );
  BUFFD0 U456 ( .I(n540), .Z(n538) );
  BUFFD0 U457 ( .I(n541), .Z(n539) );
  BUFFD0 U458 ( .I(n542), .Z(n540) );
  BUFFD0 U459 ( .I(n543), .Z(n541) );
  BUFFD0 U460 ( .I(n544), .Z(n542) );
  BUFFD0 U461 ( .I(n545), .Z(n543) );
  BUFFD0 U462 ( .I(n546), .Z(n544) );
  BUFFD0 U463 ( .I(N49), .Z(n545) );
  BUFFD0 U464 ( .I(n547), .Z(n546) );
  BUFFD0 U465 ( .I(n548), .Z(n547) );
  BUFFD0 U466 ( .I(n549), .Z(n548) );
  BUFFD0 U467 ( .I(n550), .Z(n549) );
  BUFFD0 U468 ( .I(n551), .Z(n550) );
  BUFFD0 U469 ( .I(n552), .Z(n551) );
  BUFFD0 U470 ( .I(n553), .Z(n552) );
  BUFFD0 U471 ( .I(n554), .Z(n553) );
  BUFFD0 U472 ( .I(n555), .Z(n554) );
  BUFFD0 U473 ( .I(n556), .Z(n555) );
  BUFFD0 U474 ( .I(n557), .Z(n556) );
  BUFFD0 U475 ( .I(n558), .Z(n557) );
  BUFFD0 U476 ( .I(n559), .Z(n558) );
  BUFFD0 U477 ( .I(n560), .Z(n559) );
  BUFFD0 U478 ( .I(n561), .Z(n560) );
  BUFFD0 U479 ( .I(n562), .Z(n561) );
  BUFFD0 U480 ( .I(n563), .Z(n562) );
  BUFFD0 U481 ( .I(n564), .Z(n563) );
  BUFFD0 U482 ( .I(n565), .Z(n564) );
  BUFFD0 U483 ( .I(n866), .Z(n565) );
  BUFFD0 U484 ( .I(n834), .Z(n566) );
  BUFFD0 U485 ( .I(n569), .Z(n567) );
  BUFFD0 U486 ( .I(n570), .Z(n568) );
  BUFFD0 U487 ( .I(n571), .Z(n569) );
  BUFFD0 U488 ( .I(n572), .Z(n570) );
  BUFFD0 U489 ( .I(n573), .Z(n571) );
  BUFFD0 U490 ( .I(n574), .Z(n572) );
  BUFFD0 U491 ( .I(n575), .Z(n573) );
  BUFFD0 U492 ( .I(n576), .Z(n574) );
  BUFFD0 U493 ( .I(N47), .Z(n575) );
  BUFFD0 U494 ( .I(n577), .Z(n576) );
  BUFFD0 U495 ( .I(n578), .Z(n577) );
  BUFFD0 U496 ( .I(n579), .Z(n578) );
  BUFFD0 U497 ( .I(n580), .Z(n579) );
  BUFFD0 U498 ( .I(n581), .Z(n580) );
  BUFFD0 U499 ( .I(n582), .Z(n581) );
  BUFFD0 U500 ( .I(n583), .Z(n582) );
  BUFFD0 U501 ( .I(n584), .Z(n583) );
  BUFFD0 U502 ( .I(n585), .Z(n584) );
  BUFFD0 U503 ( .I(n586), .Z(n585) );
  BUFFD0 U504 ( .I(n587), .Z(n586) );
  BUFFD0 U505 ( .I(n588), .Z(n587) );
  BUFFD0 U506 ( .I(n589), .Z(n588) );
  BUFFD0 U507 ( .I(n590), .Z(n589) );
  BUFFD0 U508 ( .I(n591), .Z(n590) );
  BUFFD0 U509 ( .I(n592), .Z(n591) );
  BUFFD0 U510 ( .I(n593), .Z(n592) );
  BUFFD0 U511 ( .I(n594), .Z(n593) );
  BUFFD0 U512 ( .I(n595), .Z(n594) );
  BUFFD0 U513 ( .I(n596), .Z(n595) );
  BUFFD0 U514 ( .I(n852), .Z(n596) );
  XNR2D0 U515 ( .A1(n598), .A2(ReadAddr[1]), .ZN(n852) );
  BUFFD0 U516 ( .I(n599), .Z(n597) );
  BUFFD0 U517 ( .I(n600), .Z(n598) );
  BUFFD0 U518 ( .I(n601), .Z(n599) );
  BUFFD0 U519 ( .I(n602), .Z(n600) );
  BUFFD0 U520 ( .I(n603), .Z(n601) );
  BUFFD0 U521 ( .I(n604), .Z(n602) );
  BUFFD0 U522 ( .I(n605), .Z(n603) );
  BUFFD0 U523 ( .I(n606), .Z(n604) );
  BUFFD0 U524 ( .I(n607), .Z(n605) );
  BUFFD0 U525 ( .I(n608), .Z(n606) );
  BUFFD0 U526 ( .I(n609), .Z(n607) );
  BUFFD0 U527 ( .I(n610), .Z(n608) );
  BUFFD0 U528 ( .I(n611), .Z(n609) );
  BUFFD0 U529 ( .I(n612), .Z(n610) );
  BUFFD0 U530 ( .I(n613), .Z(n611) );
  BUFFD0 U531 ( .I(n614), .Z(n612) );
  BUFFD0 U532 ( .I(N46), .Z(n613) );
  BUFFD0 U533 ( .I(n615), .Z(n614) );
  BUFFD0 U534 ( .I(n616), .Z(n615) );
  BUFFD0 U535 ( .I(n617), .Z(n616) );
  BUFFD0 U536 ( .I(n618), .Z(n617) );
  BUFFD0 U537 ( .I(n619), .Z(n618) );
  BUFFD0 U538 ( .I(n620), .Z(n619) );
  BUFFD0 U539 ( .I(n621), .Z(n620) );
  BUFFD0 U540 ( .I(n622), .Z(n621) );
  BUFFD0 U541 ( .I(n623), .Z(n622) );
  BUFFD0 U542 ( .I(n624), .Z(n623) );
  BUFFD0 U543 ( .I(n625), .Z(n624) );
  BUFFD0 U544 ( .I(n626), .Z(n625) );
  BUFFD0 U545 ( .I(ReadAddr[0]), .Z(n626) );
  BUFFD0 U546 ( .I(n649), .Z(n627) );
  BUFFD0 U547 ( .I(n630), .Z(n628) );
  BUFFD0 U548 ( .I(N48), .Z(n629) );
  BUFFD0 U549 ( .I(n632), .Z(n630) );
  BUFFD0 U550 ( .I(n629), .Z(n631) );
  BUFFD0 U551 ( .I(n633), .Z(n632) );
  BUFFD0 U552 ( .I(n635), .Z(n633) );
  BUFFD0 U553 ( .I(n631), .Z(n634) );
  BUFFD0 U554 ( .I(n636), .Z(n635) );
  BUFFD0 U555 ( .I(n637), .Z(n636) );
  BUFFD0 U556 ( .I(n638), .Z(n637) );
  BUFFD0 U557 ( .I(n639), .Z(n638) );
  BUFFD0 U558 ( .I(n640), .Z(n639) );
  BUFFD0 U559 ( .I(n641), .Z(n640) );
  BUFFD0 U560 ( .I(n642), .Z(n641) );
  BUFFD0 U561 ( .I(n643), .Z(n642) );
  BUFFD0 U562 ( .I(n644), .Z(n643) );
  BUFFD0 U563 ( .I(n646), .Z(n644) );
  BUFFD0 U564 ( .I(n926), .Z(n645) );
  BUFFD0 U565 ( .I(n647), .Z(n646) );
  BUFFD0 U566 ( .I(n648), .Z(n647) );
  BUFFD0 U567 ( .I(n1), .Z(n648) );
  CKBXD0 U568 ( .I(n634), .Z(n649) );
  BUFFD0 U569 ( .I(n654), .Z(n650) );
  BUFFD0 U570 ( .I(N63), .Z(n651) );
  BUFFD0 U571 ( .I(n651), .Z(n652) );
  BUFFD0 U572 ( .I(n652), .Z(n653) );
  BUFFD0 U573 ( .I(n655), .Z(n654) );
  BUFFD0 U574 ( .I(n656), .Z(n655) );
  BUFFD0 U575 ( .I(n657), .Z(n656) );
  BUFFD0 U576 ( .I(n658), .Z(n657) );
  BUFFD0 U577 ( .I(n659), .Z(n658) );
  BUFFD0 U578 ( .I(n660), .Z(n659) );
  BUFFD0 U579 ( .I(n661), .Z(n660) );
  BUFFD0 U580 ( .I(n662), .Z(n661) );
  BUFFD0 U581 ( .I(n663), .Z(n662) );
  BUFFD0 U582 ( .I(n664), .Z(n663) );
  BUFFD0 U583 ( .I(n665), .Z(n664) );
  BUFFD0 U584 ( .I(n666), .Z(n665) );
  BUFFD0 U585 ( .I(n667), .Z(n666) );
  BUFFD0 U586 ( .I(n668), .Z(n667) );
  BUFFD0 U587 ( .I(n669), .Z(n668) );
  BUFFD0 U588 ( .I(n670), .Z(n669) );
  BUFFD0 U589 ( .I(n671), .Z(n670) );
  BUFFD0 U590 ( .I(n672), .Z(n671) );
  BUFFD0 U591 ( .I(n673), .Z(n672) );
  BUFFD0 U592 ( .I(n674), .Z(n673) );
  BUFFD0 U593 ( .I(n675), .Z(n674) );
  BUFFD0 U594 ( .I(n676), .Z(n675) );
  BUFFD0 U595 ( .I(n677), .Z(n676) );
  BUFFD0 U596 ( .I(n678), .Z(n677) );
  BUFFD0 U597 ( .I(n679), .Z(n678) );
  BUFFD0 U598 ( .I(n680), .Z(n679) );
  BUFFD0 U599 ( .I(n681), .Z(n680) );
  BUFFD0 U600 ( .I(n682), .Z(n681) );
  BUFFD0 U601 ( .I(n683), .Z(n682) );
  BUFFD0 U602 ( .I(n684), .Z(n683) );
  BUFFD0 U603 ( .I(n653), .Z(n684) );
  BUFFD0 U604 ( .I(n709), .Z(n685) );
  CKBD0 U605 ( .CLK(N66), .C(n686) );
  CKBD0 U606 ( .CLK(n686), .C(n687) );
  CKBD0 U607 ( .CLK(n687), .C(n688) );
  CKBD0 U608 ( .CLK(n688), .C(n689) );
  CKBD0 U609 ( .CLK(n689), .C(n690) );
  CKBD0 U610 ( .CLK(n690), .C(n691) );
  CKBD0 U611 ( .CLK(n691), .C(n692) );
  CKBD0 U612 ( .CLK(n692), .C(n693) );
  CKBD0 U613 ( .CLK(n693), .C(n694) );
  CKBD0 U614 ( .CLK(n694), .C(n695) );
  CKBD0 U615 ( .CLK(n695), .C(n696) );
  CKBD0 U616 ( .CLK(n696), .C(n697) );
  CKBD0 U617 ( .CLK(n697), .C(n698) );
  BUFFD0 U618 ( .I(n924), .Z(n699) );
  BUFFD0 U619 ( .I(n698), .Z(n700) );
  BUFFD0 U620 ( .I(n700), .Z(n701) );
  BUFFD0 U621 ( .I(n701), .Z(n702) );
  BUFFD0 U622 ( .I(n702), .Z(n703) );
  BUFFD0 U623 ( .I(n703), .Z(n704) );
  BUFFD0 U624 ( .I(n704), .Z(n705) );
  BUFFD0 U625 ( .I(n705), .Z(n706) );
  BUFFD0 U626 ( .I(n706), .Z(n707) );
  BUFFD0 U627 ( .I(n707), .Z(n708) );
  CKBD0 U628 ( .CLK(n708), .C(n709) );
  BUFFD0 U629 ( .I(n712), .Z(n710) );
  CKBD0 U630 ( .CLK(CurState[1]), .C(n711) );
  BUFFD0 U631 ( .I(n645), .Z(n712) );
  CKND2D0 U632 ( .A1(n711), .A2(n922), .ZN(n924) );
  BUFFD0 U633 ( .I(n714), .Z(n713) );
  BUFFD0 U634 ( .I(n716), .Z(n714) );
  BUFFD0 U635 ( .I(n717), .Z(n715) );
  BUFFD0 U636 ( .I(n718), .Z(n716) );
  BUFFD0 U637 ( .I(n719), .Z(n717) );
  BUFFD0 U638 ( .I(n720), .Z(n718) );
  BUFFD0 U639 ( .I(n721), .Z(n719) );
  BUFFD0 U640 ( .I(n722), .Z(n720) );
  BUFFD0 U641 ( .I(n723), .Z(n721) );
  BUFFD0 U642 ( .I(n724), .Z(n722) );
  BUFFD0 U643 ( .I(n725), .Z(n723) );
  BUFFD0 U644 ( .I(n726), .Z(n724) );
  BUFFD0 U645 ( .I(n727), .Z(n725) );
  BUFFD0 U646 ( .I(n728), .Z(n726) );
  BUFFD0 U647 ( .I(n729), .Z(n727) );
  BUFFD0 U648 ( .I(n730), .Z(n728) );
  BUFFD0 U649 ( .I(n731), .Z(n729) );
  BUFFD0 U650 ( .I(n732), .Z(n730) );
  BUFFD0 U651 ( .I(n733), .Z(n731) );
  BUFFD0 U652 ( .I(n734), .Z(n732) );
  BUFFD0 U653 ( .I(n735), .Z(n733) );
  BUFFD0 U654 ( .I(n736), .Z(n734) );
  BUFFD0 U655 ( .I(n737), .Z(n735) );
  BUFFD0 U656 ( .I(n738), .Z(n736) );
  BUFFD0 U657 ( .I(n739), .Z(n737) );
  BUFFD0 U658 ( .I(n740), .Z(n738) );
  BUFFD0 U659 ( .I(n741), .Z(n739) );
  BUFFD0 U660 ( .I(n839), .Z(n740) );
  BUFFD0 U661 ( .I(n742), .Z(n741) );
  BUFFD0 U662 ( .I(n743), .Z(n742) );
  BUFFD0 U663 ( .I(n744), .Z(n743) );
  BUFFD0 U664 ( .I(n745), .Z(n744) );
  BUFFD0 U665 ( .I(n746), .Z(n745) );
  BUFFD0 U666 ( .I(n747), .Z(n746) );
  BUFFD0 U667 ( .I(n748), .Z(n747) );
  BUFFD0 U668 ( .I(n849), .Z(n748) );
  BUFFD0 U669 ( .I(n750), .Z(n749) );
  BUFFD0 U670 ( .I(n752), .Z(n750) );
  BUFFD0 U671 ( .I(n753), .Z(n751) );
  BUFFD0 U672 ( .I(n754), .Z(n752) );
  BUFFD0 U673 ( .I(n755), .Z(n753) );
  BUFFD0 U674 ( .I(n756), .Z(n754) );
  BUFFD0 U675 ( .I(n757), .Z(n755) );
  BUFFD0 U676 ( .I(n758), .Z(n756) );
  BUFFD0 U677 ( .I(n759), .Z(n757) );
  BUFFD0 U678 ( .I(n760), .Z(n758) );
  BUFFD0 U679 ( .I(n761), .Z(n759) );
  BUFFD0 U680 ( .I(n762), .Z(n760) );
  BUFFD0 U681 ( .I(n763), .Z(n761) );
  BUFFD0 U682 ( .I(n764), .Z(n762) );
  BUFFD0 U683 ( .I(n765), .Z(n763) );
  BUFFD0 U684 ( .I(n766), .Z(n764) );
  BUFFD0 U685 ( .I(n767), .Z(n765) );
  BUFFD0 U686 ( .I(n768), .Z(n766) );
  BUFFD0 U687 ( .I(n769), .Z(n767) );
  BUFFD0 U688 ( .I(n770), .Z(n768) );
  BUFFD0 U689 ( .I(n771), .Z(n769) );
  BUFFD0 U690 ( .I(n772), .Z(n770) );
  BUFFD0 U691 ( .I(n773), .Z(n771) );
  BUFFD0 U692 ( .I(n774), .Z(n772) );
  BUFFD0 U693 ( .I(n775), .Z(n773) );
  BUFFD0 U694 ( .I(n776), .Z(n774) );
  BUFFD0 U695 ( .I(n777), .Z(n775) );
  BUFFD0 U696 ( .I(n837), .Z(n776) );
  BUFFD0 U697 ( .I(n778), .Z(n777) );
  BUFFD0 U698 ( .I(n779), .Z(n778) );
  BUFFD0 U699 ( .I(n780), .Z(n779) );
  BUFFD0 U700 ( .I(n781), .Z(n780) );
  BUFFD0 U701 ( .I(n782), .Z(n781) );
  BUFFD0 U702 ( .I(n783), .Z(n782) );
  BUFFD0 U703 ( .I(n784), .Z(n783) );
  BUFFD0 U704 ( .I(n848), .Z(n784) );
  BUFFD0 U705 ( .I(n786), .Z(n785) );
  BUFFD0 U706 ( .I(n788), .Z(n786) );
  BUFFD0 U707 ( .I(n789), .Z(n787) );
  BUFFD0 U708 ( .I(n790), .Z(n788) );
  BUFFD0 U709 ( .I(n791), .Z(n789) );
  BUFFD0 U710 ( .I(n792), .Z(n790) );
  BUFFD0 U711 ( .I(n793), .Z(n791) );
  BUFFD0 U712 ( .I(n794), .Z(n792) );
  BUFFD0 U713 ( .I(n795), .Z(n793) );
  BUFFD0 U714 ( .I(n796), .Z(n794) );
  BUFFD0 U715 ( .I(n797), .Z(n795) );
  BUFFD0 U716 ( .I(n798), .Z(n796) );
  BUFFD0 U717 ( .I(n799), .Z(n797) );
  BUFFD0 U718 ( .I(n800), .Z(n798) );
  BUFFD0 U719 ( .I(n801), .Z(n799) );
  BUFFD0 U720 ( .I(n802), .Z(n800) );
  BUFFD0 U721 ( .I(n803), .Z(n801) );
  BUFFD0 U722 ( .I(n804), .Z(n802) );
  BUFFD0 U723 ( .I(n805), .Z(n803) );
  BUFFD0 U724 ( .I(n806), .Z(n804) );
  BUFFD0 U725 ( .I(n807), .Z(n805) );
  BUFFD0 U726 ( .I(n808), .Z(n806) );
  BUFFD0 U727 ( .I(n809), .Z(n807) );
  BUFFD0 U728 ( .I(n810), .Z(n808) );
  BUFFD0 U729 ( .I(n811), .Z(n809) );
  BUFFD0 U730 ( .I(n812), .Z(n810) );
  BUFFD0 U731 ( .I(n813), .Z(n811) );
  BUFFD0 U732 ( .I(n814), .Z(n812) );
  BUFFD0 U733 ( .I(n815), .Z(n813) );
  BUFFD0 U734 ( .I(n816), .Z(n814) );
  BUFFD0 U735 ( .I(n817), .Z(n815) );
  BUFFD0 U736 ( .I(n818), .Z(n816) );
  BUFFD0 U737 ( .I(n819), .Z(n817) );
  BUFFD0 U738 ( .I(n840), .Z(n818) );
  BUFFD0 U739 ( .I(n820), .Z(n819) );
  BUFFD0 U740 ( .I(n821), .Z(n820) );
  BUFFD0 U741 ( .I(n850), .Z(n821) );
  INVD1 U742 ( .I(Reset), .ZN(n829) );
  INVD1 U743 ( .I(Reset), .ZN(n830) );
  INVD1 U744 ( .I(n887), .ZN(n880) );
  INVD1 U745 ( .I(n915), .ZN(n909) );
  MAOI22D0 U746 ( .A1(ReadAddr[0]), .A2(n889), .B1(n918), .B2(n867), .ZN(n864)
         );
  INVD1 U747 ( .I(n889), .ZN(n883) );
  XNR2D1 U748 ( .A1(n880), .A2(ReadAddr[2]), .ZN(n906) );
  ND2D1 U749 ( .A1(n881), .A2(n924), .ZN(n878) );
  NR2D1 U750 ( .A1(n894), .A2(n885), .ZN(n922) );
  ND2D1 U751 ( .A1(n881), .A2(n926), .ZN(n916) );
  NR2D1 U752 ( .A1(n598), .A2(n856), .ZN(N46) );
  NR2D1 U753 ( .A1(n538), .A2(n856), .ZN(N49) );
  NR2D1 U754 ( .A1(n568), .A2(n856), .ZN(N47) );
  OAI211D1 U755 ( .A1(CurState[1]), .A2(n885), .B(n881), .C(n861), .ZN(n915)
         );
  AOI21D1 U756 ( .A1(WriteReq), .A2(n921), .B(n860), .ZN(n861) );
  AOI21D1 U757 ( .A1(CurState[0]), .A2(n859), .B(n894), .ZN(n860) );
  OAI33D1 U758 ( .A1(n879), .A2(n921), .A3(n878), .B1(n877), .B2(n876), .B3(
        n875), .ZN(n838) );
  INVD1 U759 ( .I(WriteCmd), .ZN(n879) );
  XNR2D1 U760 ( .A1(n917), .A2(n291), .ZN(n875) );
  XNR2D1 U761 ( .A1(n918), .A2(n290), .ZN(n876) );
  ND2D1 U762 ( .A1(WriteReq), .A2(n916), .ZN(n919) );
  OAI22D0 U763 ( .A1(n915), .A2(n715), .B1(n909), .B2(n903), .ZN(n839) );
  AOI31D0 U764 ( .A1(n902), .A2(n901), .A3(n900), .B(n921), .ZN(n903) );
  IIND4D1 U765 ( .A1(n893), .A2(n891), .B1(n886), .B2(n885), .ZN(n901) );
  AOI31D0 U766 ( .A1(n832), .A2(CurState[0]), .A3(n899), .B(n898), .ZN(n900)
         );
  OAI22D0 U767 ( .A1(n915), .A2(n751), .B1(n909), .B2(n873), .ZN(n837) );
  AOI21D1 U768 ( .A1(CurState[1]), .A2(n872), .B(n922), .ZN(n873) );
  OAI21D1 U769 ( .A1(CurState[2]), .A2(n871), .B(n870), .ZN(n872) );
  AOI22D0 U770 ( .A1(n907), .A2(ReadAddr[2]), .B1(n834), .B2(n908), .ZN(n871)
         );
  OAI31D0 U771 ( .A1(n926), .A2(WriteReq), .A3(Reset), .B(n925), .ZN(n847) );
  OAI31D0 U772 ( .A1(CurState[0]), .A2(Reset), .A3(CurState[2]), .B(EmptyFIFO), 
        .ZN(n925) );
  OAI21D1 U773 ( .A1(n915), .A2(n787), .B(n914), .ZN(n840) );
  OAI211D1 U774 ( .A1(CurState[2]), .A2(n913), .B(CurState[0]), .C(n912), .ZN(
        n914) );
  NR4D0 U775 ( .A1(n906), .A2(n905), .A3(n910), .A4(n904), .ZN(n913) );
  AOI21D1 U776 ( .A1(n911), .A2(n910), .B(n909), .ZN(n912) );
  ND3D1 U777 ( .A1(n874), .A2(n916), .A3(WriteReq), .ZN(n877) );
  XNR2D1 U778 ( .A1(WriteAddr[0]), .A2(n292), .ZN(n874) );
  MAOI22D0 U779 ( .A1(WriteAddr[0]), .A2(n862), .B1(n833), .B2(n867), .ZN(n863) );
  OAI33D1 U780 ( .A1(ReadAddr[1]), .A2(WriteAddr[2]), .A3(n864), .B1(n917), 
        .B2(WriteAddr[1]), .B3(n863), .ZN(n908) );
  OAI33D1 U781 ( .A1(ReadAddr[1]), .A2(n864), .A3(n917), .B1(n863), .B2(
        WriteAddr[2]), .B3(WriteAddr[1]), .ZN(n907) );
  NR2D1 U782 ( .A1(n918), .A2(n831), .ZN(n889) );
  XOR2D1 U783 ( .A1(n865), .A2(n833), .Z(n905) );
  AOI31D0 U784 ( .A1(n831), .A2(CurState[0]), .A3(n882), .B(n881), .ZN(n902)
         );
  NR3D0 U785 ( .A1(n905), .A2(n832), .A3(n906), .ZN(n882) );
  OAI31D0 U786 ( .A1(n869), .A2(n868), .A3(n904), .B(CurState[0]), .ZN(n870)
         );
  XNR2D1 U787 ( .A1(WriteAddr[2]), .A2(n866), .ZN(n868) );
  INVD1 U788 ( .I(n905), .ZN(n869) );
  NR3D0 U789 ( .A1(n905), .A2(n831), .A3(n890), .ZN(n899) );
  AOI21D1 U790 ( .A1(n893), .A2(n889), .B(n888), .ZN(n890) );
  OAI32D1 U791 ( .A1(n917), .A2(n834), .A3(n889), .B1(ReadAddr[2]), .B2(n887), 
        .ZN(n888) );
  AO22D0 U792 ( .A1(ReadAddr[2]), .A2(n908), .B1(n907), .B2(n834), .Z(n911) );
  OAI222D0 U793 ( .A1(n917), .A2(ReadAddr[2]), .B1(n918), .B2(ReadAddr[1]), 
        .C1(n831), .C2(ReadAddr[0]), .ZN(n891) );
  AOI22D0 U794 ( .A1(n894), .A2(CurState[1]), .B1(n910), .B2(n922), .ZN(n881)
         );
  NR3D0 U795 ( .A1(n711), .A2(CurState[2]), .A3(CurState[0]), .ZN(n921) );
  OAI21D1 U796 ( .A1(n831), .A2(n832), .B(n867), .ZN(n904) );
  OAI32D0 U797 ( .A1(n924), .A2(Reset), .A3(ReadReq), .B1(n923), .B2(n7), .ZN(
        n846) );
  ND2D1 U798 ( .A1(n929), .A2(n699), .ZN(n853) );
  OAI211D1 U799 ( .A1(n831), .A2(ReadAddr[1]), .B(n884), .C(n883), .ZN(n886)
         );
  OAI21D1 U800 ( .A1(WriteAddr[1]), .A2(n833), .B(n832), .ZN(n884) );
  CKND2D0 U801 ( .A1(ReadReq), .A2(n878), .ZN(n920) );
  NR2D1 U802 ( .A1(WriteAddr[2]), .A2(n834), .ZN(n893) );
  ND2D1 U803 ( .A1(n831), .A2(n832), .ZN(n867) );
  OAI22D0 U804 ( .A1(n832), .A2(n699), .B1(WriteAddr[0]), .B2(n853), .ZN(N63)
         );
  OAI22D0 U805 ( .A1(n535), .A2(n699), .B1(n880), .B2(n853), .ZN(N65) );
  OAI22D0 U806 ( .A1(n534), .A2(n699), .B1(n865), .B2(n853), .ZN(N64) );
  AOI31D0 U807 ( .A1(n897), .A2(n896), .A3(n895), .B(n894), .ZN(n898) );
  AOI22D0 U808 ( .A1(n893), .A2(ReadAddr[1]), .B1(n831), .B2(ReadAddr[0]), 
        .ZN(n895) );
  OAI21D1 U809 ( .A1(n893), .A2(n891), .B(n918), .ZN(n897) );
  OAI21D1 U810 ( .A1(ReadAddr[1]), .A2(n892), .B(n891), .ZN(n896) );
  OAI32D1 U811 ( .A1(n858), .A2(n857), .A3(n859), .B1(n878), .B2(n856), .ZN(
        n836) );
  XNR2D1 U812 ( .A1(n833), .A2(n269), .ZN(n857) );
  ND3D1 U813 ( .A1(n855), .A2(n878), .A3(n854), .ZN(n858) );
  XNR2D1 U814 ( .A1(ReadAddr[2]), .A2(n271), .ZN(n855) );
  NR2D1 U815 ( .A1(n832), .A2(n534), .ZN(n862) );
  XOR2D1 U816 ( .A1(n862), .A2(n535), .Z(n866) );
  XNR2D1 U817 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n892) );
  XNR2D1 U818 ( .A1(ReadAddr[0]), .A2(n270), .ZN(n854) );
  ND2D1 U819 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  INVD0 U820 ( .I(ReadReq), .ZN(n859) );
endmodule


module DPMem1kx32_AWid3_DWid32_1 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [2:0] AddrR;
  input [2:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N48, N49, N50, ClockW, Dreadyr, \Storage[7][32] , \Storage[7][31] ,
         \Storage[7][30] , \Storage[7][29] , \Storage[7][28] ,
         \Storage[7][27] , \Storage[7][26] , \Storage[7][25] ,
         \Storage[7][24] , \Storage[7][23] , \Storage[7][22] ,
         \Storage[7][21] , \Storage[7][20] , \Storage[7][19] ,
         \Storage[7][18] , \Storage[7][17] , \Storage[7][16] ,
         \Storage[7][15] , \Storage[7][14] , \Storage[7][13] ,
         \Storage[7][12] , \Storage[7][11] , \Storage[7][10] , \Storage[7][9] ,
         \Storage[7][8] , \Storage[7][7] , \Storage[7][6] , \Storage[7][5] ,
         \Storage[7][4] , \Storage[7][3] , \Storage[7][2] , \Storage[7][1] ,
         \Storage[7][0] , \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N87, N99, N194, N227, N293, N359, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373;
  wire   [31:0] DataOr;
  assign N48 = AddrR[0];
  assign N49 = AddrR[1];
  assign N50 = AddrR[2];

  XNR4D1 U13 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n4361) );
  XOR4D1 U14 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n4362) );
  XOR4D1 U15 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n4365) );
  XOR4D1 U16 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n4368) );
  XNR4D1 U17 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n4371) );
  XOR4D1 U21 ( .A1(n4356), .A2(N74), .A3(n4355), .A4(N77), .Z(n4357) );
  XNR4D1 U22 ( .A1(N71), .A2(N70), .A3(N73), .A4(N72), .ZN(n4355) );
  XNR4D1 U27 ( .A1(N53), .A2(N52), .A3(N55), .A4(N54), .ZN(n4349) );
  XOR4D1 U28 ( .A1(N57), .A2(N56), .A3(N59), .A4(N58), .Z(n4350) );
  XNR4D1 U29 ( .A1(N64), .A2(N63), .A3(N66), .A4(N65), .ZN(n4353) );
  XNR4D1 U30 ( .A1(N82), .A2(N80), .A3(N84), .A4(N83), .ZN(n4359) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(n4302), .CP(n4315), .CDN(
        n4340), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n4304), .CP(n4311), .CDN(
        n4343), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n4304), .CP(n4311), .CDN(
        n4337), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n4304), .CP(n4311), .CDN(
        n4339), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(n4304), .CP(n4315), .CDN(
        n4339), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n4304), .CP(n4318), .CDN(
        n4338), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n4304), .CP(n4322), .CDN(
        n4339), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n4302), .CP(n4310), .CDN(
        n4337), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n4302), .CP(n4315), .CDN(
        n4339), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n4302), .CP(n4314), .CDN(
        n4339), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n4302), .CP(n4320), .CDN(
        n4339), .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n4302), .CP(n4321), .CDN(
        n4337), .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(n4302), .CP(ClockW), .CDN(
        n4339), .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n4302), .CP(n4320), .CDN(
        n4338), .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(n4302), .CP(ClockW), .CDN(
        n4339), .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n4302), .CP(n4320), .CDN(
        n4339), .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(n4302), .CP(n4313), .CDN(
        n4339), .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n4302), .CP(n4318), .CDN(
        n4337), .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(n4302), .CP(n4310), .CDN(
        n4339), .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(n4302), .CP(n4311), .CDN(
        n4338), .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n4308), .CP(n4317), .CDN(
        n4336), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(n4307), .CP(n4317), .CDN(
        n4340), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n4307), .CP(n4318), .CDN(
        n4330), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n4307), .CP(n4318), .CDN(
        n4335), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(n4307), .CP(n4318), .CDN(
        n4340), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(n4307), .CP(n4318), .CDN(
        n4344), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(n4307), .CP(n4318), .CDN(
        n4336), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n4308), .CP(n4318), .CDN(
        n4344), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(n4308), .CP(n4313), .CDN(
        n4343), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(n4308), .CP(n4320), .CDN(
        n4335), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n4308), .CP(n4315), .CDN(
        n4340), .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(n4308), .CP(n4316), .CDN(
        n4334), .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(n4308), .CP(n4317), .CDN(
        n4343), .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(n4308), .CP(n4313), .CDN(
        n4342), .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(n4308), .CP(n4310), .CDN(
        n4343), .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n4308), .CP(n4322), .CDN(
        n4331), .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(n4308), .CP(n4321), .CDN(
        n4341), .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(N99), .CP(n4319), .CDN(n4341), .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(N99), .CP(n4319), .CDN(n4331), .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(N99), .CP(n4319), .CDN(n4331), .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n4292), .CP(n4311), .CDN(
        n4332), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n4292), .CP(ClockW), .CDN(
        n4332), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n4292), .CP(n4313), .CDN(
        n4332), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n4292), .CP(n4314), .CDN(
        n4332), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n4292), .CP(n4310), .CDN(
        n4332), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(n4292), .CP(ClockW), .CDN(
        n4332), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(n4292), .CP(n4321), .CDN(
        n4332), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n4293), .CP(n4319), .CDN(
        n4332), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n4293), .CP(n4319), .CDN(
        n4332), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n4293), .CP(n4320), .CDN(
        n4332), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n4293), .CP(n4322), .CDN(
        n4344), .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(n4293), .CP(n4321), .CDN(
        n4341), .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(n4293), .CP(n4310), .CDN(
        n4344), .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(n4293), .CP(n4313), .CDN(
        n4341), .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(n4293), .CP(n4318), .CDN(
        n4344), .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n4293), .CP(n4315), .CDN(
        n4341), .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n4293), .CP(n4316), .CDN(
        n4344), .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n4293), .CP(n4314), .CDN(
        n4341), .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n4292), .CP(n4314), .CDN(
        n4344), .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n4293), .CP(n4314), .CDN(
        n4341), .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(N293), .CP(n4321), .CDN(
        n4334), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n4295), .CP(n4320), .CDN(
        n4344), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n4295), .CP(n4315), .CDN(
        n4330), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n4295), .CP(n4312), .CDN(
        n4342), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n4295), .CP(n4322), .CDN(
        n4337), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(n4295), .CP(n4320), .CDN(
        n4344), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n4295), .CP(ClockW), .CDN(
        n4334), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n4296), .CP(n4312), .CDN(
        n4330), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n4296), .CP(n4315), .CDN(
        n4342), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n4296), .CP(n4312), .CDN(
        n4336), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n4296), .CP(n4318), .CDN(
        n4331), .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(n4296), .CP(n4310), .CDN(
        n4331), .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(n4296), .CP(n4310), .CDN(
        n4331), .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n4296), .CP(n4316), .CDN(
        n4331), .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(n4296), .CP(n4319), .CDN(
        n4331), .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n4296), .CP(n4312), .CDN(
        n4331), .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n4296), .CP(n4322), .CDN(
        n4331), .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(N293), .CP(n4314), .CDN(
        n4331), .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(n4296), .CP(n4321), .CDN(
        n4331), .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n4295), .CP(n4315), .CDN(
        n4331), .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(n4298), .CP(n4312), .CDN(
        n4330), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n4297), .CP(n4317), .CDN(
        n4330), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n4297), .CP(n4314), .CDN(
        n4342), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n4297), .CP(n4314), .CDN(
        n4341), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(n4298), .CP(n4312), .CDN(
        n4340), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(n4297), .CP(n4319), .CDN(
        n4341), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(n4298), .CP(n4318), .CDN(
        n4337), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n4297), .CP(n4311), .CDN(
        n4335), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n4297), .CP(n4317), .CDN(
        n4337), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n4297), .CP(n4314), .CDN(
        n4334), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n4297), .CP(n4319), .CDN(
        n4341), .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(n4297), .CP(n4322), .CDN(
        n4336), .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(n4297), .CP(ClockW), .CDN(
        n4338), .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(n4297), .CP(n4311), .CDN(
        n4331), .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(n4297), .CP(n4310), .CDN(
        n4338), .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n4297), .CP(n4321), .CDN(
        n4344), .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(n4297), .CP(n4311), .CDN(
        n4345), .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n4298), .CP(n4317), .CDN(
        n4344), .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(n4298), .CP(n4321), .CDN(
        n4331), .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(n4298), .CP(ClockW), .CDN(
        n4331), .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(N227), .CP(n4314), .CDN(
        n4333), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n4299), .CP(n4320), .CDN(
        n4343), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n4299), .CP(n4321), .CDN(
        n4343), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n4299), .CP(n4317), .CDN(
        n4342), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(n4299), .CP(ClockW), .CDN(
        n4342), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n4299), .CP(n4314), .CDN(
        n4345), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(n4299), .CP(n4319), .CDN(
        n4340), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n4300), .CP(n4315), .CDN(
        n4345), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n4300), .CP(n4310), .CDN(
        n4336), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n4300), .CP(n4311), .CDN(
        n4342), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n4300), .CP(n4320), .CDN(
        n4338), .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n4300), .CP(n4322), .CDN(
        n4344), .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(n4300), .CP(n4311), .CDN(
        n4340), .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(n4300), .CP(n4319), .CDN(
        n4340), .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(n4300), .CP(n4321), .CDN(
        n4340), .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n4300), .CP(n4310), .CDN(
        n4343), .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(n4300), .CP(n4322), .CDN(
        n4340), .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n4300), .CP(n4321), .CDN(
        n4334), .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(N227), .CP(n4320), .CDN(
        n4340), .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(N227), .CP(n4319), .CDN(
        n4341), .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n4305), .CP(n4310), .CDN(
        n4345), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n4305), .CP(n4317), .CDN(
        n4345), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n4305), .CP(n4310), .CDN(
        n4342), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n4305), .CP(n4317), .CDN(
        n4344), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n4305), .CP(n4318), .CDN(
        n4334), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(n4305), .CP(n4315), .CDN(
        n4332), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(n4305), .CP(n4315), .CDN(
        n4333), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n4306), .CP(n4315), .CDN(
        n4337), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n4306), .CP(n4315), .CDN(
        n4341), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n4306), .CP(n4315), .CDN(
        n4342), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n4306), .CP(n4315), .CDN(
        n4343), .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(n4306), .CP(n4315), .CDN(
        n4339), .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(n4306), .CP(n4315), .CDN(
        n4336), .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(n4306), .CP(n4315), .CDN(
        n4344), .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(n4306), .CP(n4316), .CDN(
        n4341), .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n4306), .CP(n4316), .CDN(
        n4342), .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n4306), .CP(n4316), .CDN(
        n4340), .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n4305), .CP(n4316), .CDN(
        n4340), .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n4305), .CP(n4316), .CDN(
        n4342), .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n4306), .CP(n4316), .CDN(
        n4345), .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(N359), .CP(n4313), .CDN(
        n4335), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n4289), .CP(n4313), .CDN(
        n4335), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n4289), .CP(n4313), .CDN(
        n4334), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(n4289), .CP(n4313), .CDN(
        n4334), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(n4289), .CP(n4313), .CDN(
        n4334), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(n4289), .CP(n4319), .CDN(
        n4334), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(n4289), .CP(n4313), .CDN(
        n4334), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n4290), .CP(n4318), .CDN(
        n4334), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n4290), .CP(n4312), .CDN(
        n4334), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n4290), .CP(n4311), .CDN(
        n4334), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n4290), .CP(n4317), .CDN(
        n4333), .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(n4290), .CP(n4318), .CDN(
        n4333), .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(n4290), .CP(n4315), .CDN(
        n4333), .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(n4290), .CP(n4316), .CDN(
        n4333), .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(n4290), .CP(n4312), .CDN(
        n4333), .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n4290), .CP(n4320), .CDN(
        n4333), .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n4290), .CP(n4310), .CDN(
        n4333), .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n4290), .CP(n4318), .CDN(
        n4333), .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(N359), .CP(n4319), .CDN(
        n4333), .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(N359), .CP(n4320), .CDN(
        n4333), .Q(\Storage[7][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n1768), .CP(n4323), .CDN(n4342), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N87), .E(n4302), .CP(n4313), .CDN(n4340), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(n4302), .CP(n4310), .CDN(
        n4344), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(N194), .CP(n4316), .CDN(
        n4340), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(N194), .CP(n4316), .CDN(
        n4343), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(N194), .CP(ClockW), .CDN(
        n4342), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(N194), .CP(n4322), .CDN(
        n4341), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(N194), .CP(n4316), .CDN(
        n4334), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(N194), .CP(n4320), .CDN(
        n4343), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(N194), .CP(n4322), .CDN(
        n4336), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n4304), .CP(n4321), .CDN(
        n4343), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n4304), .CP(n4320), .CDN(
        n4339), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n4304), .CP(ClockW), .CDN(
        n4338), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n4304), .CP(n4310), .CDN(
        n4339), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N87), .E(n4307), .CP(n4316), .CDN(n4335), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(n4308), .CP(n4316), .CDN(
        n4343), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n4307), .CP(n4316), .CDN(
        n4335), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(n4308), .CP(n4317), .CDN(
        n4341), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(N99), .CP(n4317), .CDN(
        n4333), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(N99), .CP(n4317), .CDN(
        n4330), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(N99), .CP(n4317), .CDN(
        n4336), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(N99), .CP(n4317), .CDN(
        n4341), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n4307), .CP(n4317), .CDN(
        n4342), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n4307), .CP(n4317), .CDN(
        n4345), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(n4307), .CP(n4318), .CDN(
        n4340), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(n4307), .CP(n4318), .CDN(
        n4339), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(n4307), .CP(n4318), .CDN(
        n4344), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N87), .E(n4292), .CP(n4311), .CDN(n4333), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(n4293), .CP(ClockW), .CDN(
        n4332), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(n4292), .CP(n4321), .CDN(
        n4332), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n4293), .CP(n4322), .CDN(
        n4332), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(n4292), .CP(n4321), .CDN(
        n4332), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(n4293), .CP(n4312), .CDN(
        n4332), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(n4292), .CP(n4314), .CDN(
        n4332), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(n4293), .CP(n4318), .CDN(
        n4332), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n4292), .CP(n4312), .CDN(
        n4332), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(n4292), .CP(n4311), .CDN(
        n4332), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n4292), .CP(n4320), .CDN(
        n4333), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n4292), .CP(n4311), .CDN(
        n4333), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n4292), .CP(n4322), .CDN(
        n4333), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N87), .E(n4295), .CP(n4314), .CDN(n4344), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(n4296), .CP(n4314), .CDN(
        n4333), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(n4295), .CP(n4314), .CDN(
        n4330), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(n4296), .CP(n4314), .CDN(
        n4342), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(N293), .CP(n4314), .CDN(
        n4335), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(N293), .CP(n4314), .CDN(
        n4333), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(N293), .CP(n4319), .CDN(
        n4342), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(N293), .CP(n4317), .CDN(
        n4330), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(N293), .CP(n4310), .CDN(
        n4335), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(n4295), .CP(n4310), .CDN(
        n4334), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n4295), .CP(n4317), .CDN(
        n4330), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n4295), .CP(ClockW), .CDN(
        n4341), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n4295), .CP(n4311), .CDN(
        n4330), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N87), .E(n4298), .CP(n4313), .CDN(n4331), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(n4298), .CP(ClockW), .CDN(
        n4330), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(n4298), .CP(n4320), .CDN(
        n4330), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(n4298), .CP(n4319), .CDN(
        n4330), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n4298), .CP(n4314), .CDN(
        n4330), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n4298), .CP(n4322), .CDN(
        n4330), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n4298), .CP(n4311), .CDN(
        n4330), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(n4298), .CP(n4321), .CDN(
        n4330), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n4298), .CP(n4322), .CDN(
        n4330), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(n4297), .CP(n4311), .CDN(
        n4330), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n4298), .CP(n4322), .CDN(
        n4342), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n4297), .CP(n4319), .CDN(
        n4339), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n4298), .CP(n4317), .CDN(
        n4331), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N87), .E(n4299), .CP(n4321), .CDN(n4331), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(n4300), .CP(n4318), .CDN(
        n4340), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(n4299), .CP(n4320), .CDN(
        n4343), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(n4300), .CP(n4315), .CDN(
        n4343), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(n4299), .CP(ClockW), .CDN(
        n4331), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(N227), .CP(n4320), .CDN(
        n4345), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(N227), .CP(n4321), .CDN(
        n4342), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(N227), .CP(n4316), .CDN(
        n4341), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(N227), .CP(n4311), .CDN(
        n4345), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n4299), .CP(n4319), .CDN(
        n4343), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n4299), .CP(n4322), .CDN(
        n4343), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n4299), .CP(n4313), .CDN(
        n4340), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n4299), .CP(n4319), .CDN(
        n4343), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N87), .E(n4306), .CP(n4313), .CDN(n4339), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(n4306), .CP(n4312), .CDN(
        n4345), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(n4305), .CP(n4321), .CDN(
        n4345), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(n4306), .CP(n4322), .CDN(
        n4345), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(n4305), .CP(n4316), .CDN(
        n4345), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(n4306), .CP(n4316), .CDN(
        n4345), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(n4305), .CP(n4313), .CDN(
        n4345), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(n4306), .CP(n4320), .CDN(
        n4345), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n4305), .CP(n4316), .CDN(
        n4345), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(n4305), .CP(n4311), .CDN(
        n4345), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n4305), .CP(n4322), .CDN(
        n4342), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n4305), .CP(n4319), .CDN(
        n4330), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n4305), .CP(ClockW), .CDN(
        n4335), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N87), .E(n4289), .CP(n4312), .CDN(n4336), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(n4290), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(n4289), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n4290), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n4289), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(N359), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(N359), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(N359), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(N359), .CP(n4312), .CDN(
        n4335), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(n4289), .CP(n4313), .CDN(
        n4335), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n4289), .CP(n4313), .CDN(
        n4334), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n4289), .CP(n4313), .CDN(
        n4334), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n4289), .CP(n4313), .CDN(
        n4334), .Q(\Storage[7][18] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n1831), .E(n4326), .CP(n4324), .CDN(n4339), 
        .Q(DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n1901), .E(n4326), .CP(n4324), .CDN(n4338), 
        .Q(DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n1971), .E(n4326), .CP(n4323), .CDN(n4338), 
        .Q(DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n2041), .E(n4326), .CP(n4324), .CDN(n4338), 
        .Q(DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n2111), .E(n4326), .CP(n4323), .CDN(n4338), 
        .Q(DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n2181), .E(n4326), .CP(n4324), .CDN(n4338), 
        .Q(DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n2251), .E(n4326), .CP(n4323), .CDN(n4338), 
        .Q(DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n2321), .E(n4326), .CP(n4324), .CDN(n4338), 
        .Q(DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n2391), .E(n4326), .CP(n4323), .CDN(n4338), 
        .Q(DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n2461), .E(n4326), .CP(n4323), .CDN(n4338), 
        .Q(DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n2531), .E(n4326), .CP(n4323), .CDN(n4338), 
        .Q(DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n2601), .E(n4326), .CP(n4323), .CDN(n4338), 
        .Q(DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n2671), .E(n4326), .CP(n4323), .CDN(n4337), 
        .Q(DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n2741), .E(n4326), .CP(n4323), .CDN(n4337), 
        .Q(DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n2811), .E(n4326), .CP(n4323), .CDN(n4337), 
        .Q(DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n2881), .E(n4326), .CP(n4323), .CDN(n4337), 
        .Q(DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n2951), .E(n4326), .CP(n4323), .CDN(n4337), 
        .Q(DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n3021), .E(n4325), .CP(n4323), .CDN(n4337), 
        .Q(DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n3091), .E(n4325), .CP(n4324), .CDN(n4337), 
        .Q(DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n3161), .E(n4325), .CP(n4324), .CDN(n4337), 
        .Q(DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n3231), .E(n4325), .CP(n4324), .CDN(n4337), 
        .Q(DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n3301), .E(n4325), .CP(n4324), .CDN(n4337), 
        .Q(DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n3371), .E(n4325), .CP(n4324), .CDN(n4337), 
        .Q(DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n3441), .E(n4325), .CP(n4324), .CDN(n4336), 
        .Q(DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n3510), .E(n4325), .CP(n4324), .CDN(n4336), 
        .Q(DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n3580), .E(n4325), .CP(n4324), .CDN(n4336), 
        .Q(DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n3650), .E(n4325), .CP(n4324), .CDN(n4336), 
        .Q(DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n3720), .E(n4325), .CP(n4324), .CDN(n4336), 
        .Q(DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n1), .E(n4325), .CP(n4323), .CDN(n4336), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n3857), .E(n4325), .CP(n4323), .CDN(n4336), 
        .Q(DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n3926), .E(n4325), .CP(n4324), .CDN(n4336), 
        .Q(DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n3995), .E(n4325), .CP(n4324), .CDN(n4336), 
        .Q(DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(n4066), .E(n4325), .CP(n4323), .CDN(n4336), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(n1713), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(n1658), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(n1603), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(n1548), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(n1493), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(n1439), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(n1385), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(n1331), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(n1277), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(n1223), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(n1169), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(n1115), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(n1061), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(n1007), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(n953), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(n899), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(n845), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(n791), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(n737), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(n683), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(n629), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(n575), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(n521), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(n467), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(n413), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(n359), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(n305), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(n251), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(n197), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(n143), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(n61), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(n7), .OE(ChipEna), .Z(DataO[31]) );
  BUFFD0 U3 ( .I(n3789), .Z(n1) );
  BUFFD0 U4 ( .I(n4132), .Z(n2) );
  OR3D1 U5 ( .A1(n4348), .A2(AddrW[0]), .A3(n4347), .Z(n3) );
  CKND2D0 U6 ( .A1(ClkR), .A2(ChipEna), .ZN(n4) );
  OR3D1 U7 ( .A1(n4346), .A2(AddrW[1]), .A3(n4373), .Z(n5) );
  OR3D1 U8 ( .A1(n4347), .A2(AddrW[1]), .A3(AddrW[0]), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(n10), .Z(n9) );
  BUFFD0 U12 ( .I(n11), .Z(n10) );
  BUFFD0 U18 ( .I(n12), .Z(n11) );
  BUFFD0 U19 ( .I(n13), .Z(n12) );
  BUFFD0 U20 ( .I(n14), .Z(n13) );
  BUFFD0 U23 ( .I(n15), .Z(n14) );
  BUFFD0 U24 ( .I(n16), .Z(n15) );
  BUFFD0 U25 ( .I(n17), .Z(n16) );
  BUFFD0 U26 ( .I(n18), .Z(n17) );
  BUFFD0 U31 ( .I(n19), .Z(n18) );
  BUFFD0 U32 ( .I(n20), .Z(n19) );
  BUFFD0 U33 ( .I(n21), .Z(n20) );
  BUFFD0 U34 ( .I(n22), .Z(n21) );
  BUFFD0 U35 ( .I(n23), .Z(n22) );
  BUFFD0 U36 ( .I(n24), .Z(n23) );
  BUFFD0 U37 ( .I(n25), .Z(n24) );
  BUFFD0 U38 ( .I(n26), .Z(n25) );
  BUFFD0 U39 ( .I(n27), .Z(n26) );
  BUFFD0 U40 ( .I(n28), .Z(n27) );
  BUFFD0 U41 ( .I(n29), .Z(n28) );
  BUFFD0 U42 ( .I(n30), .Z(n29) );
  BUFFD0 U43 ( .I(n31), .Z(n30) );
  BUFFD0 U44 ( .I(n32), .Z(n31) );
  BUFFD0 U45 ( .I(n33), .Z(n32) );
  BUFFD0 U46 ( .I(n34), .Z(n33) );
  BUFFD0 U47 ( .I(n35), .Z(n34) );
  BUFFD0 U48 ( .I(n36), .Z(n35) );
  BUFFD0 U49 ( .I(n37), .Z(n36) );
  BUFFD0 U50 ( .I(n38), .Z(n37) );
  BUFFD0 U51 ( .I(n39), .Z(n38) );
  BUFFD0 U52 ( .I(n40), .Z(n39) );
  BUFFD0 U53 ( .I(n41), .Z(n40) );
  BUFFD0 U54 ( .I(n42), .Z(n41) );
  BUFFD0 U55 ( .I(n43), .Z(n42) );
  BUFFD0 U56 ( .I(n44), .Z(n43) );
  BUFFD0 U57 ( .I(n45), .Z(n44) );
  BUFFD0 U58 ( .I(n46), .Z(n45) );
  BUFFD0 U59 ( .I(n47), .Z(n46) );
  BUFFD0 U60 ( .I(n48), .Z(n47) );
  BUFFD0 U61 ( .I(n49), .Z(n48) );
  BUFFD0 U62 ( .I(n50), .Z(n49) );
  BUFFD0 U63 ( .I(n51), .Z(n50) );
  BUFFD0 U64 ( .I(n52), .Z(n51) );
  BUFFD0 U65 ( .I(n53), .Z(n52) );
  BUFFD0 U66 ( .I(n54), .Z(n53) );
  BUFFD0 U67 ( .I(n55), .Z(n54) );
  BUFFD0 U68 ( .I(n56), .Z(n55) );
  BUFFD0 U69 ( .I(n57), .Z(n56) );
  BUFFD0 U70 ( .I(n58), .Z(n57) );
  BUFFD0 U71 ( .I(n59), .Z(n58) );
  BUFFD0 U72 ( .I(n60), .Z(n59) );
  BUFFD0 U73 ( .I(DataOr[31]), .Z(n60) );
  BUFFD0 U74 ( .I(n62), .Z(n61) );
  BUFFD0 U75 ( .I(n63), .Z(n62) );
  BUFFD0 U76 ( .I(n64), .Z(n63) );
  BUFFD0 U77 ( .I(n65), .Z(n64) );
  BUFFD0 U78 ( .I(n94), .Z(n65) );
  BUFFD0 U79 ( .I(n95), .Z(n94) );
  BUFFD0 U80 ( .I(n96), .Z(n95) );
  BUFFD0 U81 ( .I(n97), .Z(n96) );
  BUFFD0 U82 ( .I(n98), .Z(n97) );
  BUFFD0 U83 ( .I(n99), .Z(n98) );
  BUFFD0 U84 ( .I(n100), .Z(n99) );
  BUFFD0 U85 ( .I(n101), .Z(n100) );
  BUFFD0 U86 ( .I(n102), .Z(n101) );
  BUFFD0 U87 ( .I(n103), .Z(n102) );
  BUFFD0 U88 ( .I(n104), .Z(n103) );
  BUFFD0 U89 ( .I(n105), .Z(n104) );
  BUFFD0 U90 ( .I(n106), .Z(n105) );
  BUFFD0 U91 ( .I(n107), .Z(n106) );
  BUFFD0 U92 ( .I(n108), .Z(n107) );
  BUFFD0 U93 ( .I(n109), .Z(n108) );
  BUFFD0 U94 ( .I(n110), .Z(n109) );
  BUFFD0 U95 ( .I(n111), .Z(n110) );
  BUFFD0 U96 ( .I(n112), .Z(n111) );
  BUFFD0 U97 ( .I(n113), .Z(n112) );
  BUFFD0 U98 ( .I(n114), .Z(n113) );
  BUFFD0 U99 ( .I(n115), .Z(n114) );
  BUFFD0 U100 ( .I(n116), .Z(n115) );
  BUFFD0 U101 ( .I(n117), .Z(n116) );
  BUFFD0 U102 ( .I(n118), .Z(n117) );
  BUFFD0 U103 ( .I(n119), .Z(n118) );
  BUFFD0 U104 ( .I(n120), .Z(n119) );
  BUFFD0 U105 ( .I(n121), .Z(n120) );
  BUFFD0 U106 ( .I(n122), .Z(n121) );
  BUFFD0 U107 ( .I(n123), .Z(n122) );
  BUFFD0 U108 ( .I(n124), .Z(n123) );
  BUFFD0 U109 ( .I(n125), .Z(n124) );
  BUFFD0 U110 ( .I(n126), .Z(n125) );
  BUFFD0 U111 ( .I(n127), .Z(n126) );
  BUFFD0 U112 ( .I(n128), .Z(n127) );
  BUFFD0 U113 ( .I(n129), .Z(n128) );
  BUFFD0 U114 ( .I(n130), .Z(n129) );
  BUFFD0 U115 ( .I(n131), .Z(n130) );
  BUFFD0 U116 ( .I(n132), .Z(n131) );
  BUFFD0 U117 ( .I(n133), .Z(n132) );
  BUFFD0 U118 ( .I(n134), .Z(n133) );
  BUFFD0 U119 ( .I(n135), .Z(n134) );
  BUFFD0 U120 ( .I(n136), .Z(n135) );
  BUFFD0 U121 ( .I(n137), .Z(n136) );
  BUFFD0 U122 ( .I(n138), .Z(n137) );
  BUFFD0 U123 ( .I(n139), .Z(n138) );
  BUFFD0 U124 ( .I(n140), .Z(n139) );
  BUFFD0 U125 ( .I(n141), .Z(n140) );
  BUFFD0 U126 ( .I(n142), .Z(n141) );
  BUFFD0 U127 ( .I(DataOr[30]), .Z(n142) );
  BUFFD0 U128 ( .I(n144), .Z(n143) );
  BUFFD0 U129 ( .I(n145), .Z(n144) );
  BUFFD0 U130 ( .I(n146), .Z(n145) );
  BUFFD0 U131 ( .I(n147), .Z(n146) );
  BUFFD0 U132 ( .I(n148), .Z(n147) );
  BUFFD0 U133 ( .I(n149), .Z(n148) );
  BUFFD0 U134 ( .I(n150), .Z(n149) );
  BUFFD0 U135 ( .I(n151), .Z(n150) );
  BUFFD0 U136 ( .I(n152), .Z(n151) );
  BUFFD0 U137 ( .I(n153), .Z(n152) );
  BUFFD0 U138 ( .I(n154), .Z(n153) );
  BUFFD0 U139 ( .I(n155), .Z(n154) );
  BUFFD0 U140 ( .I(n156), .Z(n155) );
  BUFFD0 U141 ( .I(n157), .Z(n156) );
  BUFFD0 U142 ( .I(n158), .Z(n157) );
  BUFFD0 U143 ( .I(n159), .Z(n158) );
  BUFFD0 U144 ( .I(n160), .Z(n159) );
  BUFFD0 U145 ( .I(n161), .Z(n160) );
  BUFFD0 U146 ( .I(n162), .Z(n161) );
  BUFFD0 U147 ( .I(n163), .Z(n162) );
  BUFFD0 U148 ( .I(n164), .Z(n163) );
  BUFFD0 U149 ( .I(n165), .Z(n164) );
  BUFFD0 U150 ( .I(n166), .Z(n165) );
  BUFFD0 U151 ( .I(n167), .Z(n166) );
  BUFFD0 U152 ( .I(n168), .Z(n167) );
  BUFFD0 U153 ( .I(n169), .Z(n168) );
  BUFFD0 U154 ( .I(n170), .Z(n169) );
  BUFFD0 U155 ( .I(n171), .Z(n170) );
  BUFFD0 U156 ( .I(n172), .Z(n171) );
  BUFFD0 U157 ( .I(n173), .Z(n172) );
  BUFFD0 U158 ( .I(n174), .Z(n173) );
  BUFFD0 U159 ( .I(n175), .Z(n174) );
  BUFFD0 U160 ( .I(n176), .Z(n175) );
  BUFFD0 U161 ( .I(n177), .Z(n176) );
  BUFFD0 U162 ( .I(n178), .Z(n177) );
  BUFFD0 U163 ( .I(n179), .Z(n178) );
  BUFFD0 U164 ( .I(n180), .Z(n179) );
  BUFFD0 U165 ( .I(n181), .Z(n180) );
  BUFFD0 U166 ( .I(n182), .Z(n181) );
  BUFFD0 U167 ( .I(n183), .Z(n182) );
  BUFFD0 U168 ( .I(n184), .Z(n183) );
  BUFFD0 U169 ( .I(n185), .Z(n184) );
  BUFFD0 U170 ( .I(n186), .Z(n185) );
  BUFFD0 U171 ( .I(n187), .Z(n186) );
  BUFFD0 U172 ( .I(n188), .Z(n187) );
  BUFFD0 U173 ( .I(n189), .Z(n188) );
  BUFFD0 U174 ( .I(n190), .Z(n189) );
  BUFFD0 U175 ( .I(n191), .Z(n190) );
  BUFFD0 U176 ( .I(n192), .Z(n191) );
  BUFFD0 U177 ( .I(n193), .Z(n192) );
  BUFFD0 U178 ( .I(n194), .Z(n193) );
  BUFFD0 U179 ( .I(n195), .Z(n194) );
  BUFFD0 U180 ( .I(n196), .Z(n195) );
  BUFFD0 U181 ( .I(DataOr[29]), .Z(n196) );
  BUFFD0 U182 ( .I(n198), .Z(n197) );
  BUFFD0 U183 ( .I(n199), .Z(n198) );
  BUFFD0 U184 ( .I(n200), .Z(n199) );
  BUFFD0 U185 ( .I(n201), .Z(n200) );
  BUFFD0 U186 ( .I(n202), .Z(n201) );
  BUFFD0 U187 ( .I(n203), .Z(n202) );
  BUFFD0 U188 ( .I(n204), .Z(n203) );
  BUFFD0 U189 ( .I(n205), .Z(n204) );
  BUFFD0 U190 ( .I(n206), .Z(n205) );
  BUFFD0 U191 ( .I(n207), .Z(n206) );
  BUFFD0 U192 ( .I(n208), .Z(n207) );
  BUFFD0 U193 ( .I(n209), .Z(n208) );
  BUFFD0 U194 ( .I(n210), .Z(n209) );
  BUFFD0 U195 ( .I(n211), .Z(n210) );
  BUFFD0 U196 ( .I(n212), .Z(n211) );
  BUFFD0 U197 ( .I(n213), .Z(n212) );
  BUFFD0 U198 ( .I(n214), .Z(n213) );
  BUFFD0 U199 ( .I(n215), .Z(n214) );
  BUFFD0 U200 ( .I(n216), .Z(n215) );
  BUFFD0 U201 ( .I(n217), .Z(n216) );
  BUFFD0 U202 ( .I(n218), .Z(n217) );
  BUFFD0 U203 ( .I(n219), .Z(n218) );
  BUFFD0 U204 ( .I(n220), .Z(n219) );
  BUFFD0 U205 ( .I(n221), .Z(n220) );
  BUFFD0 U206 ( .I(n222), .Z(n221) );
  BUFFD0 U207 ( .I(n223), .Z(n222) );
  BUFFD0 U208 ( .I(n224), .Z(n223) );
  BUFFD0 U209 ( .I(n225), .Z(n224) );
  BUFFD0 U210 ( .I(n226), .Z(n225) );
  BUFFD0 U211 ( .I(n227), .Z(n226) );
  BUFFD0 U212 ( .I(n228), .Z(n227) );
  BUFFD0 U213 ( .I(n229), .Z(n228) );
  BUFFD0 U214 ( .I(n230), .Z(n229) );
  BUFFD0 U215 ( .I(n231), .Z(n230) );
  BUFFD0 U216 ( .I(n232), .Z(n231) );
  BUFFD0 U217 ( .I(n233), .Z(n232) );
  BUFFD0 U218 ( .I(n234), .Z(n233) );
  BUFFD0 U219 ( .I(n235), .Z(n234) );
  BUFFD0 U220 ( .I(n236), .Z(n235) );
  BUFFD0 U221 ( .I(n237), .Z(n236) );
  BUFFD0 U222 ( .I(n238), .Z(n237) );
  BUFFD0 U223 ( .I(n239), .Z(n238) );
  BUFFD0 U224 ( .I(n240), .Z(n239) );
  BUFFD0 U225 ( .I(n241), .Z(n240) );
  BUFFD0 U226 ( .I(n242), .Z(n241) );
  BUFFD0 U227 ( .I(n243), .Z(n242) );
  BUFFD0 U228 ( .I(n244), .Z(n243) );
  BUFFD0 U229 ( .I(n245), .Z(n244) );
  BUFFD0 U230 ( .I(n246), .Z(n245) );
  BUFFD0 U231 ( .I(n247), .Z(n246) );
  BUFFD0 U232 ( .I(n248), .Z(n247) );
  BUFFD0 U233 ( .I(n249), .Z(n248) );
  BUFFD0 U234 ( .I(n250), .Z(n249) );
  BUFFD0 U235 ( .I(DataOr[28]), .Z(n250) );
  BUFFD0 U236 ( .I(n252), .Z(n251) );
  BUFFD0 U237 ( .I(n253), .Z(n252) );
  BUFFD0 U238 ( .I(n254), .Z(n253) );
  BUFFD0 U239 ( .I(n255), .Z(n254) );
  BUFFD0 U240 ( .I(n256), .Z(n255) );
  BUFFD0 U241 ( .I(n257), .Z(n256) );
  BUFFD0 U242 ( .I(n258), .Z(n257) );
  BUFFD0 U243 ( .I(n259), .Z(n258) );
  BUFFD0 U244 ( .I(n260), .Z(n259) );
  BUFFD0 U245 ( .I(n261), .Z(n260) );
  BUFFD0 U246 ( .I(n262), .Z(n261) );
  BUFFD0 U247 ( .I(n263), .Z(n262) );
  BUFFD0 U248 ( .I(n264), .Z(n263) );
  BUFFD0 U249 ( .I(n265), .Z(n264) );
  BUFFD0 U250 ( .I(n266), .Z(n265) );
  BUFFD0 U251 ( .I(n267), .Z(n266) );
  BUFFD0 U252 ( .I(n268), .Z(n267) );
  BUFFD0 U253 ( .I(n269), .Z(n268) );
  BUFFD0 U254 ( .I(n270), .Z(n269) );
  BUFFD0 U255 ( .I(n271), .Z(n270) );
  BUFFD0 U256 ( .I(n272), .Z(n271) );
  BUFFD0 U257 ( .I(n273), .Z(n272) );
  BUFFD0 U258 ( .I(n274), .Z(n273) );
  BUFFD0 U259 ( .I(n275), .Z(n274) );
  BUFFD0 U260 ( .I(n276), .Z(n275) );
  BUFFD0 U261 ( .I(n277), .Z(n276) );
  BUFFD0 U262 ( .I(n278), .Z(n277) );
  BUFFD0 U263 ( .I(n279), .Z(n278) );
  BUFFD0 U264 ( .I(n280), .Z(n279) );
  BUFFD0 U265 ( .I(n281), .Z(n280) );
  BUFFD0 U266 ( .I(n282), .Z(n281) );
  BUFFD0 U267 ( .I(n283), .Z(n282) );
  BUFFD0 U268 ( .I(n284), .Z(n283) );
  BUFFD0 U269 ( .I(n285), .Z(n284) );
  BUFFD0 U270 ( .I(n286), .Z(n285) );
  BUFFD0 U271 ( .I(n287), .Z(n286) );
  BUFFD0 U272 ( .I(n288), .Z(n287) );
  BUFFD0 U273 ( .I(n289), .Z(n288) );
  BUFFD0 U274 ( .I(n290), .Z(n289) );
  BUFFD0 U275 ( .I(n291), .Z(n290) );
  BUFFD0 U276 ( .I(n292), .Z(n291) );
  BUFFD0 U277 ( .I(n293), .Z(n292) );
  BUFFD0 U278 ( .I(n294), .Z(n293) );
  BUFFD0 U279 ( .I(n295), .Z(n294) );
  BUFFD0 U280 ( .I(n296), .Z(n295) );
  BUFFD0 U281 ( .I(n297), .Z(n296) );
  BUFFD0 U282 ( .I(n298), .Z(n297) );
  BUFFD0 U283 ( .I(n299), .Z(n298) );
  BUFFD0 U284 ( .I(n300), .Z(n299) );
  BUFFD0 U285 ( .I(n301), .Z(n300) );
  BUFFD0 U286 ( .I(n302), .Z(n301) );
  BUFFD0 U287 ( .I(n303), .Z(n302) );
  BUFFD0 U288 ( .I(n304), .Z(n303) );
  BUFFD0 U289 ( .I(DataOr[27]), .Z(n304) );
  BUFFD0 U290 ( .I(n306), .Z(n305) );
  BUFFD0 U291 ( .I(n307), .Z(n306) );
  BUFFD0 U292 ( .I(n308), .Z(n307) );
  BUFFD0 U293 ( .I(n309), .Z(n308) );
  BUFFD0 U294 ( .I(n310), .Z(n309) );
  BUFFD0 U295 ( .I(n311), .Z(n310) );
  BUFFD0 U296 ( .I(n312), .Z(n311) );
  BUFFD0 U297 ( .I(n313), .Z(n312) );
  BUFFD0 U298 ( .I(n314), .Z(n313) );
  BUFFD0 U299 ( .I(n315), .Z(n314) );
  BUFFD0 U300 ( .I(n316), .Z(n315) );
  BUFFD0 U301 ( .I(n317), .Z(n316) );
  BUFFD0 U302 ( .I(n318), .Z(n317) );
  BUFFD0 U303 ( .I(n319), .Z(n318) );
  BUFFD0 U304 ( .I(n320), .Z(n319) );
  BUFFD0 U305 ( .I(n321), .Z(n320) );
  BUFFD0 U306 ( .I(n322), .Z(n321) );
  BUFFD0 U307 ( .I(n323), .Z(n322) );
  BUFFD0 U308 ( .I(n324), .Z(n323) );
  BUFFD0 U309 ( .I(n325), .Z(n324) );
  BUFFD0 U310 ( .I(n326), .Z(n325) );
  BUFFD0 U311 ( .I(n327), .Z(n326) );
  BUFFD0 U312 ( .I(n328), .Z(n327) );
  BUFFD0 U313 ( .I(n329), .Z(n328) );
  BUFFD0 U314 ( .I(n330), .Z(n329) );
  BUFFD0 U315 ( .I(n331), .Z(n330) );
  BUFFD0 U316 ( .I(n332), .Z(n331) );
  BUFFD0 U317 ( .I(n333), .Z(n332) );
  BUFFD0 U318 ( .I(n334), .Z(n333) );
  BUFFD0 U319 ( .I(n335), .Z(n334) );
  BUFFD0 U320 ( .I(n336), .Z(n335) );
  BUFFD0 U321 ( .I(n337), .Z(n336) );
  BUFFD0 U322 ( .I(n338), .Z(n337) );
  BUFFD0 U323 ( .I(n339), .Z(n338) );
  BUFFD0 U324 ( .I(n340), .Z(n339) );
  BUFFD0 U325 ( .I(n341), .Z(n340) );
  BUFFD0 U326 ( .I(n342), .Z(n341) );
  BUFFD0 U327 ( .I(n343), .Z(n342) );
  BUFFD0 U328 ( .I(n344), .Z(n343) );
  BUFFD0 U329 ( .I(n345), .Z(n344) );
  BUFFD0 U330 ( .I(n346), .Z(n345) );
  BUFFD0 U331 ( .I(n347), .Z(n346) );
  BUFFD0 U332 ( .I(n348), .Z(n347) );
  BUFFD0 U333 ( .I(n349), .Z(n348) );
  BUFFD0 U334 ( .I(n350), .Z(n349) );
  BUFFD0 U335 ( .I(n351), .Z(n350) );
  BUFFD0 U336 ( .I(n352), .Z(n351) );
  BUFFD0 U337 ( .I(n353), .Z(n352) );
  BUFFD0 U338 ( .I(n354), .Z(n353) );
  BUFFD0 U339 ( .I(n355), .Z(n354) );
  BUFFD0 U340 ( .I(n356), .Z(n355) );
  BUFFD0 U341 ( .I(n357), .Z(n356) );
  BUFFD0 U342 ( .I(n358), .Z(n357) );
  BUFFD0 U343 ( .I(DataOr[26]), .Z(n358) );
  BUFFD0 U344 ( .I(n360), .Z(n359) );
  BUFFD0 U345 ( .I(n361), .Z(n360) );
  BUFFD0 U346 ( .I(n362), .Z(n361) );
  BUFFD0 U347 ( .I(n363), .Z(n362) );
  BUFFD0 U348 ( .I(n364), .Z(n363) );
  BUFFD0 U349 ( .I(n365), .Z(n364) );
  BUFFD0 U350 ( .I(n366), .Z(n365) );
  BUFFD0 U351 ( .I(n367), .Z(n366) );
  BUFFD0 U352 ( .I(n368), .Z(n367) );
  BUFFD0 U353 ( .I(n369), .Z(n368) );
  BUFFD0 U354 ( .I(n370), .Z(n369) );
  BUFFD0 U355 ( .I(n371), .Z(n370) );
  BUFFD0 U356 ( .I(n372), .Z(n371) );
  BUFFD0 U357 ( .I(n373), .Z(n372) );
  BUFFD0 U358 ( .I(n374), .Z(n373) );
  BUFFD0 U359 ( .I(n375), .Z(n374) );
  BUFFD0 U360 ( .I(n376), .Z(n375) );
  BUFFD0 U361 ( .I(n377), .Z(n376) );
  BUFFD0 U362 ( .I(n378), .Z(n377) );
  BUFFD0 U363 ( .I(n379), .Z(n378) );
  BUFFD0 U364 ( .I(n380), .Z(n379) );
  BUFFD0 U365 ( .I(n381), .Z(n380) );
  BUFFD0 U366 ( .I(n382), .Z(n381) );
  BUFFD0 U367 ( .I(n383), .Z(n382) );
  BUFFD0 U368 ( .I(n384), .Z(n383) );
  BUFFD0 U369 ( .I(n385), .Z(n384) );
  BUFFD0 U370 ( .I(n386), .Z(n385) );
  BUFFD0 U371 ( .I(n387), .Z(n386) );
  BUFFD0 U372 ( .I(n388), .Z(n387) );
  BUFFD0 U373 ( .I(n389), .Z(n388) );
  BUFFD0 U374 ( .I(n390), .Z(n389) );
  BUFFD0 U375 ( .I(n391), .Z(n390) );
  BUFFD0 U376 ( .I(n392), .Z(n391) );
  BUFFD0 U377 ( .I(n393), .Z(n392) );
  BUFFD0 U378 ( .I(n394), .Z(n393) );
  BUFFD0 U379 ( .I(n395), .Z(n394) );
  BUFFD0 U380 ( .I(n396), .Z(n395) );
  BUFFD0 U381 ( .I(n397), .Z(n396) );
  BUFFD0 U382 ( .I(n398), .Z(n397) );
  BUFFD0 U383 ( .I(n399), .Z(n398) );
  BUFFD0 U384 ( .I(n400), .Z(n399) );
  BUFFD0 U385 ( .I(n401), .Z(n400) );
  BUFFD0 U386 ( .I(n402), .Z(n401) );
  BUFFD0 U387 ( .I(n403), .Z(n402) );
  BUFFD0 U388 ( .I(n404), .Z(n403) );
  BUFFD0 U389 ( .I(n405), .Z(n404) );
  BUFFD0 U390 ( .I(n406), .Z(n405) );
  BUFFD0 U391 ( .I(n407), .Z(n406) );
  BUFFD0 U392 ( .I(n408), .Z(n407) );
  BUFFD0 U393 ( .I(n409), .Z(n408) );
  BUFFD0 U394 ( .I(n410), .Z(n409) );
  BUFFD0 U395 ( .I(n411), .Z(n410) );
  BUFFD0 U396 ( .I(n412), .Z(n411) );
  BUFFD0 U397 ( .I(DataOr[25]), .Z(n412) );
  BUFFD0 U398 ( .I(n414), .Z(n413) );
  BUFFD0 U399 ( .I(n415), .Z(n414) );
  BUFFD0 U400 ( .I(n416), .Z(n415) );
  BUFFD0 U401 ( .I(n417), .Z(n416) );
  BUFFD0 U402 ( .I(n418), .Z(n417) );
  BUFFD0 U403 ( .I(n419), .Z(n418) );
  BUFFD0 U404 ( .I(n420), .Z(n419) );
  BUFFD0 U405 ( .I(n421), .Z(n420) );
  BUFFD0 U406 ( .I(n422), .Z(n421) );
  BUFFD0 U407 ( .I(n423), .Z(n422) );
  BUFFD0 U408 ( .I(n424), .Z(n423) );
  BUFFD0 U409 ( .I(n425), .Z(n424) );
  BUFFD0 U410 ( .I(n426), .Z(n425) );
  BUFFD0 U411 ( .I(n427), .Z(n426) );
  BUFFD0 U412 ( .I(n428), .Z(n427) );
  BUFFD0 U413 ( .I(n429), .Z(n428) );
  BUFFD0 U414 ( .I(n430), .Z(n429) );
  BUFFD0 U415 ( .I(n431), .Z(n430) );
  BUFFD0 U416 ( .I(n432), .Z(n431) );
  BUFFD0 U417 ( .I(n433), .Z(n432) );
  BUFFD0 U418 ( .I(n434), .Z(n433) );
  BUFFD0 U419 ( .I(n435), .Z(n434) );
  BUFFD0 U420 ( .I(n436), .Z(n435) );
  BUFFD0 U421 ( .I(n437), .Z(n436) );
  BUFFD0 U422 ( .I(n438), .Z(n437) );
  BUFFD0 U423 ( .I(n439), .Z(n438) );
  BUFFD0 U424 ( .I(n440), .Z(n439) );
  BUFFD0 U425 ( .I(n441), .Z(n440) );
  BUFFD0 U426 ( .I(n442), .Z(n441) );
  BUFFD0 U427 ( .I(n443), .Z(n442) );
  BUFFD0 U428 ( .I(n444), .Z(n443) );
  BUFFD0 U429 ( .I(n445), .Z(n444) );
  BUFFD0 U430 ( .I(n446), .Z(n445) );
  BUFFD0 U431 ( .I(n447), .Z(n446) );
  BUFFD0 U432 ( .I(n448), .Z(n447) );
  BUFFD0 U433 ( .I(n449), .Z(n448) );
  BUFFD0 U434 ( .I(n450), .Z(n449) );
  BUFFD0 U435 ( .I(n451), .Z(n450) );
  BUFFD0 U436 ( .I(n452), .Z(n451) );
  BUFFD0 U437 ( .I(n453), .Z(n452) );
  BUFFD0 U438 ( .I(n454), .Z(n453) );
  BUFFD0 U439 ( .I(n455), .Z(n454) );
  BUFFD0 U440 ( .I(n456), .Z(n455) );
  BUFFD0 U441 ( .I(n457), .Z(n456) );
  BUFFD0 U442 ( .I(n458), .Z(n457) );
  BUFFD0 U443 ( .I(n459), .Z(n458) );
  BUFFD0 U444 ( .I(n460), .Z(n459) );
  BUFFD0 U445 ( .I(n461), .Z(n460) );
  BUFFD0 U446 ( .I(n462), .Z(n461) );
  BUFFD0 U447 ( .I(n463), .Z(n462) );
  BUFFD0 U448 ( .I(n464), .Z(n463) );
  BUFFD0 U449 ( .I(n465), .Z(n464) );
  BUFFD0 U450 ( .I(n466), .Z(n465) );
  BUFFD0 U451 ( .I(DataOr[24]), .Z(n466) );
  BUFFD0 U452 ( .I(n468), .Z(n467) );
  BUFFD0 U453 ( .I(n469), .Z(n468) );
  BUFFD0 U454 ( .I(n470), .Z(n469) );
  BUFFD0 U455 ( .I(n471), .Z(n470) );
  BUFFD0 U456 ( .I(n472), .Z(n471) );
  BUFFD0 U457 ( .I(n473), .Z(n472) );
  BUFFD0 U458 ( .I(n474), .Z(n473) );
  BUFFD0 U459 ( .I(n475), .Z(n474) );
  BUFFD0 U460 ( .I(n476), .Z(n475) );
  BUFFD0 U461 ( .I(n477), .Z(n476) );
  BUFFD0 U462 ( .I(n478), .Z(n477) );
  BUFFD0 U463 ( .I(n479), .Z(n478) );
  BUFFD0 U464 ( .I(n480), .Z(n479) );
  BUFFD0 U465 ( .I(n481), .Z(n480) );
  BUFFD0 U466 ( .I(n482), .Z(n481) );
  BUFFD0 U467 ( .I(n483), .Z(n482) );
  BUFFD0 U468 ( .I(n484), .Z(n483) );
  BUFFD0 U469 ( .I(n485), .Z(n484) );
  BUFFD0 U470 ( .I(n486), .Z(n485) );
  BUFFD0 U471 ( .I(n487), .Z(n486) );
  BUFFD0 U472 ( .I(n488), .Z(n487) );
  BUFFD0 U473 ( .I(n489), .Z(n488) );
  BUFFD0 U474 ( .I(n490), .Z(n489) );
  BUFFD0 U475 ( .I(n491), .Z(n490) );
  BUFFD0 U476 ( .I(n492), .Z(n491) );
  BUFFD0 U477 ( .I(n493), .Z(n492) );
  BUFFD0 U478 ( .I(n494), .Z(n493) );
  BUFFD0 U479 ( .I(n495), .Z(n494) );
  BUFFD0 U480 ( .I(n496), .Z(n495) );
  BUFFD0 U481 ( .I(n497), .Z(n496) );
  BUFFD0 U482 ( .I(n498), .Z(n497) );
  BUFFD0 U483 ( .I(n499), .Z(n498) );
  BUFFD0 U484 ( .I(n500), .Z(n499) );
  BUFFD0 U485 ( .I(n501), .Z(n500) );
  BUFFD0 U486 ( .I(n502), .Z(n501) );
  BUFFD0 U487 ( .I(n503), .Z(n502) );
  BUFFD0 U488 ( .I(n504), .Z(n503) );
  BUFFD0 U489 ( .I(n505), .Z(n504) );
  BUFFD0 U490 ( .I(n506), .Z(n505) );
  BUFFD0 U491 ( .I(n507), .Z(n506) );
  BUFFD0 U492 ( .I(n508), .Z(n507) );
  BUFFD0 U493 ( .I(n509), .Z(n508) );
  BUFFD0 U494 ( .I(n510), .Z(n509) );
  BUFFD0 U495 ( .I(n511), .Z(n510) );
  BUFFD0 U496 ( .I(n512), .Z(n511) );
  BUFFD0 U497 ( .I(n513), .Z(n512) );
  BUFFD0 U498 ( .I(n514), .Z(n513) );
  BUFFD0 U499 ( .I(n515), .Z(n514) );
  BUFFD0 U500 ( .I(n516), .Z(n515) );
  BUFFD0 U501 ( .I(n517), .Z(n516) );
  BUFFD0 U502 ( .I(n518), .Z(n517) );
  BUFFD0 U503 ( .I(n519), .Z(n518) );
  BUFFD0 U504 ( .I(n520), .Z(n519) );
  BUFFD0 U505 ( .I(DataOr[23]), .Z(n520) );
  BUFFD0 U506 ( .I(n522), .Z(n521) );
  BUFFD0 U507 ( .I(n523), .Z(n522) );
  BUFFD0 U508 ( .I(n524), .Z(n523) );
  BUFFD0 U509 ( .I(n525), .Z(n524) );
  BUFFD0 U510 ( .I(n526), .Z(n525) );
  BUFFD0 U511 ( .I(n527), .Z(n526) );
  BUFFD0 U512 ( .I(n528), .Z(n527) );
  BUFFD0 U513 ( .I(n529), .Z(n528) );
  BUFFD0 U514 ( .I(n530), .Z(n529) );
  BUFFD0 U515 ( .I(n531), .Z(n530) );
  BUFFD0 U516 ( .I(n532), .Z(n531) );
  BUFFD0 U517 ( .I(n533), .Z(n532) );
  BUFFD0 U518 ( .I(n534), .Z(n533) );
  BUFFD0 U519 ( .I(n535), .Z(n534) );
  BUFFD0 U520 ( .I(n536), .Z(n535) );
  BUFFD0 U521 ( .I(n537), .Z(n536) );
  BUFFD0 U522 ( .I(n538), .Z(n537) );
  BUFFD0 U523 ( .I(n539), .Z(n538) );
  BUFFD0 U524 ( .I(n540), .Z(n539) );
  BUFFD0 U525 ( .I(n541), .Z(n540) );
  BUFFD0 U526 ( .I(n542), .Z(n541) );
  BUFFD0 U527 ( .I(n543), .Z(n542) );
  BUFFD0 U528 ( .I(n544), .Z(n543) );
  BUFFD0 U529 ( .I(n545), .Z(n544) );
  BUFFD0 U530 ( .I(n546), .Z(n545) );
  BUFFD0 U531 ( .I(n547), .Z(n546) );
  BUFFD0 U532 ( .I(n548), .Z(n547) );
  BUFFD0 U533 ( .I(n549), .Z(n548) );
  BUFFD0 U534 ( .I(n550), .Z(n549) );
  BUFFD0 U535 ( .I(n551), .Z(n550) );
  BUFFD0 U536 ( .I(n552), .Z(n551) );
  BUFFD0 U537 ( .I(n553), .Z(n552) );
  BUFFD0 U538 ( .I(n554), .Z(n553) );
  BUFFD0 U539 ( .I(n555), .Z(n554) );
  BUFFD0 U540 ( .I(n556), .Z(n555) );
  BUFFD0 U541 ( .I(n557), .Z(n556) );
  BUFFD0 U542 ( .I(n558), .Z(n557) );
  BUFFD0 U543 ( .I(n559), .Z(n558) );
  BUFFD0 U544 ( .I(n560), .Z(n559) );
  BUFFD0 U545 ( .I(n561), .Z(n560) );
  BUFFD0 U546 ( .I(n562), .Z(n561) );
  BUFFD0 U547 ( .I(n563), .Z(n562) );
  BUFFD0 U548 ( .I(n564), .Z(n563) );
  BUFFD0 U549 ( .I(n565), .Z(n564) );
  BUFFD0 U550 ( .I(n566), .Z(n565) );
  BUFFD0 U551 ( .I(n567), .Z(n566) );
  BUFFD0 U552 ( .I(n568), .Z(n567) );
  BUFFD0 U553 ( .I(n569), .Z(n568) );
  BUFFD0 U554 ( .I(n570), .Z(n569) );
  BUFFD0 U555 ( .I(n571), .Z(n570) );
  BUFFD0 U556 ( .I(n572), .Z(n571) );
  BUFFD0 U557 ( .I(n573), .Z(n572) );
  BUFFD0 U558 ( .I(n574), .Z(n573) );
  BUFFD0 U559 ( .I(DataOr[22]), .Z(n574) );
  BUFFD0 U560 ( .I(n576), .Z(n575) );
  BUFFD0 U561 ( .I(n577), .Z(n576) );
  BUFFD0 U562 ( .I(n578), .Z(n577) );
  BUFFD0 U563 ( .I(n579), .Z(n578) );
  BUFFD0 U564 ( .I(n580), .Z(n579) );
  BUFFD0 U565 ( .I(n581), .Z(n580) );
  BUFFD0 U566 ( .I(n582), .Z(n581) );
  BUFFD0 U567 ( .I(n583), .Z(n582) );
  BUFFD0 U568 ( .I(n584), .Z(n583) );
  BUFFD0 U569 ( .I(n585), .Z(n584) );
  BUFFD0 U570 ( .I(n586), .Z(n585) );
  BUFFD0 U571 ( .I(n587), .Z(n586) );
  BUFFD0 U572 ( .I(n588), .Z(n587) );
  BUFFD0 U573 ( .I(n589), .Z(n588) );
  BUFFD0 U574 ( .I(n590), .Z(n589) );
  BUFFD0 U575 ( .I(n591), .Z(n590) );
  BUFFD0 U576 ( .I(n592), .Z(n591) );
  BUFFD0 U577 ( .I(n593), .Z(n592) );
  BUFFD0 U578 ( .I(n594), .Z(n593) );
  BUFFD0 U579 ( .I(n595), .Z(n594) );
  BUFFD0 U580 ( .I(n596), .Z(n595) );
  BUFFD0 U581 ( .I(n597), .Z(n596) );
  BUFFD0 U582 ( .I(n598), .Z(n597) );
  BUFFD0 U583 ( .I(n599), .Z(n598) );
  BUFFD0 U584 ( .I(n600), .Z(n599) );
  BUFFD0 U585 ( .I(n601), .Z(n600) );
  BUFFD0 U586 ( .I(n602), .Z(n601) );
  BUFFD0 U587 ( .I(n603), .Z(n602) );
  BUFFD0 U588 ( .I(n604), .Z(n603) );
  BUFFD0 U589 ( .I(n605), .Z(n604) );
  BUFFD0 U590 ( .I(n606), .Z(n605) );
  BUFFD0 U591 ( .I(n607), .Z(n606) );
  BUFFD0 U592 ( .I(n608), .Z(n607) );
  BUFFD0 U593 ( .I(n609), .Z(n608) );
  BUFFD0 U594 ( .I(n610), .Z(n609) );
  BUFFD0 U595 ( .I(n611), .Z(n610) );
  BUFFD0 U596 ( .I(n612), .Z(n611) );
  BUFFD0 U597 ( .I(n613), .Z(n612) );
  BUFFD0 U598 ( .I(n614), .Z(n613) );
  BUFFD0 U599 ( .I(n615), .Z(n614) );
  BUFFD0 U600 ( .I(n616), .Z(n615) );
  BUFFD0 U601 ( .I(n617), .Z(n616) );
  BUFFD0 U602 ( .I(n618), .Z(n617) );
  BUFFD0 U603 ( .I(n619), .Z(n618) );
  BUFFD0 U604 ( .I(n620), .Z(n619) );
  BUFFD0 U605 ( .I(n621), .Z(n620) );
  BUFFD0 U606 ( .I(n622), .Z(n621) );
  BUFFD0 U607 ( .I(n623), .Z(n622) );
  BUFFD0 U608 ( .I(n624), .Z(n623) );
  BUFFD0 U609 ( .I(n625), .Z(n624) );
  BUFFD0 U610 ( .I(n626), .Z(n625) );
  BUFFD0 U611 ( .I(n627), .Z(n626) );
  BUFFD0 U612 ( .I(n628), .Z(n627) );
  BUFFD0 U613 ( .I(DataOr[21]), .Z(n628) );
  BUFFD0 U614 ( .I(n630), .Z(n629) );
  BUFFD0 U615 ( .I(n631), .Z(n630) );
  BUFFD0 U616 ( .I(n632), .Z(n631) );
  BUFFD0 U617 ( .I(n633), .Z(n632) );
  BUFFD0 U618 ( .I(n634), .Z(n633) );
  BUFFD0 U619 ( .I(n635), .Z(n634) );
  BUFFD0 U620 ( .I(n636), .Z(n635) );
  BUFFD0 U621 ( .I(n637), .Z(n636) );
  BUFFD0 U622 ( .I(n638), .Z(n637) );
  BUFFD0 U623 ( .I(n639), .Z(n638) );
  BUFFD0 U624 ( .I(n640), .Z(n639) );
  BUFFD0 U625 ( .I(n641), .Z(n640) );
  BUFFD0 U626 ( .I(n642), .Z(n641) );
  BUFFD0 U627 ( .I(n643), .Z(n642) );
  BUFFD0 U628 ( .I(n644), .Z(n643) );
  BUFFD0 U629 ( .I(n645), .Z(n644) );
  BUFFD0 U630 ( .I(n646), .Z(n645) );
  BUFFD0 U631 ( .I(n647), .Z(n646) );
  BUFFD0 U632 ( .I(n648), .Z(n647) );
  BUFFD0 U633 ( .I(n649), .Z(n648) );
  BUFFD0 U634 ( .I(n650), .Z(n649) );
  BUFFD0 U635 ( .I(n651), .Z(n650) );
  BUFFD0 U636 ( .I(n652), .Z(n651) );
  BUFFD0 U637 ( .I(n653), .Z(n652) );
  BUFFD0 U638 ( .I(n654), .Z(n653) );
  BUFFD0 U639 ( .I(n655), .Z(n654) );
  BUFFD0 U640 ( .I(n656), .Z(n655) );
  BUFFD0 U641 ( .I(n657), .Z(n656) );
  BUFFD0 U642 ( .I(n658), .Z(n657) );
  BUFFD0 U643 ( .I(n659), .Z(n658) );
  BUFFD0 U644 ( .I(n660), .Z(n659) );
  BUFFD0 U645 ( .I(n661), .Z(n660) );
  BUFFD0 U646 ( .I(n662), .Z(n661) );
  BUFFD0 U647 ( .I(n663), .Z(n662) );
  BUFFD0 U648 ( .I(n664), .Z(n663) );
  BUFFD0 U649 ( .I(n665), .Z(n664) );
  BUFFD0 U650 ( .I(n666), .Z(n665) );
  BUFFD0 U651 ( .I(n667), .Z(n666) );
  BUFFD0 U652 ( .I(n668), .Z(n667) );
  BUFFD0 U653 ( .I(n669), .Z(n668) );
  BUFFD0 U654 ( .I(n670), .Z(n669) );
  BUFFD0 U655 ( .I(n671), .Z(n670) );
  BUFFD0 U656 ( .I(n672), .Z(n671) );
  BUFFD0 U657 ( .I(n673), .Z(n672) );
  BUFFD0 U658 ( .I(n674), .Z(n673) );
  BUFFD0 U659 ( .I(n675), .Z(n674) );
  BUFFD0 U660 ( .I(n676), .Z(n675) );
  BUFFD0 U661 ( .I(n677), .Z(n676) );
  BUFFD0 U662 ( .I(n678), .Z(n677) );
  BUFFD0 U663 ( .I(n679), .Z(n678) );
  BUFFD0 U664 ( .I(n680), .Z(n679) );
  BUFFD0 U665 ( .I(n681), .Z(n680) );
  BUFFD0 U666 ( .I(n682), .Z(n681) );
  BUFFD0 U667 ( .I(DataOr[20]), .Z(n682) );
  BUFFD0 U668 ( .I(n684), .Z(n683) );
  BUFFD0 U669 ( .I(n685), .Z(n684) );
  BUFFD0 U670 ( .I(n686), .Z(n685) );
  BUFFD0 U671 ( .I(n687), .Z(n686) );
  BUFFD0 U672 ( .I(n688), .Z(n687) );
  BUFFD0 U673 ( .I(n689), .Z(n688) );
  BUFFD0 U674 ( .I(n690), .Z(n689) );
  BUFFD0 U675 ( .I(n691), .Z(n690) );
  BUFFD0 U676 ( .I(n692), .Z(n691) );
  BUFFD0 U677 ( .I(n693), .Z(n692) );
  BUFFD0 U678 ( .I(n694), .Z(n693) );
  BUFFD0 U679 ( .I(n695), .Z(n694) );
  BUFFD0 U680 ( .I(n696), .Z(n695) );
  BUFFD0 U681 ( .I(n697), .Z(n696) );
  BUFFD0 U682 ( .I(n698), .Z(n697) );
  BUFFD0 U683 ( .I(n699), .Z(n698) );
  BUFFD0 U684 ( .I(n700), .Z(n699) );
  BUFFD0 U685 ( .I(n701), .Z(n700) );
  BUFFD0 U686 ( .I(n702), .Z(n701) );
  BUFFD0 U687 ( .I(n703), .Z(n702) );
  BUFFD0 U688 ( .I(n704), .Z(n703) );
  BUFFD0 U689 ( .I(n705), .Z(n704) );
  BUFFD0 U690 ( .I(n706), .Z(n705) );
  BUFFD0 U691 ( .I(n707), .Z(n706) );
  BUFFD0 U692 ( .I(n708), .Z(n707) );
  BUFFD0 U693 ( .I(n709), .Z(n708) );
  BUFFD0 U694 ( .I(n710), .Z(n709) );
  BUFFD0 U695 ( .I(n711), .Z(n710) );
  BUFFD0 U696 ( .I(n712), .Z(n711) );
  BUFFD0 U697 ( .I(n713), .Z(n712) );
  BUFFD0 U698 ( .I(n714), .Z(n713) );
  BUFFD0 U699 ( .I(n715), .Z(n714) );
  BUFFD0 U700 ( .I(n716), .Z(n715) );
  BUFFD0 U701 ( .I(n717), .Z(n716) );
  BUFFD0 U702 ( .I(n718), .Z(n717) );
  BUFFD0 U703 ( .I(n719), .Z(n718) );
  BUFFD0 U704 ( .I(n720), .Z(n719) );
  BUFFD0 U705 ( .I(n721), .Z(n720) );
  BUFFD0 U706 ( .I(n722), .Z(n721) );
  BUFFD0 U707 ( .I(n723), .Z(n722) );
  BUFFD0 U708 ( .I(n724), .Z(n723) );
  BUFFD0 U709 ( .I(n725), .Z(n724) );
  BUFFD0 U710 ( .I(n726), .Z(n725) );
  BUFFD0 U711 ( .I(n727), .Z(n726) );
  BUFFD0 U712 ( .I(n728), .Z(n727) );
  BUFFD0 U713 ( .I(n729), .Z(n728) );
  BUFFD0 U714 ( .I(n730), .Z(n729) );
  BUFFD0 U715 ( .I(n731), .Z(n730) );
  BUFFD0 U716 ( .I(n732), .Z(n731) );
  BUFFD0 U717 ( .I(n733), .Z(n732) );
  BUFFD0 U718 ( .I(n734), .Z(n733) );
  BUFFD0 U719 ( .I(n735), .Z(n734) );
  BUFFD0 U720 ( .I(n736), .Z(n735) );
  BUFFD0 U721 ( .I(DataOr[19]), .Z(n736) );
  BUFFD0 U722 ( .I(n738), .Z(n737) );
  BUFFD0 U723 ( .I(n739), .Z(n738) );
  BUFFD0 U724 ( .I(n740), .Z(n739) );
  BUFFD0 U725 ( .I(n741), .Z(n740) );
  BUFFD0 U726 ( .I(n742), .Z(n741) );
  BUFFD0 U727 ( .I(n743), .Z(n742) );
  BUFFD0 U728 ( .I(n744), .Z(n743) );
  BUFFD0 U729 ( .I(n745), .Z(n744) );
  BUFFD0 U730 ( .I(n746), .Z(n745) );
  BUFFD0 U731 ( .I(n747), .Z(n746) );
  BUFFD0 U732 ( .I(n748), .Z(n747) );
  BUFFD0 U733 ( .I(n749), .Z(n748) );
  BUFFD0 U734 ( .I(n750), .Z(n749) );
  BUFFD0 U735 ( .I(n751), .Z(n750) );
  BUFFD0 U736 ( .I(n752), .Z(n751) );
  BUFFD0 U737 ( .I(n753), .Z(n752) );
  BUFFD0 U738 ( .I(n754), .Z(n753) );
  BUFFD0 U739 ( .I(n755), .Z(n754) );
  BUFFD0 U740 ( .I(n756), .Z(n755) );
  BUFFD0 U741 ( .I(n757), .Z(n756) );
  BUFFD0 U742 ( .I(n758), .Z(n757) );
  BUFFD0 U743 ( .I(n759), .Z(n758) );
  BUFFD0 U744 ( .I(n760), .Z(n759) );
  BUFFD0 U745 ( .I(n761), .Z(n760) );
  BUFFD0 U746 ( .I(n762), .Z(n761) );
  BUFFD0 U747 ( .I(n763), .Z(n762) );
  BUFFD0 U748 ( .I(n764), .Z(n763) );
  BUFFD0 U749 ( .I(n765), .Z(n764) );
  BUFFD0 U750 ( .I(n766), .Z(n765) );
  BUFFD0 U751 ( .I(n767), .Z(n766) );
  BUFFD0 U752 ( .I(n768), .Z(n767) );
  BUFFD0 U753 ( .I(n769), .Z(n768) );
  BUFFD0 U754 ( .I(n770), .Z(n769) );
  BUFFD0 U755 ( .I(n771), .Z(n770) );
  BUFFD0 U756 ( .I(n772), .Z(n771) );
  BUFFD0 U757 ( .I(n773), .Z(n772) );
  BUFFD0 U758 ( .I(n774), .Z(n773) );
  BUFFD0 U759 ( .I(n775), .Z(n774) );
  BUFFD0 U760 ( .I(n776), .Z(n775) );
  BUFFD0 U761 ( .I(n777), .Z(n776) );
  BUFFD0 U762 ( .I(n778), .Z(n777) );
  BUFFD0 U763 ( .I(n779), .Z(n778) );
  BUFFD0 U764 ( .I(n780), .Z(n779) );
  BUFFD0 U765 ( .I(n781), .Z(n780) );
  BUFFD0 U766 ( .I(n782), .Z(n781) );
  BUFFD0 U767 ( .I(n783), .Z(n782) );
  BUFFD0 U768 ( .I(n784), .Z(n783) );
  BUFFD0 U769 ( .I(n785), .Z(n784) );
  BUFFD0 U770 ( .I(n786), .Z(n785) );
  BUFFD0 U771 ( .I(n787), .Z(n786) );
  BUFFD0 U772 ( .I(n788), .Z(n787) );
  BUFFD0 U773 ( .I(n789), .Z(n788) );
  BUFFD0 U774 ( .I(n790), .Z(n789) );
  BUFFD0 U775 ( .I(DataOr[18]), .Z(n790) );
  BUFFD0 U776 ( .I(n792), .Z(n791) );
  BUFFD0 U777 ( .I(n793), .Z(n792) );
  BUFFD0 U778 ( .I(n794), .Z(n793) );
  BUFFD0 U779 ( .I(n795), .Z(n794) );
  BUFFD0 U780 ( .I(n796), .Z(n795) );
  BUFFD0 U781 ( .I(n797), .Z(n796) );
  BUFFD0 U782 ( .I(n798), .Z(n797) );
  BUFFD0 U783 ( .I(n799), .Z(n798) );
  BUFFD0 U784 ( .I(n800), .Z(n799) );
  BUFFD0 U785 ( .I(n801), .Z(n800) );
  BUFFD0 U786 ( .I(n802), .Z(n801) );
  BUFFD0 U787 ( .I(n803), .Z(n802) );
  BUFFD0 U788 ( .I(n804), .Z(n803) );
  BUFFD0 U789 ( .I(n805), .Z(n804) );
  BUFFD0 U790 ( .I(n806), .Z(n805) );
  BUFFD0 U791 ( .I(n807), .Z(n806) );
  BUFFD0 U792 ( .I(n808), .Z(n807) );
  BUFFD0 U793 ( .I(n809), .Z(n808) );
  BUFFD0 U794 ( .I(n810), .Z(n809) );
  BUFFD0 U795 ( .I(n811), .Z(n810) );
  BUFFD0 U796 ( .I(n812), .Z(n811) );
  BUFFD0 U797 ( .I(n813), .Z(n812) );
  BUFFD0 U798 ( .I(n814), .Z(n813) );
  BUFFD0 U799 ( .I(n815), .Z(n814) );
  BUFFD0 U800 ( .I(n816), .Z(n815) );
  BUFFD0 U801 ( .I(n817), .Z(n816) );
  BUFFD0 U802 ( .I(n818), .Z(n817) );
  BUFFD0 U803 ( .I(n819), .Z(n818) );
  BUFFD0 U804 ( .I(n820), .Z(n819) );
  BUFFD0 U805 ( .I(n821), .Z(n820) );
  BUFFD0 U806 ( .I(n822), .Z(n821) );
  BUFFD0 U807 ( .I(n823), .Z(n822) );
  BUFFD0 U808 ( .I(n824), .Z(n823) );
  BUFFD0 U809 ( .I(n825), .Z(n824) );
  BUFFD0 U810 ( .I(n826), .Z(n825) );
  BUFFD0 U811 ( .I(n827), .Z(n826) );
  BUFFD0 U812 ( .I(n828), .Z(n827) );
  BUFFD0 U813 ( .I(n829), .Z(n828) );
  BUFFD0 U814 ( .I(n830), .Z(n829) );
  BUFFD0 U815 ( .I(n831), .Z(n830) );
  BUFFD0 U816 ( .I(n832), .Z(n831) );
  BUFFD0 U817 ( .I(n833), .Z(n832) );
  BUFFD0 U818 ( .I(n834), .Z(n833) );
  BUFFD0 U819 ( .I(n835), .Z(n834) );
  BUFFD0 U820 ( .I(n836), .Z(n835) );
  BUFFD0 U821 ( .I(n837), .Z(n836) );
  BUFFD0 U822 ( .I(n838), .Z(n837) );
  BUFFD0 U823 ( .I(n839), .Z(n838) );
  BUFFD0 U824 ( .I(n840), .Z(n839) );
  BUFFD0 U825 ( .I(n841), .Z(n840) );
  BUFFD0 U826 ( .I(n842), .Z(n841) );
  BUFFD0 U827 ( .I(n843), .Z(n842) );
  BUFFD0 U828 ( .I(n844), .Z(n843) );
  BUFFD0 U829 ( .I(DataOr[17]), .Z(n844) );
  BUFFD0 U830 ( .I(n846), .Z(n845) );
  BUFFD0 U831 ( .I(n847), .Z(n846) );
  BUFFD0 U832 ( .I(n848), .Z(n847) );
  BUFFD0 U833 ( .I(n849), .Z(n848) );
  BUFFD0 U834 ( .I(n850), .Z(n849) );
  BUFFD0 U835 ( .I(n851), .Z(n850) );
  BUFFD0 U836 ( .I(n852), .Z(n851) );
  BUFFD0 U837 ( .I(n853), .Z(n852) );
  BUFFD0 U838 ( .I(n854), .Z(n853) );
  BUFFD0 U839 ( .I(n855), .Z(n854) );
  BUFFD0 U840 ( .I(n856), .Z(n855) );
  BUFFD0 U841 ( .I(n857), .Z(n856) );
  BUFFD0 U842 ( .I(n858), .Z(n857) );
  BUFFD0 U843 ( .I(n859), .Z(n858) );
  BUFFD0 U844 ( .I(n860), .Z(n859) );
  BUFFD0 U845 ( .I(n861), .Z(n860) );
  BUFFD0 U846 ( .I(n862), .Z(n861) );
  BUFFD0 U847 ( .I(n863), .Z(n862) );
  BUFFD0 U848 ( .I(n864), .Z(n863) );
  BUFFD0 U849 ( .I(n865), .Z(n864) );
  BUFFD0 U850 ( .I(n866), .Z(n865) );
  BUFFD0 U851 ( .I(n867), .Z(n866) );
  BUFFD0 U852 ( .I(n868), .Z(n867) );
  BUFFD0 U853 ( .I(n869), .Z(n868) );
  BUFFD0 U854 ( .I(n870), .Z(n869) );
  BUFFD0 U855 ( .I(n871), .Z(n870) );
  BUFFD0 U856 ( .I(n872), .Z(n871) );
  BUFFD0 U857 ( .I(n873), .Z(n872) );
  BUFFD0 U858 ( .I(n874), .Z(n873) );
  BUFFD0 U859 ( .I(n875), .Z(n874) );
  BUFFD0 U860 ( .I(n876), .Z(n875) );
  BUFFD0 U861 ( .I(n877), .Z(n876) );
  BUFFD0 U862 ( .I(n878), .Z(n877) );
  BUFFD0 U863 ( .I(n879), .Z(n878) );
  BUFFD0 U864 ( .I(n880), .Z(n879) );
  BUFFD0 U865 ( .I(n881), .Z(n880) );
  BUFFD0 U866 ( .I(n882), .Z(n881) );
  BUFFD0 U867 ( .I(n883), .Z(n882) );
  BUFFD0 U868 ( .I(n884), .Z(n883) );
  BUFFD0 U869 ( .I(n885), .Z(n884) );
  BUFFD0 U870 ( .I(n886), .Z(n885) );
  BUFFD0 U871 ( .I(n887), .Z(n886) );
  BUFFD0 U872 ( .I(n888), .Z(n887) );
  BUFFD0 U873 ( .I(n889), .Z(n888) );
  BUFFD0 U874 ( .I(n890), .Z(n889) );
  BUFFD0 U875 ( .I(n891), .Z(n890) );
  BUFFD0 U876 ( .I(n892), .Z(n891) );
  BUFFD0 U877 ( .I(n893), .Z(n892) );
  BUFFD0 U878 ( .I(n894), .Z(n893) );
  BUFFD0 U879 ( .I(n895), .Z(n894) );
  BUFFD0 U880 ( .I(n896), .Z(n895) );
  BUFFD0 U881 ( .I(n897), .Z(n896) );
  BUFFD0 U882 ( .I(n898), .Z(n897) );
  BUFFD0 U883 ( .I(DataOr[16]), .Z(n898) );
  BUFFD0 U884 ( .I(n900), .Z(n899) );
  BUFFD0 U885 ( .I(n901), .Z(n900) );
  BUFFD0 U886 ( .I(n902), .Z(n901) );
  BUFFD0 U887 ( .I(n903), .Z(n902) );
  BUFFD0 U888 ( .I(n904), .Z(n903) );
  BUFFD0 U889 ( .I(n905), .Z(n904) );
  BUFFD0 U890 ( .I(n906), .Z(n905) );
  BUFFD0 U891 ( .I(n907), .Z(n906) );
  BUFFD0 U892 ( .I(n908), .Z(n907) );
  BUFFD0 U893 ( .I(n909), .Z(n908) );
  BUFFD0 U894 ( .I(n910), .Z(n909) );
  BUFFD0 U895 ( .I(n911), .Z(n910) );
  BUFFD0 U896 ( .I(n912), .Z(n911) );
  BUFFD0 U897 ( .I(n913), .Z(n912) );
  BUFFD0 U898 ( .I(n914), .Z(n913) );
  BUFFD0 U899 ( .I(n915), .Z(n914) );
  BUFFD0 U900 ( .I(n916), .Z(n915) );
  BUFFD0 U901 ( .I(n917), .Z(n916) );
  BUFFD0 U902 ( .I(n918), .Z(n917) );
  BUFFD0 U903 ( .I(n919), .Z(n918) );
  BUFFD0 U904 ( .I(n920), .Z(n919) );
  BUFFD0 U905 ( .I(n921), .Z(n920) );
  BUFFD0 U906 ( .I(n922), .Z(n921) );
  BUFFD0 U907 ( .I(n923), .Z(n922) );
  BUFFD0 U908 ( .I(n924), .Z(n923) );
  BUFFD0 U909 ( .I(n925), .Z(n924) );
  BUFFD0 U910 ( .I(n926), .Z(n925) );
  BUFFD0 U911 ( .I(n927), .Z(n926) );
  BUFFD0 U912 ( .I(n928), .Z(n927) );
  BUFFD0 U913 ( .I(n929), .Z(n928) );
  BUFFD0 U914 ( .I(n930), .Z(n929) );
  BUFFD0 U915 ( .I(n931), .Z(n930) );
  BUFFD0 U916 ( .I(n932), .Z(n931) );
  BUFFD0 U917 ( .I(n933), .Z(n932) );
  BUFFD0 U918 ( .I(n934), .Z(n933) );
  BUFFD0 U919 ( .I(n935), .Z(n934) );
  BUFFD0 U920 ( .I(n936), .Z(n935) );
  BUFFD0 U921 ( .I(n937), .Z(n936) );
  BUFFD0 U922 ( .I(n938), .Z(n937) );
  BUFFD0 U923 ( .I(n939), .Z(n938) );
  BUFFD0 U924 ( .I(n940), .Z(n939) );
  BUFFD0 U925 ( .I(n941), .Z(n940) );
  BUFFD0 U926 ( .I(n942), .Z(n941) );
  BUFFD0 U927 ( .I(n943), .Z(n942) );
  BUFFD0 U928 ( .I(n944), .Z(n943) );
  BUFFD0 U929 ( .I(n945), .Z(n944) );
  BUFFD0 U930 ( .I(n946), .Z(n945) );
  BUFFD0 U931 ( .I(n947), .Z(n946) );
  BUFFD0 U932 ( .I(n948), .Z(n947) );
  BUFFD0 U933 ( .I(n949), .Z(n948) );
  BUFFD0 U934 ( .I(n950), .Z(n949) );
  BUFFD0 U935 ( .I(n951), .Z(n950) );
  BUFFD0 U936 ( .I(n952), .Z(n951) );
  BUFFD0 U937 ( .I(DataOr[15]), .Z(n952) );
  BUFFD0 U938 ( .I(n954), .Z(n953) );
  BUFFD0 U939 ( .I(n955), .Z(n954) );
  BUFFD0 U940 ( .I(n956), .Z(n955) );
  BUFFD0 U941 ( .I(n957), .Z(n956) );
  BUFFD0 U942 ( .I(n958), .Z(n957) );
  BUFFD0 U943 ( .I(n959), .Z(n958) );
  BUFFD0 U944 ( .I(n960), .Z(n959) );
  BUFFD0 U945 ( .I(n961), .Z(n960) );
  BUFFD0 U946 ( .I(n962), .Z(n961) );
  BUFFD0 U947 ( .I(n963), .Z(n962) );
  BUFFD0 U948 ( .I(n964), .Z(n963) );
  BUFFD0 U949 ( .I(n965), .Z(n964) );
  BUFFD0 U950 ( .I(n966), .Z(n965) );
  BUFFD0 U951 ( .I(n967), .Z(n966) );
  BUFFD0 U952 ( .I(n968), .Z(n967) );
  BUFFD0 U953 ( .I(n969), .Z(n968) );
  BUFFD0 U954 ( .I(n970), .Z(n969) );
  BUFFD0 U955 ( .I(n971), .Z(n970) );
  BUFFD0 U956 ( .I(n972), .Z(n971) );
  BUFFD0 U957 ( .I(n973), .Z(n972) );
  BUFFD0 U958 ( .I(n974), .Z(n973) );
  BUFFD0 U959 ( .I(n975), .Z(n974) );
  BUFFD0 U960 ( .I(n976), .Z(n975) );
  BUFFD0 U961 ( .I(n977), .Z(n976) );
  BUFFD0 U962 ( .I(n978), .Z(n977) );
  BUFFD0 U963 ( .I(n979), .Z(n978) );
  BUFFD0 U964 ( .I(n980), .Z(n979) );
  BUFFD0 U965 ( .I(n981), .Z(n980) );
  BUFFD0 U966 ( .I(n982), .Z(n981) );
  BUFFD0 U967 ( .I(n983), .Z(n982) );
  BUFFD0 U968 ( .I(n984), .Z(n983) );
  BUFFD0 U969 ( .I(n985), .Z(n984) );
  BUFFD0 U970 ( .I(n986), .Z(n985) );
  BUFFD0 U971 ( .I(n987), .Z(n986) );
  BUFFD0 U972 ( .I(n988), .Z(n987) );
  BUFFD0 U973 ( .I(n989), .Z(n988) );
  BUFFD0 U974 ( .I(n990), .Z(n989) );
  BUFFD0 U975 ( .I(n991), .Z(n990) );
  BUFFD0 U976 ( .I(n992), .Z(n991) );
  BUFFD0 U977 ( .I(n993), .Z(n992) );
  BUFFD0 U978 ( .I(n994), .Z(n993) );
  BUFFD0 U979 ( .I(n995), .Z(n994) );
  BUFFD0 U980 ( .I(n996), .Z(n995) );
  BUFFD0 U981 ( .I(n997), .Z(n996) );
  BUFFD0 U982 ( .I(n998), .Z(n997) );
  BUFFD0 U983 ( .I(n999), .Z(n998) );
  BUFFD0 U984 ( .I(n1000), .Z(n999) );
  BUFFD0 U985 ( .I(n1001), .Z(n1000) );
  BUFFD0 U986 ( .I(n1002), .Z(n1001) );
  BUFFD0 U987 ( .I(n1003), .Z(n1002) );
  BUFFD0 U988 ( .I(n1004), .Z(n1003) );
  BUFFD0 U989 ( .I(n1005), .Z(n1004) );
  BUFFD0 U990 ( .I(n1006), .Z(n1005) );
  BUFFD0 U991 ( .I(DataOr[14]), .Z(n1006) );
  BUFFD0 U992 ( .I(n1008), .Z(n1007) );
  BUFFD0 U993 ( .I(n1009), .Z(n1008) );
  BUFFD0 U994 ( .I(n1010), .Z(n1009) );
  BUFFD0 U995 ( .I(n1011), .Z(n1010) );
  BUFFD0 U996 ( .I(n1012), .Z(n1011) );
  BUFFD0 U997 ( .I(n1013), .Z(n1012) );
  BUFFD0 U998 ( .I(n1014), .Z(n1013) );
  BUFFD0 U999 ( .I(n1015), .Z(n1014) );
  BUFFD0 U1000 ( .I(n1016), .Z(n1015) );
  BUFFD0 U1001 ( .I(n1017), .Z(n1016) );
  BUFFD0 U1002 ( .I(n1018), .Z(n1017) );
  BUFFD0 U1003 ( .I(n1019), .Z(n1018) );
  BUFFD0 U1004 ( .I(n1020), .Z(n1019) );
  BUFFD0 U1005 ( .I(n1021), .Z(n1020) );
  BUFFD0 U1006 ( .I(n1022), .Z(n1021) );
  BUFFD0 U1007 ( .I(n1023), .Z(n1022) );
  BUFFD0 U1008 ( .I(n1024), .Z(n1023) );
  BUFFD0 U1009 ( .I(n1025), .Z(n1024) );
  BUFFD0 U1010 ( .I(n1026), .Z(n1025) );
  BUFFD0 U1011 ( .I(n1027), .Z(n1026) );
  BUFFD0 U1012 ( .I(n1028), .Z(n1027) );
  BUFFD0 U1013 ( .I(n1029), .Z(n1028) );
  BUFFD0 U1014 ( .I(n1030), .Z(n1029) );
  BUFFD0 U1015 ( .I(n1031), .Z(n1030) );
  BUFFD0 U1016 ( .I(n1032), .Z(n1031) );
  BUFFD0 U1017 ( .I(n1033), .Z(n1032) );
  BUFFD0 U1018 ( .I(n1034), .Z(n1033) );
  BUFFD0 U1019 ( .I(n1035), .Z(n1034) );
  BUFFD0 U1020 ( .I(n1036), .Z(n1035) );
  BUFFD0 U1021 ( .I(n1037), .Z(n1036) );
  BUFFD0 U1022 ( .I(n1038), .Z(n1037) );
  BUFFD0 U1023 ( .I(n1039), .Z(n1038) );
  BUFFD0 U1024 ( .I(n1040), .Z(n1039) );
  BUFFD0 U1025 ( .I(n1041), .Z(n1040) );
  BUFFD0 U1026 ( .I(n1042), .Z(n1041) );
  BUFFD0 U1027 ( .I(n1043), .Z(n1042) );
  BUFFD0 U1028 ( .I(n1044), .Z(n1043) );
  BUFFD0 U1029 ( .I(n1045), .Z(n1044) );
  BUFFD0 U1030 ( .I(n1046), .Z(n1045) );
  BUFFD0 U1031 ( .I(n1047), .Z(n1046) );
  BUFFD0 U1032 ( .I(n1048), .Z(n1047) );
  BUFFD0 U1033 ( .I(n1049), .Z(n1048) );
  BUFFD0 U1034 ( .I(n1050), .Z(n1049) );
  BUFFD0 U1035 ( .I(n1051), .Z(n1050) );
  BUFFD0 U1036 ( .I(n1052), .Z(n1051) );
  BUFFD0 U1037 ( .I(n1053), .Z(n1052) );
  BUFFD0 U1038 ( .I(n1054), .Z(n1053) );
  BUFFD0 U1039 ( .I(n1055), .Z(n1054) );
  BUFFD0 U1040 ( .I(n1056), .Z(n1055) );
  BUFFD0 U1041 ( .I(n1057), .Z(n1056) );
  BUFFD0 U1042 ( .I(n1058), .Z(n1057) );
  BUFFD0 U1043 ( .I(n1059), .Z(n1058) );
  BUFFD0 U1044 ( .I(n1060), .Z(n1059) );
  BUFFD0 U1045 ( .I(DataOr[13]), .Z(n1060) );
  BUFFD0 U1046 ( .I(n1062), .Z(n1061) );
  BUFFD0 U1047 ( .I(n1063), .Z(n1062) );
  BUFFD0 U1048 ( .I(n1064), .Z(n1063) );
  BUFFD0 U1049 ( .I(n1065), .Z(n1064) );
  BUFFD0 U1050 ( .I(n1066), .Z(n1065) );
  BUFFD0 U1051 ( .I(n1067), .Z(n1066) );
  BUFFD0 U1052 ( .I(n1068), .Z(n1067) );
  BUFFD0 U1053 ( .I(n1069), .Z(n1068) );
  BUFFD0 U1054 ( .I(n1070), .Z(n1069) );
  BUFFD0 U1055 ( .I(n1071), .Z(n1070) );
  BUFFD0 U1056 ( .I(n1072), .Z(n1071) );
  BUFFD0 U1057 ( .I(n1073), .Z(n1072) );
  BUFFD0 U1058 ( .I(n1074), .Z(n1073) );
  BUFFD0 U1059 ( .I(n1075), .Z(n1074) );
  BUFFD0 U1060 ( .I(n1076), .Z(n1075) );
  BUFFD0 U1061 ( .I(n1077), .Z(n1076) );
  BUFFD0 U1062 ( .I(n1078), .Z(n1077) );
  BUFFD0 U1063 ( .I(n1079), .Z(n1078) );
  BUFFD0 U1064 ( .I(n1080), .Z(n1079) );
  BUFFD0 U1065 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1066 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1067 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1068 ( .I(n1084), .Z(n1083) );
  BUFFD0 U1069 ( .I(n1085), .Z(n1084) );
  BUFFD0 U1070 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1071 ( .I(n1087), .Z(n1086) );
  BUFFD0 U1072 ( .I(n1088), .Z(n1087) );
  BUFFD0 U1073 ( .I(n1089), .Z(n1088) );
  BUFFD0 U1074 ( .I(n1090), .Z(n1089) );
  BUFFD0 U1075 ( .I(n1091), .Z(n1090) );
  BUFFD0 U1076 ( .I(n1092), .Z(n1091) );
  BUFFD0 U1077 ( .I(n1093), .Z(n1092) );
  BUFFD0 U1078 ( .I(n1094), .Z(n1093) );
  BUFFD0 U1079 ( .I(n1095), .Z(n1094) );
  BUFFD0 U1080 ( .I(n1096), .Z(n1095) );
  BUFFD0 U1081 ( .I(n1097), .Z(n1096) );
  BUFFD0 U1082 ( .I(n1098), .Z(n1097) );
  BUFFD0 U1083 ( .I(n1099), .Z(n1098) );
  BUFFD0 U1084 ( .I(n1100), .Z(n1099) );
  BUFFD0 U1085 ( .I(n1101), .Z(n1100) );
  BUFFD0 U1086 ( .I(n1102), .Z(n1101) );
  BUFFD0 U1087 ( .I(n1103), .Z(n1102) );
  BUFFD0 U1088 ( .I(n1104), .Z(n1103) );
  BUFFD0 U1089 ( .I(n1105), .Z(n1104) );
  BUFFD0 U1090 ( .I(n1106), .Z(n1105) );
  BUFFD0 U1091 ( .I(n1107), .Z(n1106) );
  BUFFD0 U1092 ( .I(n1108), .Z(n1107) );
  BUFFD0 U1093 ( .I(n1109), .Z(n1108) );
  BUFFD0 U1094 ( .I(n1110), .Z(n1109) );
  BUFFD0 U1095 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1096 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1097 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1098 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1099 ( .I(DataOr[12]), .Z(n1114) );
  BUFFD0 U1100 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1101 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1102 ( .I(n1118), .Z(n1117) );
  BUFFD0 U1103 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1104 ( .I(n1120), .Z(n1119) );
  BUFFD0 U1105 ( .I(n1121), .Z(n1120) );
  BUFFD0 U1106 ( .I(n1122), .Z(n1121) );
  BUFFD0 U1107 ( .I(n1123), .Z(n1122) );
  BUFFD0 U1108 ( .I(n1124), .Z(n1123) );
  BUFFD0 U1109 ( .I(n1125), .Z(n1124) );
  BUFFD0 U1110 ( .I(n1126), .Z(n1125) );
  BUFFD0 U1111 ( .I(n1127), .Z(n1126) );
  BUFFD0 U1112 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1113 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1114 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1115 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1116 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1117 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1118 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1119 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1120 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1121 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1122 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1123 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1124 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1125 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1126 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1127 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1128 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1129 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1130 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1131 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1132 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1133 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1134 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1135 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1136 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1137 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1138 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1139 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1140 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1141 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1142 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1143 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1144 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1145 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1146 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1147 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1148 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1149 ( .I(n1165), .Z(n1164) );
  BUFFD0 U1150 ( .I(n1166), .Z(n1165) );
  BUFFD0 U1151 ( .I(n1167), .Z(n1166) );
  BUFFD0 U1152 ( .I(n1168), .Z(n1167) );
  BUFFD0 U1153 ( .I(DataOr[11]), .Z(n1168) );
  BUFFD0 U1154 ( .I(n1170), .Z(n1169) );
  BUFFD0 U1155 ( .I(n1171), .Z(n1170) );
  BUFFD0 U1156 ( .I(n1172), .Z(n1171) );
  BUFFD0 U1157 ( .I(n1173), .Z(n1172) );
  BUFFD0 U1158 ( .I(n1174), .Z(n1173) );
  BUFFD0 U1159 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1160 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1161 ( .I(n1177), .Z(n1176) );
  BUFFD0 U1162 ( .I(n1178), .Z(n1177) );
  BUFFD0 U1163 ( .I(n1179), .Z(n1178) );
  BUFFD0 U1164 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1165 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1166 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1167 ( .I(n1183), .Z(n1182) );
  BUFFD0 U1168 ( .I(n1184), .Z(n1183) );
  BUFFD0 U1169 ( .I(n1185), .Z(n1184) );
  BUFFD0 U1170 ( .I(n1186), .Z(n1185) );
  BUFFD0 U1171 ( .I(n1187), .Z(n1186) );
  BUFFD0 U1172 ( .I(n1188), .Z(n1187) );
  BUFFD0 U1173 ( .I(n1189), .Z(n1188) );
  BUFFD0 U1174 ( .I(n1190), .Z(n1189) );
  BUFFD0 U1175 ( .I(n1191), .Z(n1190) );
  BUFFD0 U1176 ( .I(n1192), .Z(n1191) );
  BUFFD0 U1177 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1178 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1179 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1180 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1181 ( .I(n1197), .Z(n1196) );
  BUFFD0 U1182 ( .I(n1198), .Z(n1197) );
  BUFFD0 U1183 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1184 ( .I(n1200), .Z(n1199) );
  BUFFD0 U1185 ( .I(n1201), .Z(n1200) );
  BUFFD0 U1186 ( .I(n1202), .Z(n1201) );
  BUFFD0 U1187 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1188 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1189 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1190 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1191 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1192 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1193 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1194 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1195 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1196 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1197 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1198 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1199 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1200 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1201 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1202 ( .I(n1218), .Z(n1217) );
  BUFFD0 U1203 ( .I(n1219), .Z(n1218) );
  BUFFD0 U1204 ( .I(n1220), .Z(n1219) );
  BUFFD0 U1205 ( .I(n1221), .Z(n1220) );
  BUFFD0 U1206 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1207 ( .I(DataOr[10]), .Z(n1222) );
  BUFFD0 U1208 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1209 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1210 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1211 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1212 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1213 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1214 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1215 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1216 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1217 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1218 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1219 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1220 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1221 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1222 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1223 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1224 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1225 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1226 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1227 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1228 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1229 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1230 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1231 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1232 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1233 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1234 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1235 ( .I(n1251), .Z(n1250) );
  BUFFD0 U1236 ( .I(n1252), .Z(n1251) );
  BUFFD0 U1237 ( .I(n1253), .Z(n1252) );
  BUFFD0 U1238 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1239 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1240 ( .I(n1256), .Z(n1255) );
  BUFFD0 U1241 ( .I(n1257), .Z(n1256) );
  BUFFD0 U1242 ( .I(n1258), .Z(n1257) );
  BUFFD0 U1243 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1244 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1245 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1246 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1247 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1248 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1249 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1250 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1251 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1252 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1253 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1254 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1255 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1256 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1257 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1258 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1259 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1260 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1261 ( .I(DataOr[9]), .Z(n1276) );
  BUFFD0 U1262 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1263 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1264 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1265 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1266 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1267 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1268 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1269 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1270 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1271 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1272 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1273 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1274 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1275 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1276 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1277 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1278 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1279 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1280 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1281 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1282 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1283 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1284 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1285 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1286 ( .I(n1302), .Z(n1301) );
  BUFFD0 U1287 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1288 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1289 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1290 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1291 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1292 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1293 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1294 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1295 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1296 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1297 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1298 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1299 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1300 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1301 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1302 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1303 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1304 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1305 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1306 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1307 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1308 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1309 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1310 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1311 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1312 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1313 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1314 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1315 ( .I(DataOr[8]), .Z(n1330) );
  BUFFD0 U1316 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1317 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1318 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1319 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1320 ( .I(n1336), .Z(n1335) );
  BUFFD0 U1321 ( .I(n1337), .Z(n1336) );
  BUFFD0 U1322 ( .I(n1338), .Z(n1337) );
  BUFFD0 U1323 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1324 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1325 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1326 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1327 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1328 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1329 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1330 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1331 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1332 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1333 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1334 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1335 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1336 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1337 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1338 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1339 ( .I(n1355), .Z(n1354) );
  BUFFD0 U1340 ( .I(n1356), .Z(n1355) );
  BUFFD0 U1341 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1342 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1343 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1344 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1345 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1346 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1347 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1348 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1349 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1350 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1351 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1352 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1353 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1354 ( .I(n1370), .Z(n1369) );
  BUFFD0 U1355 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1356 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1357 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1358 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1359 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1360 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1361 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1362 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1363 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1364 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1365 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1366 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1367 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1368 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1369 ( .I(DataOr[7]), .Z(n1384) );
  BUFFD0 U1370 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1371 ( .I(n1387), .Z(n1386) );
  BUFFD0 U1372 ( .I(n1388), .Z(n1387) );
  BUFFD0 U1373 ( .I(n1389), .Z(n1388) );
  BUFFD0 U1374 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1375 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1376 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1377 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1378 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1379 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1380 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1381 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1382 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1383 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1384 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1385 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1386 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1387 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1388 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1389 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1390 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1391 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1392 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1393 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1394 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1395 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1396 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1397 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1398 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1399 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1400 ( .I(n1416), .Z(n1415) );
  BUFFD0 U1401 ( .I(n1417), .Z(n1416) );
  BUFFD0 U1402 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1403 ( .I(n1419), .Z(n1418) );
  BUFFD0 U1404 ( .I(n1420), .Z(n1419) );
  BUFFD0 U1405 ( .I(n1421), .Z(n1420) );
  BUFFD0 U1406 ( .I(n1422), .Z(n1421) );
  BUFFD0 U1407 ( .I(n1423), .Z(n1422) );
  BUFFD0 U1408 ( .I(n1424), .Z(n1423) );
  BUFFD0 U1409 ( .I(n1425), .Z(n1424) );
  BUFFD0 U1410 ( .I(n1426), .Z(n1425) );
  BUFFD0 U1411 ( .I(n1427), .Z(n1426) );
  BUFFD0 U1412 ( .I(n1428), .Z(n1427) );
  BUFFD0 U1413 ( .I(n1429), .Z(n1428) );
  BUFFD0 U1414 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1415 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1416 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1417 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1418 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1419 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1420 ( .I(n1436), .Z(n1435) );
  BUFFD0 U1421 ( .I(n1437), .Z(n1436) );
  BUFFD0 U1422 ( .I(n1438), .Z(n1437) );
  BUFFD0 U1423 ( .I(DataOr[6]), .Z(n1438) );
  BUFFD0 U1424 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1425 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1426 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1427 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1428 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1429 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1430 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1431 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1432 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1433 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1434 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1435 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1436 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1437 ( .I(n1453), .Z(n1452) );
  BUFFD0 U1438 ( .I(n1454), .Z(n1453) );
  BUFFD0 U1439 ( .I(n1455), .Z(n1454) );
  BUFFD0 U1440 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1441 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1442 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1443 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1444 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1445 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1446 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1447 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1448 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1449 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1450 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1451 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1452 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1453 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1454 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1455 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1456 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1457 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1458 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1459 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1460 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1461 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1462 ( .I(n1478), .Z(n1477) );
  BUFFD0 U1463 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1464 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1465 ( .I(n1481), .Z(n1480) );
  BUFFD0 U1466 ( .I(n1482), .Z(n1481) );
  BUFFD0 U1467 ( .I(n1483), .Z(n1482) );
  BUFFD0 U1468 ( .I(n1484), .Z(n1483) );
  BUFFD0 U1469 ( .I(n1485), .Z(n1484) );
  BUFFD0 U1470 ( .I(n1486), .Z(n1485) );
  BUFFD0 U1471 ( .I(n1487), .Z(n1486) );
  BUFFD0 U1472 ( .I(n1488), .Z(n1487) );
  BUFFD0 U1473 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1474 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1475 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1476 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1477 ( .I(DataOr[5]), .Z(n1492) );
  BUFFD0 U1478 ( .I(n1494), .Z(n1493) );
  BUFFD0 U1479 ( .I(n1495), .Z(n1494) );
  BUFFD0 U1480 ( .I(n1496), .Z(n1495) );
  BUFFD0 U1481 ( .I(n1497), .Z(n1496) );
  BUFFD0 U1482 ( .I(n1498), .Z(n1497) );
  BUFFD0 U1483 ( .I(n1499), .Z(n1498) );
  BUFFD0 U1484 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1485 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1486 ( .I(n1502), .Z(n1501) );
  BUFFD0 U1487 ( .I(n1503), .Z(n1502) );
  BUFFD0 U1488 ( .I(n1504), .Z(n1503) );
  BUFFD0 U1489 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1490 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1491 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1492 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1493 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1494 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1495 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1496 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1497 ( .I(n1513), .Z(n1512) );
  BUFFD0 U1498 ( .I(n1514), .Z(n1513) );
  BUFFD0 U1499 ( .I(n1515), .Z(n1514) );
  BUFFD0 U1500 ( .I(n1516), .Z(n1515) );
  BUFFD0 U1501 ( .I(n1517), .Z(n1516) );
  BUFFD0 U1502 ( .I(n1518), .Z(n1517) );
  BUFFD0 U1503 ( .I(n1519), .Z(n1518) );
  BUFFD0 U1504 ( .I(n1520), .Z(n1519) );
  BUFFD0 U1505 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1506 ( .I(n1522), .Z(n1521) );
  BUFFD0 U1507 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1508 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1509 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1510 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1511 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1512 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1513 ( .I(n1529), .Z(n1528) );
  BUFFD0 U1514 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1515 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1516 ( .I(n1532), .Z(n1531) );
  BUFFD0 U1517 ( .I(n1533), .Z(n1532) );
  BUFFD0 U1518 ( .I(n1534), .Z(n1533) );
  BUFFD0 U1519 ( .I(n1535), .Z(n1534) );
  BUFFD0 U1520 ( .I(n1536), .Z(n1535) );
  BUFFD0 U1521 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1522 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1523 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1524 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1525 ( .I(n1541), .Z(n1540) );
  BUFFD0 U1526 ( .I(n1542), .Z(n1541) );
  BUFFD0 U1527 ( .I(n1543), .Z(n1542) );
  BUFFD0 U1528 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1529 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1530 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1531 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1532 ( .I(DataOr[4]), .Z(n1547) );
  BUFFD0 U1533 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1534 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1535 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1536 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1537 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1538 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1539 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1540 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1541 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1542 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1543 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1544 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1545 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1546 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1547 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1548 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1549 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1550 ( .I(n1566), .Z(n1565) );
  BUFFD0 U1551 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1552 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1553 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1554 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1555 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1556 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1557 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1558 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1559 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1560 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1561 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1562 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1563 ( .I(n1579), .Z(n1578) );
  BUFFD0 U1564 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1565 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1566 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1567 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1568 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1569 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1570 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1571 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1572 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1573 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1574 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1575 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1576 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1577 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1578 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1579 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1580 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1581 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1582 ( .I(n1598), .Z(n1597) );
  BUFFD0 U1583 ( .I(n1599), .Z(n1598) );
  BUFFD0 U1584 ( .I(n1600), .Z(n1599) );
  BUFFD0 U1585 ( .I(n1601), .Z(n1600) );
  BUFFD0 U1586 ( .I(n1602), .Z(n1601) );
  BUFFD0 U1587 ( .I(DataOr[3]), .Z(n1602) );
  BUFFD0 U1588 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1589 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1590 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1591 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1592 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1593 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1594 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1595 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1596 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1597 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1598 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1599 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1600 ( .I(n1616), .Z(n1615) );
  BUFFD0 U1601 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1602 ( .I(n1618), .Z(n1617) );
  BUFFD0 U1603 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1604 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1605 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1606 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1607 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1608 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1609 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1610 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1611 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1612 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1613 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1614 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1615 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1616 ( .I(n1632), .Z(n1631) );
  BUFFD0 U1617 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1618 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1619 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1620 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1621 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1622 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1623 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1624 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1625 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1626 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1627 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1628 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1629 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1630 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1631 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1632 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1633 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1634 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1635 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1636 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1637 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1638 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1639 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1640 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1641 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1642 ( .I(DataOr[2]), .Z(n1657) );
  BUFFD0 U1643 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1644 ( .I(n1660), .Z(n1659) );
  BUFFD0 U1645 ( .I(n1661), .Z(n1660) );
  BUFFD0 U1646 ( .I(n1662), .Z(n1661) );
  BUFFD0 U1647 ( .I(n1663), .Z(n1662) );
  BUFFD0 U1648 ( .I(n1664), .Z(n1663) );
  BUFFD0 U1649 ( .I(n1665), .Z(n1664) );
  BUFFD0 U1650 ( .I(n1666), .Z(n1665) );
  BUFFD0 U1651 ( .I(n1667), .Z(n1666) );
  BUFFD0 U1652 ( .I(n1668), .Z(n1667) );
  BUFFD0 U1653 ( .I(n1669), .Z(n1668) );
  BUFFD0 U1654 ( .I(n1670), .Z(n1669) );
  BUFFD0 U1655 ( .I(n1671), .Z(n1670) );
  BUFFD0 U1656 ( .I(n1672), .Z(n1671) );
  BUFFD0 U1657 ( .I(n1673), .Z(n1672) );
  BUFFD0 U1658 ( .I(n1674), .Z(n1673) );
  BUFFD0 U1659 ( .I(n1675), .Z(n1674) );
  BUFFD0 U1660 ( .I(n1676), .Z(n1675) );
  BUFFD0 U1661 ( .I(n1677), .Z(n1676) );
  BUFFD0 U1662 ( .I(n1678), .Z(n1677) );
  BUFFD0 U1663 ( .I(n1679), .Z(n1678) );
  BUFFD0 U1664 ( .I(n1680), .Z(n1679) );
  BUFFD0 U1665 ( .I(n1681), .Z(n1680) );
  BUFFD0 U1666 ( .I(n1682), .Z(n1681) );
  BUFFD0 U1667 ( .I(n1683), .Z(n1682) );
  BUFFD0 U1668 ( .I(n1684), .Z(n1683) );
  BUFFD0 U1669 ( .I(n1685), .Z(n1684) );
  BUFFD0 U1670 ( .I(n1686), .Z(n1685) );
  BUFFD0 U1671 ( .I(n1687), .Z(n1686) );
  BUFFD0 U1672 ( .I(n1688), .Z(n1687) );
  BUFFD0 U1673 ( .I(n1689), .Z(n1688) );
  BUFFD0 U1674 ( .I(n1690), .Z(n1689) );
  BUFFD0 U1675 ( .I(n1691), .Z(n1690) );
  BUFFD0 U1676 ( .I(n1692), .Z(n1691) );
  BUFFD0 U1677 ( .I(n1693), .Z(n1692) );
  BUFFD0 U1678 ( .I(n1694), .Z(n1693) );
  BUFFD0 U1679 ( .I(n1695), .Z(n1694) );
  BUFFD0 U1680 ( .I(n1696), .Z(n1695) );
  BUFFD0 U1681 ( .I(n1697), .Z(n1696) );
  BUFFD0 U1682 ( .I(n1698), .Z(n1697) );
  BUFFD0 U1683 ( .I(n1699), .Z(n1698) );
  BUFFD0 U1684 ( .I(n1700), .Z(n1699) );
  BUFFD0 U1685 ( .I(n1701), .Z(n1700) );
  BUFFD0 U1686 ( .I(n1702), .Z(n1701) );
  BUFFD0 U1687 ( .I(n1703), .Z(n1702) );
  BUFFD0 U1688 ( .I(n1704), .Z(n1703) );
  BUFFD0 U1689 ( .I(n1705), .Z(n1704) );
  BUFFD0 U1690 ( .I(n1706), .Z(n1705) );
  BUFFD0 U1691 ( .I(n1707), .Z(n1706) );
  BUFFD0 U1692 ( .I(n1708), .Z(n1707) );
  BUFFD0 U1693 ( .I(n1709), .Z(n1708) );
  BUFFD0 U1694 ( .I(n1710), .Z(n1709) );
  BUFFD0 U1695 ( .I(n1711), .Z(n1710) );
  BUFFD0 U1696 ( .I(n1712), .Z(n1711) );
  BUFFD0 U1697 ( .I(DataOr[1]), .Z(n1712) );
  BUFFD0 U1698 ( .I(n1714), .Z(n1713) );
  BUFFD0 U1699 ( .I(n1715), .Z(n1714) );
  BUFFD0 U1700 ( .I(n1716), .Z(n1715) );
  BUFFD0 U1701 ( .I(n1717), .Z(n1716) );
  BUFFD0 U1702 ( .I(n1718), .Z(n1717) );
  BUFFD0 U1703 ( .I(n1719), .Z(n1718) );
  BUFFD0 U1704 ( .I(n1720), .Z(n1719) );
  BUFFD0 U1705 ( .I(n1721), .Z(n1720) );
  BUFFD0 U1706 ( .I(n1722), .Z(n1721) );
  BUFFD0 U1707 ( .I(n1723), .Z(n1722) );
  BUFFD0 U1708 ( .I(n1724), .Z(n1723) );
  BUFFD0 U1709 ( .I(n1725), .Z(n1724) );
  BUFFD0 U1710 ( .I(n1726), .Z(n1725) );
  BUFFD0 U1711 ( .I(n1727), .Z(n1726) );
  BUFFD0 U1712 ( .I(n1728), .Z(n1727) );
  BUFFD0 U1713 ( .I(n1729), .Z(n1728) );
  BUFFD0 U1714 ( .I(n1730), .Z(n1729) );
  BUFFD0 U1715 ( .I(n1731), .Z(n1730) );
  BUFFD0 U1716 ( .I(n1732), .Z(n1731) );
  BUFFD0 U1717 ( .I(n1733), .Z(n1732) );
  BUFFD0 U1718 ( .I(n1734), .Z(n1733) );
  BUFFD0 U1719 ( .I(n1735), .Z(n1734) );
  BUFFD0 U1720 ( .I(n1736), .Z(n1735) );
  BUFFD0 U1721 ( .I(n1737), .Z(n1736) );
  BUFFD0 U1722 ( .I(n1738), .Z(n1737) );
  BUFFD0 U1723 ( .I(n1739), .Z(n1738) );
  BUFFD0 U1724 ( .I(n1740), .Z(n1739) );
  BUFFD0 U1725 ( .I(n1741), .Z(n1740) );
  BUFFD0 U1726 ( .I(n1742), .Z(n1741) );
  BUFFD0 U1727 ( .I(n1743), .Z(n1742) );
  BUFFD0 U1728 ( .I(n1744), .Z(n1743) );
  BUFFD0 U1729 ( .I(n1745), .Z(n1744) );
  BUFFD0 U1730 ( .I(n1746), .Z(n1745) );
  BUFFD0 U1731 ( .I(n1747), .Z(n1746) );
  BUFFD0 U1732 ( .I(n1748), .Z(n1747) );
  BUFFD0 U1733 ( .I(n1749), .Z(n1748) );
  BUFFD0 U1734 ( .I(n1750), .Z(n1749) );
  BUFFD0 U1735 ( .I(n1751), .Z(n1750) );
  BUFFD0 U1736 ( .I(n1752), .Z(n1751) );
  BUFFD0 U1737 ( .I(n1753), .Z(n1752) );
  BUFFD0 U1738 ( .I(n1754), .Z(n1753) );
  BUFFD0 U1739 ( .I(n1755), .Z(n1754) );
  BUFFD0 U1740 ( .I(n1756), .Z(n1755) );
  BUFFD0 U1741 ( .I(n1757), .Z(n1756) );
  BUFFD0 U1742 ( .I(n1758), .Z(n1757) );
  BUFFD0 U1743 ( .I(n1759), .Z(n1758) );
  BUFFD0 U1744 ( .I(n1760), .Z(n1759) );
  BUFFD0 U1745 ( .I(n1761), .Z(n1760) );
  BUFFD0 U1746 ( .I(n1762), .Z(n1761) );
  BUFFD0 U1747 ( .I(n1763), .Z(n1762) );
  BUFFD0 U1748 ( .I(n1764), .Z(n1763) );
  BUFFD0 U1749 ( .I(n1765), .Z(n1764) );
  BUFFD0 U1750 ( .I(n1766), .Z(n1765) );
  BUFFD0 U1751 ( .I(n1767), .Z(n1766) );
  BUFFD0 U1752 ( .I(DataOr[0]), .Z(n1767) );
  BUFFD0 U1753 ( .I(n1772), .Z(n1768) );
  BUFFD0 U1754 ( .I(n4180), .Z(n1769) );
  BUFFD0 U1755 ( .I(n1769), .Z(n1770) );
  BUFFD0 U1756 ( .I(n1770), .Z(n1771) );
  BUFFD0 U1757 ( .I(n1773), .Z(n1772) );
  BUFFD0 U1758 ( .I(n1774), .Z(n1773) );
  BUFFD0 U1759 ( .I(n1775), .Z(n1774) );
  BUFFD0 U1760 ( .I(n1776), .Z(n1775) );
  BUFFD0 U1761 ( .I(n1777), .Z(n1776) );
  BUFFD0 U1762 ( .I(n1778), .Z(n1777) );
  BUFFD0 U1763 ( .I(n1779), .Z(n1778) );
  BUFFD0 U1764 ( .I(n1780), .Z(n1779) );
  BUFFD0 U1765 ( .I(n1781), .Z(n1780) );
  BUFFD0 U1766 ( .I(n1782), .Z(n1781) );
  BUFFD0 U1767 ( .I(n1783), .Z(n1782) );
  BUFFD0 U1768 ( .I(n1784), .Z(n1783) );
  BUFFD0 U1769 ( .I(n1785), .Z(n1784) );
  BUFFD0 U1770 ( .I(n1786), .Z(n1785) );
  BUFFD0 U1771 ( .I(n1787), .Z(n1786) );
  BUFFD0 U1772 ( .I(n1788), .Z(n1787) );
  BUFFD0 U1773 ( .I(n1789), .Z(n1788) );
  BUFFD0 U1774 ( .I(n1790), .Z(n1789) );
  BUFFD0 U1775 ( .I(n1791), .Z(n1790) );
  BUFFD0 U1776 ( .I(n1792), .Z(n1791) );
  BUFFD0 U1777 ( .I(n1793), .Z(n1792) );
  BUFFD0 U1778 ( .I(n1794), .Z(n1793) );
  BUFFD0 U1779 ( .I(n1795), .Z(n1794) );
  BUFFD0 U1780 ( .I(n1796), .Z(n1795) );
  BUFFD0 U1781 ( .I(n1797), .Z(n1796) );
  BUFFD0 U1782 ( .I(n1798), .Z(n1797) );
  BUFFD0 U1783 ( .I(n1799), .Z(n1798) );
  BUFFD0 U1784 ( .I(n1800), .Z(n1799) );
  BUFFD0 U1785 ( .I(n1801), .Z(n1800) );
  BUFFD0 U1786 ( .I(n1802), .Z(n1801) );
  BUFFD0 U1787 ( .I(n1803), .Z(n1802) );
  BUFFD0 U1788 ( .I(n1804), .Z(n1803) );
  BUFFD0 U1789 ( .I(n1805), .Z(n1804) );
  BUFFD0 U1790 ( .I(n1806), .Z(n1805) );
  BUFFD0 U1791 ( .I(n1807), .Z(n1806) );
  BUFFD0 U1792 ( .I(n1808), .Z(n1807) );
  BUFFD0 U1793 ( .I(n1809), .Z(n1808) );
  BUFFD0 U1794 ( .I(n1810), .Z(n1809) );
  BUFFD0 U1795 ( .I(n1811), .Z(n1810) );
  BUFFD0 U1796 ( .I(n1812), .Z(n1811) );
  BUFFD0 U1797 ( .I(n1813), .Z(n1812) );
  BUFFD0 U1798 ( .I(n1814), .Z(n1813) );
  BUFFD0 U1799 ( .I(n1815), .Z(n1814) );
  BUFFD0 U1800 ( .I(n1816), .Z(n1815) );
  BUFFD0 U1801 ( .I(n1817), .Z(n1816) );
  BUFFD0 U1802 ( .I(n1818), .Z(n1817) );
  BUFFD0 U1803 ( .I(n1819), .Z(n1818) );
  BUFFD0 U1804 ( .I(n1820), .Z(n1819) );
  BUFFD0 U1805 ( .I(n1821), .Z(n1820) );
  BUFFD0 U1806 ( .I(n1822), .Z(n1821) );
  BUFFD0 U1807 ( .I(n1823), .Z(n1822) );
  BUFFD0 U1808 ( .I(n1824), .Z(n1823) );
  BUFFD0 U1809 ( .I(n1825), .Z(n1824) );
  BUFFD0 U1810 ( .I(n1826), .Z(n1825) );
  BUFFD0 U1811 ( .I(n1828), .Z(n1826) );
  BUFFD0 U1812 ( .I(n1830), .Z(n1827) );
  BUFFD0 U1813 ( .I(n1829), .Z(n1828) );
  BUFFD0 U1814 ( .I(n1771), .Z(n1829) );
  BUFFD0 U1815 ( .I(Dreadyr), .Z(n1830) );
  OR2D0 U1816 ( .A1(n4325), .A2(n1827), .Z(n4180) );
  BUFFD0 U1817 ( .I(n1832), .Z(n1831) );
  BUFFD0 U1818 ( .I(n1833), .Z(n1832) );
  BUFFD0 U1819 ( .I(n1834), .Z(n1833) );
  BUFFD0 U1820 ( .I(n1835), .Z(n1834) );
  BUFFD0 U1821 ( .I(n1836), .Z(n1835) );
  BUFFD0 U1822 ( .I(n1837), .Z(n1836) );
  BUFFD0 U1823 ( .I(n1838), .Z(n1837) );
  BUFFD0 U1824 ( .I(n1839), .Z(n1838) );
  BUFFD0 U1825 ( .I(n1840), .Z(n1839) );
  BUFFD0 U1826 ( .I(n1841), .Z(n1840) );
  BUFFD0 U1827 ( .I(n1842), .Z(n1841) );
  BUFFD0 U1828 ( .I(n1843), .Z(n1842) );
  BUFFD0 U1829 ( .I(n1844), .Z(n1843) );
  BUFFD0 U1830 ( .I(n1845), .Z(n1844) );
  BUFFD0 U1831 ( .I(n1846), .Z(n1845) );
  BUFFD0 U1832 ( .I(n1847), .Z(n1846) );
  BUFFD0 U1833 ( .I(n1848), .Z(n1847) );
  BUFFD0 U1834 ( .I(n1849), .Z(n1848) );
  BUFFD0 U1835 ( .I(n1850), .Z(n1849) );
  BUFFD0 U1836 ( .I(n1851), .Z(n1850) );
  BUFFD0 U1837 ( .I(n1852), .Z(n1851) );
  BUFFD0 U1838 ( .I(n1853), .Z(n1852) );
  BUFFD0 U1839 ( .I(n1854), .Z(n1853) );
  BUFFD0 U1840 ( .I(n1855), .Z(n1854) );
  BUFFD0 U1841 ( .I(n1856), .Z(n1855) );
  BUFFD0 U1842 ( .I(n1857), .Z(n1856) );
  BUFFD0 U1843 ( .I(n1858), .Z(n1857) );
  BUFFD0 U1844 ( .I(n1859), .Z(n1858) );
  BUFFD0 U1845 ( .I(n1860), .Z(n1859) );
  BUFFD0 U1846 ( .I(n1861), .Z(n1860) );
  BUFFD0 U1847 ( .I(n1862), .Z(n1861) );
  BUFFD0 U1848 ( .I(n1863), .Z(n1862) );
  BUFFD0 U1849 ( .I(n1864), .Z(n1863) );
  BUFFD0 U1850 ( .I(n1865), .Z(n1864) );
  BUFFD0 U1851 ( .I(n1866), .Z(n1865) );
  BUFFD0 U1852 ( .I(n1867), .Z(n1866) );
  BUFFD0 U1853 ( .I(n1868), .Z(n1867) );
  BUFFD0 U1854 ( .I(n1869), .Z(n1868) );
  BUFFD0 U1855 ( .I(n1870), .Z(n1869) );
  BUFFD0 U1856 ( .I(n1871), .Z(n1870) );
  BUFFD0 U1857 ( .I(n1872), .Z(n1871) );
  BUFFD0 U1858 ( .I(n1873), .Z(n1872) );
  BUFFD0 U1859 ( .I(n1874), .Z(n1873) );
  BUFFD0 U1860 ( .I(n1875), .Z(n1874) );
  BUFFD0 U1861 ( .I(n1876), .Z(n1875) );
  BUFFD0 U1862 ( .I(n1877), .Z(n1876) );
  BUFFD0 U1863 ( .I(n1878), .Z(n1877) );
  BUFFD0 U1864 ( .I(n1879), .Z(n1878) );
  BUFFD0 U1865 ( .I(n1880), .Z(n1879) );
  BUFFD0 U1866 ( .I(n1881), .Z(n1880) );
  BUFFD0 U1867 ( .I(n1882), .Z(n1881) );
  BUFFD0 U1868 ( .I(n1883), .Z(n1882) );
  BUFFD0 U1869 ( .I(n1884), .Z(n1883) );
  BUFFD0 U1870 ( .I(n1885), .Z(n1884) );
  BUFFD0 U1871 ( .I(n1886), .Z(n1885) );
  BUFFD0 U1872 ( .I(n1887), .Z(n1886) );
  BUFFD0 U1873 ( .I(n1888), .Z(n1887) );
  BUFFD0 U1874 ( .I(n1889), .Z(n1888) );
  BUFFD0 U1875 ( .I(n1890), .Z(n1889) );
  BUFFD0 U1876 ( .I(n1891), .Z(n1890) );
  BUFFD0 U1877 ( .I(n1892), .Z(n1891) );
  BUFFD0 U1878 ( .I(n1893), .Z(n1892) );
  BUFFD0 U1879 ( .I(n1894), .Z(n1893) );
  BUFFD0 U1880 ( .I(n1895), .Z(n1894) );
  BUFFD0 U1881 ( .I(n1896), .Z(n1895) );
  BUFFD0 U1882 ( .I(n1897), .Z(n1896) );
  BUFFD0 U1883 ( .I(n1898), .Z(n1897) );
  BUFFD0 U1884 ( .I(n1899), .Z(n1898) );
  BUFFD0 U1885 ( .I(n1900), .Z(n1899) );
  BUFFD0 U1886 ( .I(N53), .Z(n1900) );
  BUFFD0 U1887 ( .I(n1902), .Z(n1901) );
  BUFFD0 U1888 ( .I(n1903), .Z(n1902) );
  BUFFD0 U1889 ( .I(n1904), .Z(n1903) );
  BUFFD0 U1890 ( .I(n1905), .Z(n1904) );
  BUFFD0 U1891 ( .I(n1906), .Z(n1905) );
  BUFFD0 U1892 ( .I(n1907), .Z(n1906) );
  BUFFD0 U1893 ( .I(n1908), .Z(n1907) );
  BUFFD0 U1894 ( .I(n1909), .Z(n1908) );
  BUFFD0 U1895 ( .I(n1910), .Z(n1909) );
  BUFFD0 U1896 ( .I(n1911), .Z(n1910) );
  BUFFD0 U1897 ( .I(n1912), .Z(n1911) );
  BUFFD0 U1898 ( .I(n1913), .Z(n1912) );
  BUFFD0 U1899 ( .I(n1914), .Z(n1913) );
  BUFFD0 U1900 ( .I(n1915), .Z(n1914) );
  BUFFD0 U1901 ( .I(n1916), .Z(n1915) );
  BUFFD0 U1902 ( .I(n1917), .Z(n1916) );
  BUFFD0 U1903 ( .I(n1918), .Z(n1917) );
  BUFFD0 U1904 ( .I(n1919), .Z(n1918) );
  BUFFD0 U1905 ( .I(n1920), .Z(n1919) );
  BUFFD0 U1906 ( .I(n1921), .Z(n1920) );
  BUFFD0 U1907 ( .I(n1922), .Z(n1921) );
  BUFFD0 U1908 ( .I(n1923), .Z(n1922) );
  BUFFD0 U1909 ( .I(n1924), .Z(n1923) );
  BUFFD0 U1910 ( .I(n1925), .Z(n1924) );
  BUFFD0 U1911 ( .I(n1926), .Z(n1925) );
  BUFFD0 U1912 ( .I(n1927), .Z(n1926) );
  BUFFD0 U1913 ( .I(n1928), .Z(n1927) );
  BUFFD0 U1914 ( .I(n1929), .Z(n1928) );
  BUFFD0 U1915 ( .I(n1930), .Z(n1929) );
  BUFFD0 U1916 ( .I(n1931), .Z(n1930) );
  BUFFD0 U1917 ( .I(n1932), .Z(n1931) );
  BUFFD0 U1918 ( .I(n1933), .Z(n1932) );
  BUFFD0 U1919 ( .I(n1934), .Z(n1933) );
  BUFFD0 U1920 ( .I(n1935), .Z(n1934) );
  BUFFD0 U1921 ( .I(n1936), .Z(n1935) );
  BUFFD0 U1922 ( .I(n1937), .Z(n1936) );
  BUFFD0 U1923 ( .I(n1938), .Z(n1937) );
  BUFFD0 U1924 ( .I(n1939), .Z(n1938) );
  BUFFD0 U1925 ( .I(n1940), .Z(n1939) );
  BUFFD0 U1926 ( .I(n1941), .Z(n1940) );
  BUFFD0 U1927 ( .I(n1942), .Z(n1941) );
  BUFFD0 U1928 ( .I(n1943), .Z(n1942) );
  BUFFD0 U1929 ( .I(n1944), .Z(n1943) );
  BUFFD0 U1930 ( .I(n1945), .Z(n1944) );
  BUFFD0 U1931 ( .I(n1946), .Z(n1945) );
  BUFFD0 U1932 ( .I(n1947), .Z(n1946) );
  BUFFD0 U1933 ( .I(n1948), .Z(n1947) );
  BUFFD0 U1934 ( .I(n1949), .Z(n1948) );
  BUFFD0 U1935 ( .I(n1950), .Z(n1949) );
  BUFFD0 U1936 ( .I(n1951), .Z(n1950) );
  BUFFD0 U1937 ( .I(n1952), .Z(n1951) );
  BUFFD0 U1938 ( .I(n1953), .Z(n1952) );
  BUFFD0 U1939 ( .I(n1954), .Z(n1953) );
  BUFFD0 U1940 ( .I(n1955), .Z(n1954) );
  BUFFD0 U1941 ( .I(n1956), .Z(n1955) );
  BUFFD0 U1942 ( .I(n1957), .Z(n1956) );
  BUFFD0 U1943 ( .I(n1958), .Z(n1957) );
  BUFFD0 U1944 ( .I(n1959), .Z(n1958) );
  BUFFD0 U1945 ( .I(n1960), .Z(n1959) );
  BUFFD0 U1946 ( .I(n1961), .Z(n1960) );
  BUFFD0 U1947 ( .I(n1962), .Z(n1961) );
  BUFFD0 U1948 ( .I(n1963), .Z(n1962) );
  BUFFD0 U1949 ( .I(n1964), .Z(n1963) );
  BUFFD0 U1950 ( .I(n1965), .Z(n1964) );
  BUFFD0 U1951 ( .I(n1966), .Z(n1965) );
  BUFFD0 U1952 ( .I(n1967), .Z(n1966) );
  BUFFD0 U1953 ( .I(n1968), .Z(n1967) );
  BUFFD0 U1954 ( .I(n1969), .Z(n1968) );
  BUFFD0 U1955 ( .I(n1970), .Z(n1969) );
  BUFFD0 U1956 ( .I(N54), .Z(n1970) );
  BUFFD0 U1957 ( .I(n1972), .Z(n1971) );
  BUFFD0 U1958 ( .I(n1973), .Z(n1972) );
  BUFFD0 U1959 ( .I(n1974), .Z(n1973) );
  BUFFD0 U1960 ( .I(n1975), .Z(n1974) );
  BUFFD0 U1961 ( .I(n1976), .Z(n1975) );
  BUFFD0 U1962 ( .I(n1977), .Z(n1976) );
  BUFFD0 U1963 ( .I(n1978), .Z(n1977) );
  BUFFD0 U1964 ( .I(n1979), .Z(n1978) );
  BUFFD0 U1965 ( .I(n1980), .Z(n1979) );
  BUFFD0 U1966 ( .I(n1981), .Z(n1980) );
  BUFFD0 U1967 ( .I(n1982), .Z(n1981) );
  BUFFD0 U1968 ( .I(n1983), .Z(n1982) );
  BUFFD0 U1969 ( .I(n1984), .Z(n1983) );
  BUFFD0 U1970 ( .I(n1985), .Z(n1984) );
  BUFFD0 U1971 ( .I(n1986), .Z(n1985) );
  BUFFD0 U1972 ( .I(n1987), .Z(n1986) );
  BUFFD0 U1973 ( .I(n1988), .Z(n1987) );
  BUFFD0 U1974 ( .I(n1989), .Z(n1988) );
  BUFFD0 U1975 ( .I(n1990), .Z(n1989) );
  BUFFD0 U1976 ( .I(n1991), .Z(n1990) );
  BUFFD0 U1977 ( .I(n1992), .Z(n1991) );
  BUFFD0 U1978 ( .I(n1993), .Z(n1992) );
  BUFFD0 U1979 ( .I(n1994), .Z(n1993) );
  BUFFD0 U1980 ( .I(n1995), .Z(n1994) );
  BUFFD0 U1981 ( .I(n1996), .Z(n1995) );
  BUFFD0 U1982 ( .I(n1997), .Z(n1996) );
  BUFFD0 U1983 ( .I(n1998), .Z(n1997) );
  BUFFD0 U1984 ( .I(n1999), .Z(n1998) );
  BUFFD0 U1985 ( .I(n2000), .Z(n1999) );
  BUFFD0 U1986 ( .I(n2001), .Z(n2000) );
  BUFFD0 U1987 ( .I(n2002), .Z(n2001) );
  BUFFD0 U1988 ( .I(n2003), .Z(n2002) );
  BUFFD0 U1989 ( .I(n2004), .Z(n2003) );
  BUFFD0 U1990 ( .I(n2005), .Z(n2004) );
  BUFFD0 U1991 ( .I(n2006), .Z(n2005) );
  BUFFD0 U1992 ( .I(n2007), .Z(n2006) );
  BUFFD0 U1993 ( .I(n2008), .Z(n2007) );
  BUFFD0 U1994 ( .I(n2009), .Z(n2008) );
  BUFFD0 U1995 ( .I(n2010), .Z(n2009) );
  BUFFD0 U1996 ( .I(n2011), .Z(n2010) );
  BUFFD0 U1997 ( .I(n2012), .Z(n2011) );
  BUFFD0 U1998 ( .I(n2013), .Z(n2012) );
  BUFFD0 U1999 ( .I(n2014), .Z(n2013) );
  BUFFD0 U2000 ( .I(n2015), .Z(n2014) );
  BUFFD0 U2001 ( .I(n2016), .Z(n2015) );
  BUFFD0 U2002 ( .I(n2017), .Z(n2016) );
  BUFFD0 U2003 ( .I(n2018), .Z(n2017) );
  BUFFD0 U2004 ( .I(n2019), .Z(n2018) );
  BUFFD0 U2005 ( .I(n2020), .Z(n2019) );
  BUFFD0 U2006 ( .I(n2021), .Z(n2020) );
  BUFFD0 U2007 ( .I(n2022), .Z(n2021) );
  BUFFD0 U2008 ( .I(n2023), .Z(n2022) );
  BUFFD0 U2009 ( .I(n2024), .Z(n2023) );
  BUFFD0 U2010 ( .I(n2025), .Z(n2024) );
  BUFFD0 U2011 ( .I(n2026), .Z(n2025) );
  BUFFD0 U2012 ( .I(n2027), .Z(n2026) );
  BUFFD0 U2013 ( .I(n2028), .Z(n2027) );
  BUFFD0 U2014 ( .I(n2029), .Z(n2028) );
  BUFFD0 U2015 ( .I(n2030), .Z(n2029) );
  BUFFD0 U2016 ( .I(n2031), .Z(n2030) );
  BUFFD0 U2017 ( .I(n2032), .Z(n2031) );
  BUFFD0 U2018 ( .I(n2033), .Z(n2032) );
  BUFFD0 U2019 ( .I(n2034), .Z(n2033) );
  BUFFD0 U2020 ( .I(n2035), .Z(n2034) );
  BUFFD0 U2021 ( .I(n2036), .Z(n2035) );
  BUFFD0 U2022 ( .I(n2037), .Z(n2036) );
  BUFFD0 U2023 ( .I(n2038), .Z(n2037) );
  BUFFD0 U2024 ( .I(n2039), .Z(n2038) );
  BUFFD0 U2025 ( .I(n2040), .Z(n2039) );
  BUFFD0 U2026 ( .I(N55), .Z(n2040) );
  BUFFD0 U2027 ( .I(n2042), .Z(n2041) );
  BUFFD0 U2028 ( .I(n2043), .Z(n2042) );
  BUFFD0 U2029 ( .I(n2044), .Z(n2043) );
  BUFFD0 U2030 ( .I(n2045), .Z(n2044) );
  BUFFD0 U2031 ( .I(n2046), .Z(n2045) );
  BUFFD0 U2032 ( .I(n2047), .Z(n2046) );
  BUFFD0 U2033 ( .I(n2048), .Z(n2047) );
  BUFFD0 U2034 ( .I(n2049), .Z(n2048) );
  BUFFD0 U2035 ( .I(n2050), .Z(n2049) );
  BUFFD0 U2036 ( .I(n2051), .Z(n2050) );
  BUFFD0 U2037 ( .I(n2052), .Z(n2051) );
  BUFFD0 U2038 ( .I(n2053), .Z(n2052) );
  BUFFD0 U2039 ( .I(n2054), .Z(n2053) );
  BUFFD0 U2040 ( .I(n2055), .Z(n2054) );
  BUFFD0 U2041 ( .I(n2056), .Z(n2055) );
  BUFFD0 U2042 ( .I(n2057), .Z(n2056) );
  BUFFD0 U2043 ( .I(n2058), .Z(n2057) );
  BUFFD0 U2044 ( .I(n2059), .Z(n2058) );
  BUFFD0 U2045 ( .I(n2060), .Z(n2059) );
  BUFFD0 U2046 ( .I(n2061), .Z(n2060) );
  BUFFD0 U2047 ( .I(n2062), .Z(n2061) );
  BUFFD0 U2048 ( .I(n2063), .Z(n2062) );
  BUFFD0 U2049 ( .I(n2064), .Z(n2063) );
  BUFFD0 U2050 ( .I(n2065), .Z(n2064) );
  BUFFD0 U2051 ( .I(n2066), .Z(n2065) );
  BUFFD0 U2052 ( .I(n2067), .Z(n2066) );
  BUFFD0 U2053 ( .I(n2068), .Z(n2067) );
  BUFFD0 U2054 ( .I(n2069), .Z(n2068) );
  BUFFD0 U2055 ( .I(n2070), .Z(n2069) );
  BUFFD0 U2056 ( .I(n2071), .Z(n2070) );
  BUFFD0 U2057 ( .I(n2072), .Z(n2071) );
  BUFFD0 U2058 ( .I(n2073), .Z(n2072) );
  BUFFD0 U2059 ( .I(n2074), .Z(n2073) );
  BUFFD0 U2060 ( .I(n2075), .Z(n2074) );
  BUFFD0 U2061 ( .I(n2076), .Z(n2075) );
  BUFFD0 U2062 ( .I(n2077), .Z(n2076) );
  BUFFD0 U2063 ( .I(n2078), .Z(n2077) );
  BUFFD0 U2064 ( .I(n2079), .Z(n2078) );
  BUFFD0 U2065 ( .I(n2080), .Z(n2079) );
  BUFFD0 U2066 ( .I(n2081), .Z(n2080) );
  BUFFD0 U2067 ( .I(n2082), .Z(n2081) );
  BUFFD0 U2068 ( .I(n2083), .Z(n2082) );
  BUFFD0 U2069 ( .I(n2084), .Z(n2083) );
  BUFFD0 U2070 ( .I(n2085), .Z(n2084) );
  BUFFD0 U2071 ( .I(n2086), .Z(n2085) );
  BUFFD0 U2072 ( .I(n2087), .Z(n2086) );
  BUFFD0 U2073 ( .I(n2088), .Z(n2087) );
  BUFFD0 U2074 ( .I(n2089), .Z(n2088) );
  BUFFD0 U2075 ( .I(n2090), .Z(n2089) );
  BUFFD0 U2076 ( .I(n2091), .Z(n2090) );
  BUFFD0 U2077 ( .I(n2092), .Z(n2091) );
  BUFFD0 U2078 ( .I(n2093), .Z(n2092) );
  BUFFD0 U2079 ( .I(n2094), .Z(n2093) );
  BUFFD0 U2080 ( .I(n2095), .Z(n2094) );
  BUFFD0 U2081 ( .I(n2096), .Z(n2095) );
  BUFFD0 U2082 ( .I(n2097), .Z(n2096) );
  BUFFD0 U2083 ( .I(n2098), .Z(n2097) );
  BUFFD0 U2084 ( .I(n2099), .Z(n2098) );
  BUFFD0 U2085 ( .I(n2100), .Z(n2099) );
  BUFFD0 U2086 ( .I(n2101), .Z(n2100) );
  BUFFD0 U2087 ( .I(n2102), .Z(n2101) );
  BUFFD0 U2088 ( .I(n2103), .Z(n2102) );
  BUFFD0 U2089 ( .I(n2104), .Z(n2103) );
  BUFFD0 U2090 ( .I(n2105), .Z(n2104) );
  BUFFD0 U2091 ( .I(n2106), .Z(n2105) );
  BUFFD0 U2092 ( .I(n2107), .Z(n2106) );
  BUFFD0 U2093 ( .I(n2108), .Z(n2107) );
  BUFFD0 U2094 ( .I(n2109), .Z(n2108) );
  BUFFD0 U2095 ( .I(n2110), .Z(n2109) );
  BUFFD0 U2096 ( .I(N56), .Z(n2110) );
  BUFFD0 U2097 ( .I(n2112), .Z(n2111) );
  BUFFD0 U2098 ( .I(n2113), .Z(n2112) );
  BUFFD0 U2099 ( .I(n2114), .Z(n2113) );
  BUFFD0 U2100 ( .I(n2115), .Z(n2114) );
  BUFFD0 U2101 ( .I(n2116), .Z(n2115) );
  BUFFD0 U2102 ( .I(n2117), .Z(n2116) );
  BUFFD0 U2103 ( .I(n2118), .Z(n2117) );
  BUFFD0 U2104 ( .I(n2119), .Z(n2118) );
  BUFFD0 U2105 ( .I(n2120), .Z(n2119) );
  BUFFD0 U2106 ( .I(n2121), .Z(n2120) );
  BUFFD0 U2107 ( .I(n2122), .Z(n2121) );
  BUFFD0 U2108 ( .I(n2123), .Z(n2122) );
  BUFFD0 U2109 ( .I(n2124), .Z(n2123) );
  BUFFD0 U2110 ( .I(n2125), .Z(n2124) );
  BUFFD0 U2111 ( .I(n2126), .Z(n2125) );
  BUFFD0 U2112 ( .I(n2127), .Z(n2126) );
  BUFFD0 U2113 ( .I(n2128), .Z(n2127) );
  BUFFD0 U2114 ( .I(n2129), .Z(n2128) );
  BUFFD0 U2115 ( .I(n2130), .Z(n2129) );
  BUFFD0 U2116 ( .I(n2131), .Z(n2130) );
  BUFFD0 U2117 ( .I(n2132), .Z(n2131) );
  BUFFD0 U2118 ( .I(n2133), .Z(n2132) );
  BUFFD0 U2119 ( .I(n2134), .Z(n2133) );
  BUFFD0 U2120 ( .I(n2135), .Z(n2134) );
  BUFFD0 U2121 ( .I(n2136), .Z(n2135) );
  BUFFD0 U2122 ( .I(n2137), .Z(n2136) );
  BUFFD0 U2123 ( .I(n2138), .Z(n2137) );
  BUFFD0 U2124 ( .I(n2139), .Z(n2138) );
  BUFFD0 U2125 ( .I(n2140), .Z(n2139) );
  BUFFD0 U2126 ( .I(n2141), .Z(n2140) );
  BUFFD0 U2127 ( .I(n2142), .Z(n2141) );
  BUFFD0 U2128 ( .I(n2143), .Z(n2142) );
  BUFFD0 U2129 ( .I(n2144), .Z(n2143) );
  BUFFD0 U2130 ( .I(n2145), .Z(n2144) );
  BUFFD0 U2131 ( .I(n2146), .Z(n2145) );
  BUFFD0 U2132 ( .I(n2147), .Z(n2146) );
  BUFFD0 U2133 ( .I(n2148), .Z(n2147) );
  BUFFD0 U2134 ( .I(n2149), .Z(n2148) );
  BUFFD0 U2135 ( .I(n2150), .Z(n2149) );
  BUFFD0 U2136 ( .I(n2151), .Z(n2150) );
  BUFFD0 U2137 ( .I(n2152), .Z(n2151) );
  BUFFD0 U2138 ( .I(n2153), .Z(n2152) );
  BUFFD0 U2139 ( .I(n2154), .Z(n2153) );
  BUFFD0 U2140 ( .I(n2155), .Z(n2154) );
  BUFFD0 U2141 ( .I(n2156), .Z(n2155) );
  BUFFD0 U2142 ( .I(n2157), .Z(n2156) );
  BUFFD0 U2143 ( .I(n2158), .Z(n2157) );
  BUFFD0 U2144 ( .I(n2159), .Z(n2158) );
  BUFFD0 U2145 ( .I(n2160), .Z(n2159) );
  BUFFD0 U2146 ( .I(n2161), .Z(n2160) );
  BUFFD0 U2147 ( .I(n2162), .Z(n2161) );
  BUFFD0 U2148 ( .I(n2163), .Z(n2162) );
  BUFFD0 U2149 ( .I(n2164), .Z(n2163) );
  BUFFD0 U2150 ( .I(n2165), .Z(n2164) );
  BUFFD0 U2151 ( .I(n2166), .Z(n2165) );
  BUFFD0 U2152 ( .I(n2167), .Z(n2166) );
  BUFFD0 U2153 ( .I(n2168), .Z(n2167) );
  BUFFD0 U2154 ( .I(n2169), .Z(n2168) );
  BUFFD0 U2155 ( .I(n2170), .Z(n2169) );
  BUFFD0 U2156 ( .I(n2171), .Z(n2170) );
  BUFFD0 U2157 ( .I(n2172), .Z(n2171) );
  BUFFD0 U2158 ( .I(n2173), .Z(n2172) );
  BUFFD0 U2159 ( .I(n2174), .Z(n2173) );
  BUFFD0 U2160 ( .I(n2175), .Z(n2174) );
  BUFFD0 U2161 ( .I(n2176), .Z(n2175) );
  BUFFD0 U2162 ( .I(n2177), .Z(n2176) );
  BUFFD0 U2163 ( .I(n2178), .Z(n2177) );
  BUFFD0 U2164 ( .I(n2179), .Z(n2178) );
  BUFFD0 U2165 ( .I(n2180), .Z(n2179) );
  BUFFD0 U2166 ( .I(N57), .Z(n2180) );
  BUFFD0 U2167 ( .I(n2182), .Z(n2181) );
  BUFFD0 U2168 ( .I(n2183), .Z(n2182) );
  BUFFD0 U2169 ( .I(n2184), .Z(n2183) );
  BUFFD0 U2170 ( .I(n2185), .Z(n2184) );
  BUFFD0 U2171 ( .I(n2186), .Z(n2185) );
  BUFFD0 U2172 ( .I(n2187), .Z(n2186) );
  BUFFD0 U2173 ( .I(n2188), .Z(n2187) );
  BUFFD0 U2174 ( .I(n2189), .Z(n2188) );
  BUFFD0 U2175 ( .I(n2190), .Z(n2189) );
  BUFFD0 U2176 ( .I(n2191), .Z(n2190) );
  BUFFD0 U2177 ( .I(n2192), .Z(n2191) );
  BUFFD0 U2178 ( .I(n2193), .Z(n2192) );
  BUFFD0 U2179 ( .I(n2194), .Z(n2193) );
  BUFFD0 U2180 ( .I(n2195), .Z(n2194) );
  BUFFD0 U2181 ( .I(n2196), .Z(n2195) );
  BUFFD0 U2182 ( .I(n2197), .Z(n2196) );
  BUFFD0 U2183 ( .I(n2198), .Z(n2197) );
  BUFFD0 U2184 ( .I(n2199), .Z(n2198) );
  BUFFD0 U2185 ( .I(n2200), .Z(n2199) );
  BUFFD0 U2186 ( .I(n2201), .Z(n2200) );
  BUFFD0 U2187 ( .I(n2202), .Z(n2201) );
  BUFFD0 U2188 ( .I(n2203), .Z(n2202) );
  BUFFD0 U2189 ( .I(n2204), .Z(n2203) );
  BUFFD0 U2190 ( .I(n2205), .Z(n2204) );
  BUFFD0 U2191 ( .I(n2206), .Z(n2205) );
  BUFFD0 U2192 ( .I(n2207), .Z(n2206) );
  BUFFD0 U2193 ( .I(n2208), .Z(n2207) );
  BUFFD0 U2194 ( .I(n2209), .Z(n2208) );
  BUFFD0 U2195 ( .I(n2210), .Z(n2209) );
  BUFFD0 U2196 ( .I(n2211), .Z(n2210) );
  BUFFD0 U2197 ( .I(n2212), .Z(n2211) );
  BUFFD0 U2198 ( .I(n2213), .Z(n2212) );
  BUFFD0 U2199 ( .I(n2214), .Z(n2213) );
  BUFFD0 U2200 ( .I(n2215), .Z(n2214) );
  BUFFD0 U2201 ( .I(n2216), .Z(n2215) );
  BUFFD0 U2202 ( .I(n2217), .Z(n2216) );
  BUFFD0 U2203 ( .I(n2218), .Z(n2217) );
  BUFFD0 U2204 ( .I(n2219), .Z(n2218) );
  BUFFD0 U2205 ( .I(n2220), .Z(n2219) );
  BUFFD0 U2206 ( .I(n2221), .Z(n2220) );
  BUFFD0 U2207 ( .I(n2222), .Z(n2221) );
  BUFFD0 U2208 ( .I(n2223), .Z(n2222) );
  BUFFD0 U2209 ( .I(n2224), .Z(n2223) );
  BUFFD0 U2210 ( .I(n2225), .Z(n2224) );
  BUFFD0 U2211 ( .I(n2226), .Z(n2225) );
  BUFFD0 U2212 ( .I(n2227), .Z(n2226) );
  BUFFD0 U2213 ( .I(n2228), .Z(n2227) );
  BUFFD0 U2214 ( .I(n2229), .Z(n2228) );
  BUFFD0 U2215 ( .I(n2230), .Z(n2229) );
  BUFFD0 U2216 ( .I(n2231), .Z(n2230) );
  BUFFD0 U2217 ( .I(n2232), .Z(n2231) );
  BUFFD0 U2218 ( .I(n2233), .Z(n2232) );
  BUFFD0 U2219 ( .I(n2234), .Z(n2233) );
  BUFFD0 U2220 ( .I(n2235), .Z(n2234) );
  BUFFD0 U2221 ( .I(n2236), .Z(n2235) );
  BUFFD0 U2222 ( .I(n2237), .Z(n2236) );
  BUFFD0 U2223 ( .I(n2238), .Z(n2237) );
  BUFFD0 U2224 ( .I(n2239), .Z(n2238) );
  BUFFD0 U2225 ( .I(n2240), .Z(n2239) );
  BUFFD0 U2226 ( .I(n2241), .Z(n2240) );
  BUFFD0 U2227 ( .I(n2242), .Z(n2241) );
  BUFFD0 U2228 ( .I(n2243), .Z(n2242) );
  BUFFD0 U2229 ( .I(n2244), .Z(n2243) );
  BUFFD0 U2230 ( .I(n2245), .Z(n2244) );
  BUFFD0 U2231 ( .I(n2246), .Z(n2245) );
  BUFFD0 U2232 ( .I(n2247), .Z(n2246) );
  BUFFD0 U2233 ( .I(n2248), .Z(n2247) );
  BUFFD0 U2234 ( .I(n2249), .Z(n2248) );
  BUFFD0 U2235 ( .I(n2250), .Z(n2249) );
  BUFFD0 U2236 ( .I(N58), .Z(n2250) );
  BUFFD0 U2237 ( .I(n2252), .Z(n2251) );
  BUFFD0 U2238 ( .I(n2253), .Z(n2252) );
  BUFFD0 U2239 ( .I(n2254), .Z(n2253) );
  BUFFD0 U2240 ( .I(n2255), .Z(n2254) );
  BUFFD0 U2241 ( .I(n2256), .Z(n2255) );
  BUFFD0 U2242 ( .I(n2257), .Z(n2256) );
  BUFFD0 U2243 ( .I(n2258), .Z(n2257) );
  BUFFD0 U2244 ( .I(n2259), .Z(n2258) );
  BUFFD0 U2245 ( .I(n2260), .Z(n2259) );
  BUFFD0 U2246 ( .I(n2261), .Z(n2260) );
  BUFFD0 U2247 ( .I(n2262), .Z(n2261) );
  BUFFD0 U2248 ( .I(n2263), .Z(n2262) );
  BUFFD0 U2249 ( .I(n2264), .Z(n2263) );
  BUFFD0 U2250 ( .I(n2265), .Z(n2264) );
  BUFFD0 U2251 ( .I(n2266), .Z(n2265) );
  BUFFD0 U2252 ( .I(n2267), .Z(n2266) );
  BUFFD0 U2253 ( .I(n2268), .Z(n2267) );
  BUFFD0 U2254 ( .I(n2269), .Z(n2268) );
  BUFFD0 U2255 ( .I(n2270), .Z(n2269) );
  BUFFD0 U2256 ( .I(n2271), .Z(n2270) );
  BUFFD0 U2257 ( .I(n2272), .Z(n2271) );
  BUFFD0 U2258 ( .I(n2273), .Z(n2272) );
  BUFFD0 U2259 ( .I(n2274), .Z(n2273) );
  BUFFD0 U2260 ( .I(n2275), .Z(n2274) );
  BUFFD0 U2261 ( .I(n2276), .Z(n2275) );
  BUFFD0 U2262 ( .I(n2277), .Z(n2276) );
  BUFFD0 U2263 ( .I(n2278), .Z(n2277) );
  BUFFD0 U2264 ( .I(n2279), .Z(n2278) );
  BUFFD0 U2265 ( .I(n2280), .Z(n2279) );
  BUFFD0 U2266 ( .I(n2281), .Z(n2280) );
  BUFFD0 U2267 ( .I(n2282), .Z(n2281) );
  BUFFD0 U2268 ( .I(n2283), .Z(n2282) );
  BUFFD0 U2269 ( .I(n2284), .Z(n2283) );
  BUFFD0 U2270 ( .I(n2285), .Z(n2284) );
  BUFFD0 U2271 ( .I(n2286), .Z(n2285) );
  BUFFD0 U2272 ( .I(n2287), .Z(n2286) );
  BUFFD0 U2273 ( .I(n2288), .Z(n2287) );
  BUFFD0 U2274 ( .I(n2289), .Z(n2288) );
  BUFFD0 U2275 ( .I(n2290), .Z(n2289) );
  BUFFD0 U2276 ( .I(n2291), .Z(n2290) );
  BUFFD0 U2277 ( .I(n2292), .Z(n2291) );
  BUFFD0 U2278 ( .I(n2293), .Z(n2292) );
  BUFFD0 U2279 ( .I(n2294), .Z(n2293) );
  BUFFD0 U2280 ( .I(n2295), .Z(n2294) );
  BUFFD0 U2281 ( .I(n2296), .Z(n2295) );
  BUFFD0 U2282 ( .I(n2297), .Z(n2296) );
  BUFFD0 U2283 ( .I(n2298), .Z(n2297) );
  BUFFD0 U2284 ( .I(n2299), .Z(n2298) );
  BUFFD0 U2285 ( .I(n2300), .Z(n2299) );
  BUFFD0 U2286 ( .I(n2301), .Z(n2300) );
  BUFFD0 U2287 ( .I(n2302), .Z(n2301) );
  BUFFD0 U2288 ( .I(n2303), .Z(n2302) );
  BUFFD0 U2289 ( .I(n2304), .Z(n2303) );
  BUFFD0 U2290 ( .I(n2305), .Z(n2304) );
  BUFFD0 U2291 ( .I(n2306), .Z(n2305) );
  BUFFD0 U2292 ( .I(n2307), .Z(n2306) );
  BUFFD0 U2293 ( .I(n2308), .Z(n2307) );
  BUFFD0 U2294 ( .I(n2309), .Z(n2308) );
  BUFFD0 U2295 ( .I(n2310), .Z(n2309) );
  BUFFD0 U2296 ( .I(n2311), .Z(n2310) );
  BUFFD0 U2297 ( .I(n2312), .Z(n2311) );
  BUFFD0 U2298 ( .I(n2313), .Z(n2312) );
  BUFFD0 U2299 ( .I(n2314), .Z(n2313) );
  BUFFD0 U2300 ( .I(n2315), .Z(n2314) );
  BUFFD0 U2301 ( .I(n2316), .Z(n2315) );
  BUFFD0 U2302 ( .I(n2317), .Z(n2316) );
  BUFFD0 U2303 ( .I(n2318), .Z(n2317) );
  BUFFD0 U2304 ( .I(n2319), .Z(n2318) );
  BUFFD0 U2305 ( .I(n2320), .Z(n2319) );
  BUFFD0 U2306 ( .I(N59), .Z(n2320) );
  BUFFD0 U2307 ( .I(n2322), .Z(n2321) );
  BUFFD0 U2308 ( .I(n2323), .Z(n2322) );
  BUFFD0 U2309 ( .I(n2324), .Z(n2323) );
  BUFFD0 U2310 ( .I(n2325), .Z(n2324) );
  BUFFD0 U2311 ( .I(n2326), .Z(n2325) );
  BUFFD0 U2312 ( .I(n2327), .Z(n2326) );
  BUFFD0 U2313 ( .I(n2328), .Z(n2327) );
  BUFFD0 U2314 ( .I(n2329), .Z(n2328) );
  BUFFD0 U2315 ( .I(n2330), .Z(n2329) );
  BUFFD0 U2316 ( .I(n2331), .Z(n2330) );
  BUFFD0 U2317 ( .I(n2332), .Z(n2331) );
  BUFFD0 U2318 ( .I(n2333), .Z(n2332) );
  BUFFD0 U2319 ( .I(n2334), .Z(n2333) );
  BUFFD0 U2320 ( .I(n2335), .Z(n2334) );
  BUFFD0 U2321 ( .I(n2336), .Z(n2335) );
  BUFFD0 U2322 ( .I(n2337), .Z(n2336) );
  BUFFD0 U2323 ( .I(n2338), .Z(n2337) );
  BUFFD0 U2324 ( .I(n2339), .Z(n2338) );
  BUFFD0 U2325 ( .I(n2340), .Z(n2339) );
  BUFFD0 U2326 ( .I(n2341), .Z(n2340) );
  BUFFD0 U2327 ( .I(n2342), .Z(n2341) );
  BUFFD0 U2328 ( .I(n2343), .Z(n2342) );
  BUFFD0 U2329 ( .I(n2344), .Z(n2343) );
  BUFFD0 U2330 ( .I(n2345), .Z(n2344) );
  BUFFD0 U2331 ( .I(n2346), .Z(n2345) );
  BUFFD0 U2332 ( .I(n2347), .Z(n2346) );
  BUFFD0 U2333 ( .I(n2348), .Z(n2347) );
  BUFFD0 U2334 ( .I(n2349), .Z(n2348) );
  BUFFD0 U2335 ( .I(n2350), .Z(n2349) );
  BUFFD0 U2336 ( .I(n2351), .Z(n2350) );
  BUFFD0 U2337 ( .I(n2352), .Z(n2351) );
  BUFFD0 U2338 ( .I(n2353), .Z(n2352) );
  BUFFD0 U2339 ( .I(n2354), .Z(n2353) );
  BUFFD0 U2340 ( .I(n2355), .Z(n2354) );
  BUFFD0 U2341 ( .I(n2356), .Z(n2355) );
  BUFFD0 U2342 ( .I(n2357), .Z(n2356) );
  BUFFD0 U2343 ( .I(n2358), .Z(n2357) );
  BUFFD0 U2344 ( .I(n2359), .Z(n2358) );
  BUFFD0 U2345 ( .I(n2360), .Z(n2359) );
  BUFFD0 U2346 ( .I(n2361), .Z(n2360) );
  BUFFD0 U2347 ( .I(n2362), .Z(n2361) );
  BUFFD0 U2348 ( .I(n2363), .Z(n2362) );
  BUFFD0 U2349 ( .I(n2364), .Z(n2363) );
  BUFFD0 U2350 ( .I(n2365), .Z(n2364) );
  BUFFD0 U2351 ( .I(n2366), .Z(n2365) );
  BUFFD0 U2352 ( .I(n2367), .Z(n2366) );
  BUFFD0 U2353 ( .I(n2368), .Z(n2367) );
  BUFFD0 U2354 ( .I(n2369), .Z(n2368) );
  BUFFD0 U2355 ( .I(n2370), .Z(n2369) );
  BUFFD0 U2356 ( .I(n2371), .Z(n2370) );
  BUFFD0 U2357 ( .I(n2372), .Z(n2371) );
  BUFFD0 U2358 ( .I(n2373), .Z(n2372) );
  BUFFD0 U2359 ( .I(n2374), .Z(n2373) );
  BUFFD0 U2360 ( .I(n2375), .Z(n2374) );
  BUFFD0 U2361 ( .I(n2376), .Z(n2375) );
  BUFFD0 U2362 ( .I(n2377), .Z(n2376) );
  BUFFD0 U2363 ( .I(n2378), .Z(n2377) );
  BUFFD0 U2364 ( .I(n2379), .Z(n2378) );
  BUFFD0 U2365 ( .I(n2380), .Z(n2379) );
  BUFFD0 U2366 ( .I(n2381), .Z(n2380) );
  BUFFD0 U2367 ( .I(n2382), .Z(n2381) );
  BUFFD0 U2368 ( .I(n2383), .Z(n2382) );
  BUFFD0 U2369 ( .I(n2384), .Z(n2383) );
  BUFFD0 U2370 ( .I(n2385), .Z(n2384) );
  BUFFD0 U2371 ( .I(n2386), .Z(n2385) );
  BUFFD0 U2372 ( .I(n2387), .Z(n2386) );
  BUFFD0 U2373 ( .I(n2388), .Z(n2387) );
  BUFFD0 U2374 ( .I(n2389), .Z(n2388) );
  BUFFD0 U2375 ( .I(n2390), .Z(n2389) );
  BUFFD0 U2376 ( .I(N60), .Z(n2390) );
  BUFFD0 U2377 ( .I(n2392), .Z(n2391) );
  BUFFD0 U2378 ( .I(n2393), .Z(n2392) );
  BUFFD0 U2379 ( .I(n2394), .Z(n2393) );
  BUFFD0 U2380 ( .I(n2395), .Z(n2394) );
  BUFFD0 U2381 ( .I(n2396), .Z(n2395) );
  BUFFD0 U2382 ( .I(n2397), .Z(n2396) );
  BUFFD0 U2383 ( .I(n2398), .Z(n2397) );
  BUFFD0 U2384 ( .I(n2399), .Z(n2398) );
  BUFFD0 U2385 ( .I(n2400), .Z(n2399) );
  BUFFD0 U2386 ( .I(n2401), .Z(n2400) );
  BUFFD0 U2387 ( .I(n2402), .Z(n2401) );
  BUFFD0 U2388 ( .I(n2403), .Z(n2402) );
  BUFFD0 U2389 ( .I(n2404), .Z(n2403) );
  BUFFD0 U2390 ( .I(n2405), .Z(n2404) );
  BUFFD0 U2391 ( .I(n2406), .Z(n2405) );
  BUFFD0 U2392 ( .I(n2407), .Z(n2406) );
  BUFFD0 U2393 ( .I(n2408), .Z(n2407) );
  BUFFD0 U2394 ( .I(n2409), .Z(n2408) );
  BUFFD0 U2395 ( .I(n2410), .Z(n2409) );
  BUFFD0 U2396 ( .I(n2411), .Z(n2410) );
  BUFFD0 U2397 ( .I(n2412), .Z(n2411) );
  BUFFD0 U2398 ( .I(n2413), .Z(n2412) );
  BUFFD0 U2399 ( .I(n2414), .Z(n2413) );
  BUFFD0 U2400 ( .I(n2415), .Z(n2414) );
  BUFFD0 U2401 ( .I(n2416), .Z(n2415) );
  BUFFD0 U2402 ( .I(n2417), .Z(n2416) );
  BUFFD0 U2403 ( .I(n2418), .Z(n2417) );
  BUFFD0 U2404 ( .I(n2419), .Z(n2418) );
  BUFFD0 U2405 ( .I(n2420), .Z(n2419) );
  BUFFD0 U2406 ( .I(n2421), .Z(n2420) );
  BUFFD0 U2407 ( .I(n2422), .Z(n2421) );
  BUFFD0 U2408 ( .I(n2423), .Z(n2422) );
  BUFFD0 U2409 ( .I(n2424), .Z(n2423) );
  BUFFD0 U2410 ( .I(n2425), .Z(n2424) );
  BUFFD0 U2411 ( .I(n2426), .Z(n2425) );
  BUFFD0 U2412 ( .I(n2427), .Z(n2426) );
  BUFFD0 U2413 ( .I(n2428), .Z(n2427) );
  BUFFD0 U2414 ( .I(n2429), .Z(n2428) );
  BUFFD0 U2415 ( .I(n2430), .Z(n2429) );
  BUFFD0 U2416 ( .I(n2431), .Z(n2430) );
  BUFFD0 U2417 ( .I(n2432), .Z(n2431) );
  BUFFD0 U2418 ( .I(n2433), .Z(n2432) );
  BUFFD0 U2419 ( .I(n2434), .Z(n2433) );
  BUFFD0 U2420 ( .I(n2435), .Z(n2434) );
  BUFFD0 U2421 ( .I(n2436), .Z(n2435) );
  BUFFD0 U2422 ( .I(n2437), .Z(n2436) );
  BUFFD0 U2423 ( .I(n2438), .Z(n2437) );
  BUFFD0 U2424 ( .I(n2439), .Z(n2438) );
  BUFFD0 U2425 ( .I(n2440), .Z(n2439) );
  BUFFD0 U2426 ( .I(n2441), .Z(n2440) );
  BUFFD0 U2427 ( .I(n2442), .Z(n2441) );
  BUFFD0 U2428 ( .I(n2443), .Z(n2442) );
  BUFFD0 U2429 ( .I(n2444), .Z(n2443) );
  BUFFD0 U2430 ( .I(n2445), .Z(n2444) );
  BUFFD0 U2431 ( .I(n2446), .Z(n2445) );
  BUFFD0 U2432 ( .I(n2447), .Z(n2446) );
  BUFFD0 U2433 ( .I(n2448), .Z(n2447) );
  BUFFD0 U2434 ( .I(n2449), .Z(n2448) );
  BUFFD0 U2435 ( .I(n2450), .Z(n2449) );
  BUFFD0 U2436 ( .I(n2451), .Z(n2450) );
  BUFFD0 U2437 ( .I(n2452), .Z(n2451) );
  BUFFD0 U2438 ( .I(n2453), .Z(n2452) );
  BUFFD0 U2439 ( .I(n2454), .Z(n2453) );
  BUFFD0 U2440 ( .I(n2455), .Z(n2454) );
  BUFFD0 U2441 ( .I(n2456), .Z(n2455) );
  BUFFD0 U2442 ( .I(n2457), .Z(n2456) );
  BUFFD0 U2443 ( .I(n2458), .Z(n2457) );
  BUFFD0 U2444 ( .I(n2459), .Z(n2458) );
  BUFFD0 U2445 ( .I(n2460), .Z(n2459) );
  BUFFD0 U2446 ( .I(N61), .Z(n2460) );
  BUFFD0 U2447 ( .I(n2462), .Z(n2461) );
  BUFFD0 U2448 ( .I(n2463), .Z(n2462) );
  BUFFD0 U2449 ( .I(n2464), .Z(n2463) );
  BUFFD0 U2450 ( .I(n2465), .Z(n2464) );
  BUFFD0 U2451 ( .I(n2466), .Z(n2465) );
  BUFFD0 U2452 ( .I(n2467), .Z(n2466) );
  BUFFD0 U2453 ( .I(n2468), .Z(n2467) );
  BUFFD0 U2454 ( .I(n2469), .Z(n2468) );
  BUFFD0 U2455 ( .I(n2470), .Z(n2469) );
  BUFFD0 U2456 ( .I(n2471), .Z(n2470) );
  BUFFD0 U2457 ( .I(n2472), .Z(n2471) );
  BUFFD0 U2458 ( .I(n2473), .Z(n2472) );
  BUFFD0 U2459 ( .I(n2474), .Z(n2473) );
  BUFFD0 U2460 ( .I(n2475), .Z(n2474) );
  BUFFD0 U2461 ( .I(n2476), .Z(n2475) );
  BUFFD0 U2462 ( .I(n2477), .Z(n2476) );
  BUFFD0 U2463 ( .I(n2478), .Z(n2477) );
  BUFFD0 U2464 ( .I(n2479), .Z(n2478) );
  BUFFD0 U2465 ( .I(n2480), .Z(n2479) );
  BUFFD0 U2466 ( .I(n2481), .Z(n2480) );
  BUFFD0 U2467 ( .I(n2482), .Z(n2481) );
  BUFFD0 U2468 ( .I(n2483), .Z(n2482) );
  BUFFD0 U2469 ( .I(n2484), .Z(n2483) );
  BUFFD0 U2470 ( .I(n2485), .Z(n2484) );
  BUFFD0 U2471 ( .I(n2486), .Z(n2485) );
  BUFFD0 U2472 ( .I(n2487), .Z(n2486) );
  BUFFD0 U2473 ( .I(n2488), .Z(n2487) );
  BUFFD0 U2474 ( .I(n2489), .Z(n2488) );
  BUFFD0 U2475 ( .I(n2490), .Z(n2489) );
  BUFFD0 U2476 ( .I(n2491), .Z(n2490) );
  BUFFD0 U2477 ( .I(n2492), .Z(n2491) );
  BUFFD0 U2478 ( .I(n2493), .Z(n2492) );
  BUFFD0 U2479 ( .I(n2494), .Z(n2493) );
  BUFFD0 U2480 ( .I(n2495), .Z(n2494) );
  BUFFD0 U2481 ( .I(n2496), .Z(n2495) );
  BUFFD0 U2482 ( .I(n2497), .Z(n2496) );
  BUFFD0 U2483 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2484 ( .I(n2499), .Z(n2498) );
  BUFFD0 U2485 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2486 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2487 ( .I(n2502), .Z(n2501) );
  BUFFD0 U2488 ( .I(n2503), .Z(n2502) );
  BUFFD0 U2489 ( .I(n2504), .Z(n2503) );
  BUFFD0 U2490 ( .I(n2505), .Z(n2504) );
  BUFFD0 U2491 ( .I(n2506), .Z(n2505) );
  BUFFD0 U2492 ( .I(n2507), .Z(n2506) );
  BUFFD0 U2493 ( .I(n2508), .Z(n2507) );
  BUFFD0 U2494 ( .I(n2509), .Z(n2508) );
  BUFFD0 U2495 ( .I(n2510), .Z(n2509) );
  BUFFD0 U2496 ( .I(n2511), .Z(n2510) );
  BUFFD0 U2497 ( .I(n2512), .Z(n2511) );
  BUFFD0 U2498 ( .I(n2513), .Z(n2512) );
  BUFFD0 U2499 ( .I(n2514), .Z(n2513) );
  BUFFD0 U2500 ( .I(n2515), .Z(n2514) );
  BUFFD0 U2501 ( .I(n2516), .Z(n2515) );
  BUFFD0 U2502 ( .I(n2517), .Z(n2516) );
  BUFFD0 U2503 ( .I(n2518), .Z(n2517) );
  BUFFD0 U2504 ( .I(n2519), .Z(n2518) );
  BUFFD0 U2505 ( .I(n2520), .Z(n2519) );
  BUFFD0 U2506 ( .I(n2521), .Z(n2520) );
  BUFFD0 U2507 ( .I(n2522), .Z(n2521) );
  BUFFD0 U2508 ( .I(n2523), .Z(n2522) );
  BUFFD0 U2509 ( .I(n2524), .Z(n2523) );
  BUFFD0 U2510 ( .I(n2525), .Z(n2524) );
  BUFFD0 U2511 ( .I(n2526), .Z(n2525) );
  BUFFD0 U2512 ( .I(n2527), .Z(n2526) );
  BUFFD0 U2513 ( .I(n2528), .Z(n2527) );
  BUFFD0 U2514 ( .I(n2529), .Z(n2528) );
  BUFFD0 U2515 ( .I(n2530), .Z(n2529) );
  BUFFD0 U2516 ( .I(N62), .Z(n2530) );
  BUFFD0 U2517 ( .I(n2532), .Z(n2531) );
  BUFFD0 U2518 ( .I(n2533), .Z(n2532) );
  BUFFD0 U2519 ( .I(n2534), .Z(n2533) );
  BUFFD0 U2520 ( .I(n2535), .Z(n2534) );
  BUFFD0 U2521 ( .I(n2536), .Z(n2535) );
  BUFFD0 U2522 ( .I(n2537), .Z(n2536) );
  BUFFD0 U2523 ( .I(n2538), .Z(n2537) );
  BUFFD0 U2524 ( .I(n2539), .Z(n2538) );
  BUFFD0 U2525 ( .I(n2540), .Z(n2539) );
  BUFFD0 U2526 ( .I(n2541), .Z(n2540) );
  BUFFD0 U2527 ( .I(n2542), .Z(n2541) );
  BUFFD0 U2528 ( .I(n2543), .Z(n2542) );
  BUFFD0 U2529 ( .I(n2544), .Z(n2543) );
  BUFFD0 U2530 ( .I(n2545), .Z(n2544) );
  BUFFD0 U2531 ( .I(n2546), .Z(n2545) );
  BUFFD0 U2532 ( .I(n2547), .Z(n2546) );
  BUFFD0 U2533 ( .I(n2548), .Z(n2547) );
  BUFFD0 U2534 ( .I(n2549), .Z(n2548) );
  BUFFD0 U2535 ( .I(n2550), .Z(n2549) );
  BUFFD0 U2536 ( .I(n2551), .Z(n2550) );
  BUFFD0 U2537 ( .I(n2552), .Z(n2551) );
  BUFFD0 U2538 ( .I(n2553), .Z(n2552) );
  BUFFD0 U2539 ( .I(n2554), .Z(n2553) );
  BUFFD0 U2540 ( .I(n2555), .Z(n2554) );
  BUFFD0 U2541 ( .I(n2556), .Z(n2555) );
  BUFFD0 U2542 ( .I(n2557), .Z(n2556) );
  BUFFD0 U2543 ( .I(n2558), .Z(n2557) );
  BUFFD0 U2544 ( .I(n2559), .Z(n2558) );
  BUFFD0 U2545 ( .I(n2560), .Z(n2559) );
  BUFFD0 U2546 ( .I(n2561), .Z(n2560) );
  BUFFD0 U2547 ( .I(n2562), .Z(n2561) );
  BUFFD0 U2548 ( .I(n2563), .Z(n2562) );
  BUFFD0 U2549 ( .I(n2564), .Z(n2563) );
  BUFFD0 U2550 ( .I(n2565), .Z(n2564) );
  BUFFD0 U2551 ( .I(n2566), .Z(n2565) );
  BUFFD0 U2552 ( .I(n2567), .Z(n2566) );
  BUFFD0 U2553 ( .I(n2568), .Z(n2567) );
  BUFFD0 U2554 ( .I(n2569), .Z(n2568) );
  BUFFD0 U2555 ( .I(n2570), .Z(n2569) );
  BUFFD0 U2556 ( .I(n2571), .Z(n2570) );
  BUFFD0 U2557 ( .I(n2572), .Z(n2571) );
  BUFFD0 U2558 ( .I(n2573), .Z(n2572) );
  BUFFD0 U2559 ( .I(n2574), .Z(n2573) );
  BUFFD0 U2560 ( .I(n2575), .Z(n2574) );
  BUFFD0 U2561 ( .I(n2576), .Z(n2575) );
  BUFFD0 U2562 ( .I(n2577), .Z(n2576) );
  BUFFD0 U2563 ( .I(n2578), .Z(n2577) );
  BUFFD0 U2564 ( .I(n2579), .Z(n2578) );
  BUFFD0 U2565 ( .I(n2580), .Z(n2579) );
  BUFFD0 U2566 ( .I(n2581), .Z(n2580) );
  BUFFD0 U2567 ( .I(n2582), .Z(n2581) );
  BUFFD0 U2568 ( .I(n2583), .Z(n2582) );
  BUFFD0 U2569 ( .I(n2584), .Z(n2583) );
  BUFFD0 U2570 ( .I(n2585), .Z(n2584) );
  BUFFD0 U2571 ( .I(n2586), .Z(n2585) );
  BUFFD0 U2572 ( .I(n2587), .Z(n2586) );
  BUFFD0 U2573 ( .I(n2588), .Z(n2587) );
  BUFFD0 U2574 ( .I(n2589), .Z(n2588) );
  BUFFD0 U2575 ( .I(n2590), .Z(n2589) );
  BUFFD0 U2576 ( .I(n2591), .Z(n2590) );
  BUFFD0 U2577 ( .I(n2592), .Z(n2591) );
  BUFFD0 U2578 ( .I(n2593), .Z(n2592) );
  BUFFD0 U2579 ( .I(n2594), .Z(n2593) );
  BUFFD0 U2580 ( .I(n2595), .Z(n2594) );
  BUFFD0 U2581 ( .I(n2596), .Z(n2595) );
  BUFFD0 U2582 ( .I(n2597), .Z(n2596) );
  BUFFD0 U2583 ( .I(n2598), .Z(n2597) );
  BUFFD0 U2584 ( .I(n2599), .Z(n2598) );
  BUFFD0 U2585 ( .I(n2600), .Z(n2599) );
  BUFFD0 U2586 ( .I(N63), .Z(n2600) );
  BUFFD0 U2587 ( .I(n2602), .Z(n2601) );
  BUFFD0 U2588 ( .I(n2603), .Z(n2602) );
  BUFFD0 U2589 ( .I(n2604), .Z(n2603) );
  BUFFD0 U2590 ( .I(n2605), .Z(n2604) );
  BUFFD0 U2591 ( .I(n2606), .Z(n2605) );
  BUFFD0 U2592 ( .I(n2607), .Z(n2606) );
  BUFFD0 U2593 ( .I(n2608), .Z(n2607) );
  BUFFD0 U2594 ( .I(n2609), .Z(n2608) );
  BUFFD0 U2595 ( .I(n2610), .Z(n2609) );
  BUFFD0 U2596 ( .I(n2611), .Z(n2610) );
  BUFFD0 U2597 ( .I(n2612), .Z(n2611) );
  BUFFD0 U2598 ( .I(n2613), .Z(n2612) );
  BUFFD0 U2599 ( .I(n2614), .Z(n2613) );
  BUFFD0 U2600 ( .I(n2615), .Z(n2614) );
  BUFFD0 U2601 ( .I(n2616), .Z(n2615) );
  BUFFD0 U2602 ( .I(n2617), .Z(n2616) );
  BUFFD0 U2603 ( .I(n2618), .Z(n2617) );
  BUFFD0 U2604 ( .I(n2619), .Z(n2618) );
  BUFFD0 U2605 ( .I(n2620), .Z(n2619) );
  BUFFD0 U2606 ( .I(n2621), .Z(n2620) );
  BUFFD0 U2607 ( .I(n2622), .Z(n2621) );
  BUFFD0 U2608 ( .I(n2623), .Z(n2622) );
  BUFFD0 U2609 ( .I(n2624), .Z(n2623) );
  BUFFD0 U2610 ( .I(n2625), .Z(n2624) );
  BUFFD0 U2611 ( .I(n2626), .Z(n2625) );
  BUFFD0 U2612 ( .I(n2627), .Z(n2626) );
  BUFFD0 U2613 ( .I(n2628), .Z(n2627) );
  BUFFD0 U2614 ( .I(n2629), .Z(n2628) );
  BUFFD0 U2615 ( .I(n2630), .Z(n2629) );
  BUFFD0 U2616 ( .I(n2631), .Z(n2630) );
  BUFFD0 U2617 ( .I(n2632), .Z(n2631) );
  BUFFD0 U2618 ( .I(n2633), .Z(n2632) );
  BUFFD0 U2619 ( .I(n2634), .Z(n2633) );
  BUFFD0 U2620 ( .I(n2635), .Z(n2634) );
  BUFFD0 U2621 ( .I(n2636), .Z(n2635) );
  BUFFD0 U2622 ( .I(n2637), .Z(n2636) );
  BUFFD0 U2623 ( .I(n2638), .Z(n2637) );
  BUFFD0 U2624 ( .I(n2639), .Z(n2638) );
  BUFFD0 U2625 ( .I(n2640), .Z(n2639) );
  BUFFD0 U2626 ( .I(n2641), .Z(n2640) );
  BUFFD0 U2627 ( .I(n2642), .Z(n2641) );
  BUFFD0 U2628 ( .I(n2643), .Z(n2642) );
  BUFFD0 U2629 ( .I(n2644), .Z(n2643) );
  BUFFD0 U2630 ( .I(n2645), .Z(n2644) );
  BUFFD0 U2631 ( .I(n2646), .Z(n2645) );
  BUFFD0 U2632 ( .I(n2647), .Z(n2646) );
  BUFFD0 U2633 ( .I(n2648), .Z(n2647) );
  BUFFD0 U2634 ( .I(n2649), .Z(n2648) );
  BUFFD0 U2635 ( .I(n2650), .Z(n2649) );
  BUFFD0 U2636 ( .I(n2651), .Z(n2650) );
  BUFFD0 U2637 ( .I(n2652), .Z(n2651) );
  BUFFD0 U2638 ( .I(n2653), .Z(n2652) );
  BUFFD0 U2639 ( .I(n2654), .Z(n2653) );
  BUFFD0 U2640 ( .I(n2655), .Z(n2654) );
  BUFFD0 U2641 ( .I(n2656), .Z(n2655) );
  BUFFD0 U2642 ( .I(n2657), .Z(n2656) );
  BUFFD0 U2643 ( .I(n2658), .Z(n2657) );
  BUFFD0 U2644 ( .I(n2659), .Z(n2658) );
  BUFFD0 U2645 ( .I(n2660), .Z(n2659) );
  BUFFD0 U2646 ( .I(n2661), .Z(n2660) );
  BUFFD0 U2647 ( .I(n2662), .Z(n2661) );
  BUFFD0 U2648 ( .I(n2663), .Z(n2662) );
  BUFFD0 U2649 ( .I(n2664), .Z(n2663) );
  BUFFD0 U2650 ( .I(n2665), .Z(n2664) );
  BUFFD0 U2651 ( .I(n2666), .Z(n2665) );
  BUFFD0 U2652 ( .I(n2667), .Z(n2666) );
  BUFFD0 U2653 ( .I(n2668), .Z(n2667) );
  BUFFD0 U2654 ( .I(n2669), .Z(n2668) );
  BUFFD0 U2655 ( .I(n2670), .Z(n2669) );
  BUFFD0 U2656 ( .I(N64), .Z(n2670) );
  BUFFD0 U2657 ( .I(n2672), .Z(n2671) );
  BUFFD0 U2658 ( .I(n2673), .Z(n2672) );
  BUFFD0 U2659 ( .I(n2674), .Z(n2673) );
  BUFFD0 U2660 ( .I(n2675), .Z(n2674) );
  BUFFD0 U2661 ( .I(n2676), .Z(n2675) );
  BUFFD0 U2662 ( .I(n2677), .Z(n2676) );
  BUFFD0 U2663 ( .I(n2678), .Z(n2677) );
  BUFFD0 U2664 ( .I(n2679), .Z(n2678) );
  BUFFD0 U2665 ( .I(n2680), .Z(n2679) );
  BUFFD0 U2666 ( .I(n2681), .Z(n2680) );
  BUFFD0 U2667 ( .I(n2682), .Z(n2681) );
  BUFFD0 U2668 ( .I(n2683), .Z(n2682) );
  BUFFD0 U2669 ( .I(n2684), .Z(n2683) );
  BUFFD0 U2670 ( .I(n2685), .Z(n2684) );
  BUFFD0 U2671 ( .I(n2686), .Z(n2685) );
  BUFFD0 U2672 ( .I(n2687), .Z(n2686) );
  BUFFD0 U2673 ( .I(n2688), .Z(n2687) );
  BUFFD0 U2674 ( .I(n2689), .Z(n2688) );
  BUFFD0 U2675 ( .I(n2690), .Z(n2689) );
  BUFFD0 U2676 ( .I(n2691), .Z(n2690) );
  BUFFD0 U2677 ( .I(n2692), .Z(n2691) );
  BUFFD0 U2678 ( .I(n2693), .Z(n2692) );
  BUFFD0 U2679 ( .I(n2694), .Z(n2693) );
  BUFFD0 U2680 ( .I(n2695), .Z(n2694) );
  BUFFD0 U2681 ( .I(n2696), .Z(n2695) );
  BUFFD0 U2682 ( .I(n2697), .Z(n2696) );
  BUFFD0 U2683 ( .I(n2698), .Z(n2697) );
  BUFFD0 U2684 ( .I(n2699), .Z(n2698) );
  BUFFD0 U2685 ( .I(n2700), .Z(n2699) );
  BUFFD0 U2686 ( .I(n2701), .Z(n2700) );
  BUFFD0 U2687 ( .I(n2702), .Z(n2701) );
  BUFFD0 U2688 ( .I(n2703), .Z(n2702) );
  BUFFD0 U2689 ( .I(n2704), .Z(n2703) );
  BUFFD0 U2690 ( .I(n2705), .Z(n2704) );
  BUFFD0 U2691 ( .I(n2706), .Z(n2705) );
  BUFFD0 U2692 ( .I(n2707), .Z(n2706) );
  BUFFD0 U2693 ( .I(n2708), .Z(n2707) );
  BUFFD0 U2694 ( .I(n2709), .Z(n2708) );
  BUFFD0 U2695 ( .I(n2710), .Z(n2709) );
  BUFFD0 U2696 ( .I(n2711), .Z(n2710) );
  BUFFD0 U2697 ( .I(n2712), .Z(n2711) );
  BUFFD0 U2698 ( .I(n2713), .Z(n2712) );
  BUFFD0 U2699 ( .I(n2714), .Z(n2713) );
  BUFFD0 U2700 ( .I(n2715), .Z(n2714) );
  BUFFD0 U2701 ( .I(n2716), .Z(n2715) );
  BUFFD0 U2702 ( .I(n2717), .Z(n2716) );
  BUFFD0 U2703 ( .I(n2718), .Z(n2717) );
  BUFFD0 U2704 ( .I(n2719), .Z(n2718) );
  BUFFD0 U2705 ( .I(n2720), .Z(n2719) );
  BUFFD0 U2706 ( .I(n2721), .Z(n2720) );
  BUFFD0 U2707 ( .I(n2722), .Z(n2721) );
  BUFFD0 U2708 ( .I(n2723), .Z(n2722) );
  BUFFD0 U2709 ( .I(n2724), .Z(n2723) );
  BUFFD0 U2710 ( .I(n2725), .Z(n2724) );
  BUFFD0 U2711 ( .I(n2726), .Z(n2725) );
  BUFFD0 U2712 ( .I(n2727), .Z(n2726) );
  BUFFD0 U2713 ( .I(n2728), .Z(n2727) );
  BUFFD0 U2714 ( .I(n2729), .Z(n2728) );
  BUFFD0 U2715 ( .I(n2730), .Z(n2729) );
  BUFFD0 U2716 ( .I(n2731), .Z(n2730) );
  BUFFD0 U2717 ( .I(n2732), .Z(n2731) );
  BUFFD0 U2718 ( .I(n2733), .Z(n2732) );
  BUFFD0 U2719 ( .I(n2734), .Z(n2733) );
  BUFFD0 U2720 ( .I(n2735), .Z(n2734) );
  BUFFD0 U2721 ( .I(n2736), .Z(n2735) );
  BUFFD0 U2722 ( .I(n2737), .Z(n2736) );
  BUFFD0 U2723 ( .I(n2738), .Z(n2737) );
  BUFFD0 U2724 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2725 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2726 ( .I(N65), .Z(n2740) );
  BUFFD0 U2727 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2728 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2729 ( .I(n2744), .Z(n2743) );
  BUFFD0 U2730 ( .I(n2745), .Z(n2744) );
  BUFFD0 U2731 ( .I(n2746), .Z(n2745) );
  BUFFD0 U2732 ( .I(n2747), .Z(n2746) );
  BUFFD0 U2733 ( .I(n2748), .Z(n2747) );
  BUFFD0 U2734 ( .I(n2749), .Z(n2748) );
  BUFFD0 U2735 ( .I(n2750), .Z(n2749) );
  BUFFD0 U2736 ( .I(n2751), .Z(n2750) );
  BUFFD0 U2737 ( .I(n2752), .Z(n2751) );
  BUFFD0 U2738 ( .I(n2753), .Z(n2752) );
  BUFFD0 U2739 ( .I(n2754), .Z(n2753) );
  BUFFD0 U2740 ( .I(n2755), .Z(n2754) );
  BUFFD0 U2741 ( .I(n2756), .Z(n2755) );
  BUFFD0 U2742 ( .I(n2757), .Z(n2756) );
  BUFFD0 U2743 ( .I(n2758), .Z(n2757) );
  BUFFD0 U2744 ( .I(n2759), .Z(n2758) );
  BUFFD0 U2745 ( .I(n2760), .Z(n2759) );
  BUFFD0 U2746 ( .I(n2761), .Z(n2760) );
  BUFFD0 U2747 ( .I(n2762), .Z(n2761) );
  BUFFD0 U2748 ( .I(n2763), .Z(n2762) );
  BUFFD0 U2749 ( .I(n2764), .Z(n2763) );
  BUFFD0 U2750 ( .I(n2765), .Z(n2764) );
  BUFFD0 U2751 ( .I(n2766), .Z(n2765) );
  BUFFD0 U2752 ( .I(n2767), .Z(n2766) );
  BUFFD0 U2753 ( .I(n2768), .Z(n2767) );
  BUFFD0 U2754 ( .I(n2769), .Z(n2768) );
  BUFFD0 U2755 ( .I(n2770), .Z(n2769) );
  BUFFD0 U2756 ( .I(n2771), .Z(n2770) );
  BUFFD0 U2757 ( .I(n2772), .Z(n2771) );
  BUFFD0 U2758 ( .I(n2773), .Z(n2772) );
  BUFFD0 U2759 ( .I(n2774), .Z(n2773) );
  BUFFD0 U2760 ( .I(n2775), .Z(n2774) );
  BUFFD0 U2761 ( .I(n2776), .Z(n2775) );
  BUFFD0 U2762 ( .I(n2777), .Z(n2776) );
  BUFFD0 U2763 ( .I(n2778), .Z(n2777) );
  BUFFD0 U2764 ( .I(n2779), .Z(n2778) );
  BUFFD0 U2765 ( .I(n2780), .Z(n2779) );
  BUFFD0 U2766 ( .I(n2781), .Z(n2780) );
  BUFFD0 U2767 ( .I(n2782), .Z(n2781) );
  BUFFD0 U2768 ( .I(n2783), .Z(n2782) );
  BUFFD0 U2769 ( .I(n2784), .Z(n2783) );
  BUFFD0 U2770 ( .I(n2785), .Z(n2784) );
  BUFFD0 U2771 ( .I(n2786), .Z(n2785) );
  BUFFD0 U2772 ( .I(n2787), .Z(n2786) );
  BUFFD0 U2773 ( .I(n2788), .Z(n2787) );
  BUFFD0 U2774 ( .I(n2789), .Z(n2788) );
  BUFFD0 U2775 ( .I(n2790), .Z(n2789) );
  BUFFD0 U2776 ( .I(n2791), .Z(n2790) );
  BUFFD0 U2777 ( .I(n2792), .Z(n2791) );
  BUFFD0 U2778 ( .I(n2793), .Z(n2792) );
  BUFFD0 U2779 ( .I(n2794), .Z(n2793) );
  BUFFD0 U2780 ( .I(n2795), .Z(n2794) );
  BUFFD0 U2781 ( .I(n2796), .Z(n2795) );
  BUFFD0 U2782 ( .I(n2797), .Z(n2796) );
  BUFFD0 U2783 ( .I(n2798), .Z(n2797) );
  BUFFD0 U2784 ( .I(n2799), .Z(n2798) );
  BUFFD0 U2785 ( .I(n2800), .Z(n2799) );
  BUFFD0 U2786 ( .I(n2801), .Z(n2800) );
  BUFFD0 U2787 ( .I(n2802), .Z(n2801) );
  BUFFD0 U2788 ( .I(n2803), .Z(n2802) );
  BUFFD0 U2789 ( .I(n2804), .Z(n2803) );
  BUFFD0 U2790 ( .I(n2805), .Z(n2804) );
  BUFFD0 U2791 ( .I(n2806), .Z(n2805) );
  BUFFD0 U2792 ( .I(n2807), .Z(n2806) );
  BUFFD0 U2793 ( .I(n2808), .Z(n2807) );
  BUFFD0 U2794 ( .I(n2809), .Z(n2808) );
  BUFFD0 U2795 ( .I(n2810), .Z(n2809) );
  BUFFD0 U2796 ( .I(N66), .Z(n2810) );
  BUFFD0 U2797 ( .I(n2812), .Z(n2811) );
  BUFFD0 U2798 ( .I(n2813), .Z(n2812) );
  BUFFD0 U2799 ( .I(n2814), .Z(n2813) );
  BUFFD0 U2800 ( .I(n2815), .Z(n2814) );
  BUFFD0 U2801 ( .I(n2816), .Z(n2815) );
  BUFFD0 U2802 ( .I(n2817), .Z(n2816) );
  BUFFD0 U2803 ( .I(n2818), .Z(n2817) );
  BUFFD0 U2804 ( .I(n2819), .Z(n2818) );
  BUFFD0 U2805 ( .I(n2820), .Z(n2819) );
  BUFFD0 U2806 ( .I(n2821), .Z(n2820) );
  BUFFD0 U2807 ( .I(n2822), .Z(n2821) );
  BUFFD0 U2808 ( .I(n2823), .Z(n2822) );
  BUFFD0 U2809 ( .I(n2824), .Z(n2823) );
  BUFFD0 U2810 ( .I(n2825), .Z(n2824) );
  BUFFD0 U2811 ( .I(n2826), .Z(n2825) );
  BUFFD0 U2812 ( .I(n2827), .Z(n2826) );
  BUFFD0 U2813 ( .I(n2828), .Z(n2827) );
  BUFFD0 U2814 ( .I(n2829), .Z(n2828) );
  BUFFD0 U2815 ( .I(n2830), .Z(n2829) );
  BUFFD0 U2816 ( .I(n2831), .Z(n2830) );
  BUFFD0 U2817 ( .I(n2832), .Z(n2831) );
  BUFFD0 U2818 ( .I(n2833), .Z(n2832) );
  BUFFD0 U2819 ( .I(n2834), .Z(n2833) );
  BUFFD0 U2820 ( .I(n2835), .Z(n2834) );
  BUFFD0 U2821 ( .I(n2836), .Z(n2835) );
  BUFFD0 U2822 ( .I(n2837), .Z(n2836) );
  BUFFD0 U2823 ( .I(n2838), .Z(n2837) );
  BUFFD0 U2824 ( .I(n2839), .Z(n2838) );
  BUFFD0 U2825 ( .I(n2840), .Z(n2839) );
  BUFFD0 U2826 ( .I(n2841), .Z(n2840) );
  BUFFD0 U2827 ( .I(n2842), .Z(n2841) );
  BUFFD0 U2828 ( .I(n2843), .Z(n2842) );
  BUFFD0 U2829 ( .I(n2844), .Z(n2843) );
  BUFFD0 U2830 ( .I(n2845), .Z(n2844) );
  BUFFD0 U2831 ( .I(n2846), .Z(n2845) );
  BUFFD0 U2832 ( .I(n2847), .Z(n2846) );
  BUFFD0 U2833 ( .I(n2848), .Z(n2847) );
  BUFFD0 U2834 ( .I(n2849), .Z(n2848) );
  BUFFD0 U2835 ( .I(n2850), .Z(n2849) );
  BUFFD0 U2836 ( .I(n2851), .Z(n2850) );
  BUFFD0 U2837 ( .I(n2852), .Z(n2851) );
  BUFFD0 U2838 ( .I(n2853), .Z(n2852) );
  BUFFD0 U2839 ( .I(n2854), .Z(n2853) );
  BUFFD0 U2840 ( .I(n2855), .Z(n2854) );
  BUFFD0 U2841 ( .I(n2856), .Z(n2855) );
  BUFFD0 U2842 ( .I(n2857), .Z(n2856) );
  BUFFD0 U2843 ( .I(n2858), .Z(n2857) );
  BUFFD0 U2844 ( .I(n2859), .Z(n2858) );
  BUFFD0 U2845 ( .I(n2860), .Z(n2859) );
  BUFFD0 U2846 ( .I(n2861), .Z(n2860) );
  BUFFD0 U2847 ( .I(n2862), .Z(n2861) );
  BUFFD0 U2848 ( .I(n2863), .Z(n2862) );
  BUFFD0 U2849 ( .I(n2864), .Z(n2863) );
  BUFFD0 U2850 ( .I(n2865), .Z(n2864) );
  BUFFD0 U2851 ( .I(n2866), .Z(n2865) );
  BUFFD0 U2852 ( .I(n2867), .Z(n2866) );
  BUFFD0 U2853 ( .I(n2868), .Z(n2867) );
  BUFFD0 U2854 ( .I(n2869), .Z(n2868) );
  BUFFD0 U2855 ( .I(n2870), .Z(n2869) );
  BUFFD0 U2856 ( .I(n2871), .Z(n2870) );
  BUFFD0 U2857 ( .I(n2872), .Z(n2871) );
  BUFFD0 U2858 ( .I(n2873), .Z(n2872) );
  BUFFD0 U2859 ( .I(n2874), .Z(n2873) );
  BUFFD0 U2860 ( .I(n2875), .Z(n2874) );
  BUFFD0 U2861 ( .I(n2876), .Z(n2875) );
  BUFFD0 U2862 ( .I(n2877), .Z(n2876) );
  BUFFD0 U2863 ( .I(n2878), .Z(n2877) );
  BUFFD0 U2864 ( .I(n2879), .Z(n2878) );
  BUFFD0 U2865 ( .I(n2880), .Z(n2879) );
  BUFFD0 U2866 ( .I(N67), .Z(n2880) );
  BUFFD0 U2867 ( .I(n2882), .Z(n2881) );
  BUFFD0 U2868 ( .I(n2883), .Z(n2882) );
  BUFFD0 U2869 ( .I(n2884), .Z(n2883) );
  BUFFD0 U2870 ( .I(n2885), .Z(n2884) );
  BUFFD0 U2871 ( .I(n2886), .Z(n2885) );
  BUFFD0 U2872 ( .I(n2887), .Z(n2886) );
  BUFFD0 U2873 ( .I(n2888), .Z(n2887) );
  BUFFD0 U2874 ( .I(n2889), .Z(n2888) );
  BUFFD0 U2875 ( .I(n2890), .Z(n2889) );
  BUFFD0 U2876 ( .I(n2891), .Z(n2890) );
  BUFFD0 U2877 ( .I(n2892), .Z(n2891) );
  BUFFD0 U2878 ( .I(n2893), .Z(n2892) );
  BUFFD0 U2879 ( .I(n2894), .Z(n2893) );
  BUFFD0 U2880 ( .I(n2895), .Z(n2894) );
  BUFFD0 U2881 ( .I(n2896), .Z(n2895) );
  BUFFD0 U2882 ( .I(n2897), .Z(n2896) );
  BUFFD0 U2883 ( .I(n2898), .Z(n2897) );
  BUFFD0 U2884 ( .I(n2899), .Z(n2898) );
  BUFFD0 U2885 ( .I(n2900), .Z(n2899) );
  BUFFD0 U2886 ( .I(n2901), .Z(n2900) );
  BUFFD0 U2887 ( .I(n2902), .Z(n2901) );
  BUFFD0 U2888 ( .I(n2903), .Z(n2902) );
  BUFFD0 U2889 ( .I(n2904), .Z(n2903) );
  BUFFD0 U2890 ( .I(n2905), .Z(n2904) );
  BUFFD0 U2891 ( .I(n2906), .Z(n2905) );
  BUFFD0 U2892 ( .I(n2907), .Z(n2906) );
  BUFFD0 U2893 ( .I(n2908), .Z(n2907) );
  BUFFD0 U2894 ( .I(n2909), .Z(n2908) );
  BUFFD0 U2895 ( .I(n2910), .Z(n2909) );
  BUFFD0 U2896 ( .I(n2911), .Z(n2910) );
  BUFFD0 U2897 ( .I(n2912), .Z(n2911) );
  BUFFD0 U2898 ( .I(n2913), .Z(n2912) );
  BUFFD0 U2899 ( .I(n2914), .Z(n2913) );
  BUFFD0 U2900 ( .I(n2915), .Z(n2914) );
  BUFFD0 U2901 ( .I(n2916), .Z(n2915) );
  BUFFD0 U2902 ( .I(n2917), .Z(n2916) );
  BUFFD0 U2903 ( .I(n2918), .Z(n2917) );
  BUFFD0 U2904 ( .I(n2919), .Z(n2918) );
  BUFFD0 U2905 ( .I(n2920), .Z(n2919) );
  BUFFD0 U2906 ( .I(n2921), .Z(n2920) );
  BUFFD0 U2907 ( .I(n2922), .Z(n2921) );
  BUFFD0 U2908 ( .I(n2923), .Z(n2922) );
  BUFFD0 U2909 ( .I(n2924), .Z(n2923) );
  BUFFD0 U2910 ( .I(n2925), .Z(n2924) );
  BUFFD0 U2911 ( .I(n2926), .Z(n2925) );
  BUFFD0 U2912 ( .I(n2927), .Z(n2926) );
  BUFFD0 U2913 ( .I(n2928), .Z(n2927) );
  BUFFD0 U2914 ( .I(n2929), .Z(n2928) );
  BUFFD0 U2915 ( .I(n2930), .Z(n2929) );
  BUFFD0 U2916 ( .I(n2931), .Z(n2930) );
  BUFFD0 U2917 ( .I(n2932), .Z(n2931) );
  BUFFD0 U2918 ( .I(n2933), .Z(n2932) );
  BUFFD0 U2919 ( .I(n2934), .Z(n2933) );
  BUFFD0 U2920 ( .I(n2935), .Z(n2934) );
  BUFFD0 U2921 ( .I(n2936), .Z(n2935) );
  BUFFD0 U2922 ( .I(n2937), .Z(n2936) );
  BUFFD0 U2923 ( .I(n2938), .Z(n2937) );
  BUFFD0 U2924 ( .I(n2939), .Z(n2938) );
  BUFFD0 U2925 ( .I(n2940), .Z(n2939) );
  BUFFD0 U2926 ( .I(n2941), .Z(n2940) );
  BUFFD0 U2927 ( .I(n2942), .Z(n2941) );
  BUFFD0 U2928 ( .I(n2943), .Z(n2942) );
  BUFFD0 U2929 ( .I(n2944), .Z(n2943) );
  BUFFD0 U2930 ( .I(n2945), .Z(n2944) );
  BUFFD0 U2931 ( .I(n2946), .Z(n2945) );
  BUFFD0 U2932 ( .I(n2947), .Z(n2946) );
  BUFFD0 U2933 ( .I(n2948), .Z(n2947) );
  BUFFD0 U2934 ( .I(n2949), .Z(n2948) );
  BUFFD0 U2935 ( .I(n2950), .Z(n2949) );
  BUFFD0 U2936 ( .I(N68), .Z(n2950) );
  BUFFD0 U2937 ( .I(n2952), .Z(n2951) );
  BUFFD0 U2938 ( .I(n2953), .Z(n2952) );
  BUFFD0 U2939 ( .I(n2954), .Z(n2953) );
  BUFFD0 U2940 ( .I(n2955), .Z(n2954) );
  BUFFD0 U2941 ( .I(n2956), .Z(n2955) );
  BUFFD0 U2942 ( .I(n2957), .Z(n2956) );
  BUFFD0 U2943 ( .I(n2958), .Z(n2957) );
  BUFFD0 U2944 ( .I(n2959), .Z(n2958) );
  BUFFD0 U2945 ( .I(n2960), .Z(n2959) );
  BUFFD0 U2946 ( .I(n2961), .Z(n2960) );
  BUFFD0 U2947 ( .I(n2962), .Z(n2961) );
  BUFFD0 U2948 ( .I(n2963), .Z(n2962) );
  BUFFD0 U2949 ( .I(n2964), .Z(n2963) );
  BUFFD0 U2950 ( .I(n2965), .Z(n2964) );
  BUFFD0 U2951 ( .I(n2966), .Z(n2965) );
  BUFFD0 U2952 ( .I(n2967), .Z(n2966) );
  BUFFD0 U2953 ( .I(n2968), .Z(n2967) );
  BUFFD0 U2954 ( .I(n2969), .Z(n2968) );
  BUFFD0 U2955 ( .I(n2970), .Z(n2969) );
  BUFFD0 U2956 ( .I(n2971), .Z(n2970) );
  BUFFD0 U2957 ( .I(n2972), .Z(n2971) );
  BUFFD0 U2958 ( .I(n2973), .Z(n2972) );
  BUFFD0 U2959 ( .I(n2974), .Z(n2973) );
  BUFFD0 U2960 ( .I(n2975), .Z(n2974) );
  BUFFD0 U2961 ( .I(n2976), .Z(n2975) );
  BUFFD0 U2962 ( .I(n2977), .Z(n2976) );
  BUFFD0 U2963 ( .I(n2978), .Z(n2977) );
  BUFFD0 U2964 ( .I(n2979), .Z(n2978) );
  BUFFD0 U2965 ( .I(n2980), .Z(n2979) );
  BUFFD0 U2966 ( .I(n2981), .Z(n2980) );
  BUFFD0 U2967 ( .I(n2982), .Z(n2981) );
  BUFFD0 U2968 ( .I(n2983), .Z(n2982) );
  BUFFD0 U2969 ( .I(n2984), .Z(n2983) );
  BUFFD0 U2970 ( .I(n2985), .Z(n2984) );
  BUFFD0 U2971 ( .I(n2986), .Z(n2985) );
  BUFFD0 U2972 ( .I(n2987), .Z(n2986) );
  BUFFD0 U2973 ( .I(n2988), .Z(n2987) );
  BUFFD0 U2974 ( .I(n2989), .Z(n2988) );
  BUFFD0 U2975 ( .I(n2990), .Z(n2989) );
  BUFFD0 U2976 ( .I(n2991), .Z(n2990) );
  BUFFD0 U2977 ( .I(n2992), .Z(n2991) );
  BUFFD0 U2978 ( .I(n2993), .Z(n2992) );
  BUFFD0 U2979 ( .I(n2994), .Z(n2993) );
  BUFFD0 U2980 ( .I(n2995), .Z(n2994) );
  BUFFD0 U2981 ( .I(n2996), .Z(n2995) );
  BUFFD0 U2982 ( .I(n2997), .Z(n2996) );
  BUFFD0 U2983 ( .I(n2998), .Z(n2997) );
  BUFFD0 U2984 ( .I(n2999), .Z(n2998) );
  BUFFD0 U2985 ( .I(n3000), .Z(n2999) );
  BUFFD0 U2986 ( .I(n3001), .Z(n3000) );
  BUFFD0 U2987 ( .I(n3002), .Z(n3001) );
  BUFFD0 U2988 ( .I(n3003), .Z(n3002) );
  BUFFD0 U2989 ( .I(n3004), .Z(n3003) );
  BUFFD0 U2990 ( .I(n3005), .Z(n3004) );
  BUFFD0 U2991 ( .I(n3006), .Z(n3005) );
  BUFFD0 U2992 ( .I(n3007), .Z(n3006) );
  BUFFD0 U2993 ( .I(n3008), .Z(n3007) );
  BUFFD0 U2994 ( .I(n3009), .Z(n3008) );
  BUFFD0 U2995 ( .I(n3010), .Z(n3009) );
  BUFFD0 U2996 ( .I(n3011), .Z(n3010) );
  BUFFD0 U2997 ( .I(n3012), .Z(n3011) );
  BUFFD0 U2998 ( .I(n3013), .Z(n3012) );
  BUFFD0 U2999 ( .I(n3014), .Z(n3013) );
  BUFFD0 U3000 ( .I(n3015), .Z(n3014) );
  BUFFD0 U3001 ( .I(n3016), .Z(n3015) );
  BUFFD0 U3002 ( .I(n3017), .Z(n3016) );
  BUFFD0 U3003 ( .I(n3018), .Z(n3017) );
  BUFFD0 U3004 ( .I(n3019), .Z(n3018) );
  BUFFD0 U3005 ( .I(n3020), .Z(n3019) );
  BUFFD0 U3006 ( .I(N69), .Z(n3020) );
  BUFFD0 U3007 ( .I(n3022), .Z(n3021) );
  BUFFD0 U3008 ( .I(n3023), .Z(n3022) );
  BUFFD0 U3009 ( .I(n3024), .Z(n3023) );
  BUFFD0 U3010 ( .I(n3025), .Z(n3024) );
  BUFFD0 U3011 ( .I(n3026), .Z(n3025) );
  BUFFD0 U3012 ( .I(n3027), .Z(n3026) );
  BUFFD0 U3013 ( .I(n3028), .Z(n3027) );
  BUFFD0 U3014 ( .I(n3029), .Z(n3028) );
  BUFFD0 U3015 ( .I(n3030), .Z(n3029) );
  BUFFD0 U3016 ( .I(n3031), .Z(n3030) );
  BUFFD0 U3017 ( .I(n3032), .Z(n3031) );
  BUFFD0 U3018 ( .I(n3033), .Z(n3032) );
  BUFFD0 U3019 ( .I(n3034), .Z(n3033) );
  BUFFD0 U3020 ( .I(n3035), .Z(n3034) );
  BUFFD0 U3021 ( .I(n3036), .Z(n3035) );
  BUFFD0 U3022 ( .I(n3037), .Z(n3036) );
  BUFFD0 U3023 ( .I(n3038), .Z(n3037) );
  BUFFD0 U3024 ( .I(n3039), .Z(n3038) );
  BUFFD0 U3025 ( .I(n3040), .Z(n3039) );
  BUFFD0 U3026 ( .I(n3041), .Z(n3040) );
  BUFFD0 U3027 ( .I(n3042), .Z(n3041) );
  BUFFD0 U3028 ( .I(n3043), .Z(n3042) );
  BUFFD0 U3029 ( .I(n3044), .Z(n3043) );
  BUFFD0 U3030 ( .I(n3045), .Z(n3044) );
  BUFFD0 U3031 ( .I(n3046), .Z(n3045) );
  BUFFD0 U3032 ( .I(n3047), .Z(n3046) );
  BUFFD0 U3033 ( .I(n3048), .Z(n3047) );
  BUFFD0 U3034 ( .I(n3049), .Z(n3048) );
  BUFFD0 U3035 ( .I(n3050), .Z(n3049) );
  BUFFD0 U3036 ( .I(n3051), .Z(n3050) );
  BUFFD0 U3037 ( .I(n3052), .Z(n3051) );
  BUFFD0 U3038 ( .I(n3053), .Z(n3052) );
  BUFFD0 U3039 ( .I(n3054), .Z(n3053) );
  BUFFD0 U3040 ( .I(n3055), .Z(n3054) );
  BUFFD0 U3041 ( .I(n3056), .Z(n3055) );
  BUFFD0 U3042 ( .I(n3057), .Z(n3056) );
  BUFFD0 U3043 ( .I(n3058), .Z(n3057) );
  BUFFD0 U3044 ( .I(n3059), .Z(n3058) );
  BUFFD0 U3045 ( .I(n3060), .Z(n3059) );
  BUFFD0 U3046 ( .I(n3061), .Z(n3060) );
  BUFFD0 U3047 ( .I(n3062), .Z(n3061) );
  BUFFD0 U3048 ( .I(n3063), .Z(n3062) );
  BUFFD0 U3049 ( .I(n3064), .Z(n3063) );
  BUFFD0 U3050 ( .I(n3065), .Z(n3064) );
  BUFFD0 U3051 ( .I(n3066), .Z(n3065) );
  BUFFD0 U3052 ( .I(n3067), .Z(n3066) );
  BUFFD0 U3053 ( .I(n3068), .Z(n3067) );
  BUFFD0 U3054 ( .I(n3069), .Z(n3068) );
  BUFFD0 U3055 ( .I(n3070), .Z(n3069) );
  BUFFD0 U3056 ( .I(n3071), .Z(n3070) );
  BUFFD0 U3057 ( .I(n3072), .Z(n3071) );
  BUFFD0 U3058 ( .I(n3073), .Z(n3072) );
  BUFFD0 U3059 ( .I(n3074), .Z(n3073) );
  BUFFD0 U3060 ( .I(n3075), .Z(n3074) );
  BUFFD0 U3061 ( .I(n3076), .Z(n3075) );
  BUFFD0 U3062 ( .I(n3077), .Z(n3076) );
  BUFFD0 U3063 ( .I(n3078), .Z(n3077) );
  BUFFD0 U3064 ( .I(n3079), .Z(n3078) );
  BUFFD0 U3065 ( .I(n3080), .Z(n3079) );
  BUFFD0 U3066 ( .I(n3081), .Z(n3080) );
  BUFFD0 U3067 ( .I(n3082), .Z(n3081) );
  BUFFD0 U3068 ( .I(n3083), .Z(n3082) );
  BUFFD0 U3069 ( .I(n3084), .Z(n3083) );
  BUFFD0 U3070 ( .I(n3085), .Z(n3084) );
  BUFFD0 U3071 ( .I(n3086), .Z(n3085) );
  BUFFD0 U3072 ( .I(n3087), .Z(n3086) );
  BUFFD0 U3073 ( .I(n3088), .Z(n3087) );
  BUFFD0 U3074 ( .I(n3089), .Z(n3088) );
  BUFFD0 U3075 ( .I(n3090), .Z(n3089) );
  BUFFD0 U3076 ( .I(N70), .Z(n3090) );
  BUFFD0 U3077 ( .I(n3092), .Z(n3091) );
  BUFFD0 U3078 ( .I(n3093), .Z(n3092) );
  BUFFD0 U3079 ( .I(n3094), .Z(n3093) );
  BUFFD0 U3080 ( .I(n3095), .Z(n3094) );
  BUFFD0 U3081 ( .I(n3096), .Z(n3095) );
  BUFFD0 U3082 ( .I(n3097), .Z(n3096) );
  BUFFD0 U3083 ( .I(n3098), .Z(n3097) );
  BUFFD0 U3084 ( .I(n3099), .Z(n3098) );
  BUFFD0 U3085 ( .I(n3100), .Z(n3099) );
  BUFFD0 U3086 ( .I(n3101), .Z(n3100) );
  BUFFD0 U3087 ( .I(n3102), .Z(n3101) );
  BUFFD0 U3088 ( .I(n3103), .Z(n3102) );
  BUFFD0 U3089 ( .I(n3104), .Z(n3103) );
  BUFFD0 U3090 ( .I(n3105), .Z(n3104) );
  BUFFD0 U3091 ( .I(n3106), .Z(n3105) );
  BUFFD0 U3092 ( .I(n3107), .Z(n3106) );
  BUFFD0 U3093 ( .I(n3108), .Z(n3107) );
  BUFFD0 U3094 ( .I(n3109), .Z(n3108) );
  BUFFD0 U3095 ( .I(n3110), .Z(n3109) );
  BUFFD0 U3096 ( .I(n3111), .Z(n3110) );
  BUFFD0 U3097 ( .I(n3112), .Z(n3111) );
  BUFFD0 U3098 ( .I(n3113), .Z(n3112) );
  BUFFD0 U3099 ( .I(n3114), .Z(n3113) );
  BUFFD0 U3100 ( .I(n3115), .Z(n3114) );
  BUFFD0 U3101 ( .I(n3116), .Z(n3115) );
  BUFFD0 U3102 ( .I(n3117), .Z(n3116) );
  BUFFD0 U3103 ( .I(n3118), .Z(n3117) );
  BUFFD0 U3104 ( .I(n3119), .Z(n3118) );
  BUFFD0 U3105 ( .I(n3120), .Z(n3119) );
  BUFFD0 U3106 ( .I(n3121), .Z(n3120) );
  BUFFD0 U3107 ( .I(n3122), .Z(n3121) );
  BUFFD0 U3108 ( .I(n3123), .Z(n3122) );
  BUFFD0 U3109 ( .I(n3124), .Z(n3123) );
  BUFFD0 U3110 ( .I(n3125), .Z(n3124) );
  BUFFD0 U3111 ( .I(n3126), .Z(n3125) );
  BUFFD0 U3112 ( .I(n3127), .Z(n3126) );
  BUFFD0 U3113 ( .I(n3128), .Z(n3127) );
  BUFFD0 U3114 ( .I(n3129), .Z(n3128) );
  BUFFD0 U3115 ( .I(n3130), .Z(n3129) );
  BUFFD0 U3116 ( .I(n3131), .Z(n3130) );
  BUFFD0 U3117 ( .I(n3132), .Z(n3131) );
  BUFFD0 U3118 ( .I(n3133), .Z(n3132) );
  BUFFD0 U3119 ( .I(n3134), .Z(n3133) );
  BUFFD0 U3120 ( .I(n3135), .Z(n3134) );
  BUFFD0 U3121 ( .I(n3136), .Z(n3135) );
  BUFFD0 U3122 ( .I(n3137), .Z(n3136) );
  BUFFD0 U3123 ( .I(n3138), .Z(n3137) );
  BUFFD0 U3124 ( .I(n3139), .Z(n3138) );
  BUFFD0 U3125 ( .I(n3140), .Z(n3139) );
  BUFFD0 U3126 ( .I(n3141), .Z(n3140) );
  BUFFD0 U3127 ( .I(n3142), .Z(n3141) );
  BUFFD0 U3128 ( .I(n3143), .Z(n3142) );
  BUFFD0 U3129 ( .I(n3144), .Z(n3143) );
  BUFFD0 U3130 ( .I(n3145), .Z(n3144) );
  BUFFD0 U3131 ( .I(n3146), .Z(n3145) );
  BUFFD0 U3132 ( .I(n3147), .Z(n3146) );
  BUFFD0 U3133 ( .I(n3148), .Z(n3147) );
  BUFFD0 U3134 ( .I(n3149), .Z(n3148) );
  BUFFD0 U3135 ( .I(n3150), .Z(n3149) );
  BUFFD0 U3136 ( .I(n3151), .Z(n3150) );
  BUFFD0 U3137 ( .I(n3152), .Z(n3151) );
  BUFFD0 U3138 ( .I(n3153), .Z(n3152) );
  BUFFD0 U3139 ( .I(n3154), .Z(n3153) );
  BUFFD0 U3140 ( .I(n3155), .Z(n3154) );
  BUFFD0 U3141 ( .I(n3156), .Z(n3155) );
  BUFFD0 U3142 ( .I(n3157), .Z(n3156) );
  BUFFD0 U3143 ( .I(n3158), .Z(n3157) );
  BUFFD0 U3144 ( .I(n3159), .Z(n3158) );
  BUFFD0 U3145 ( .I(n3160), .Z(n3159) );
  BUFFD0 U3146 ( .I(N71), .Z(n3160) );
  BUFFD0 U3147 ( .I(n3162), .Z(n3161) );
  BUFFD0 U3148 ( .I(n3163), .Z(n3162) );
  BUFFD0 U3149 ( .I(n3164), .Z(n3163) );
  BUFFD0 U3150 ( .I(n3165), .Z(n3164) );
  BUFFD0 U3151 ( .I(n3166), .Z(n3165) );
  BUFFD0 U3152 ( .I(n3167), .Z(n3166) );
  BUFFD0 U3153 ( .I(n3168), .Z(n3167) );
  BUFFD0 U3154 ( .I(n3169), .Z(n3168) );
  BUFFD0 U3155 ( .I(n3170), .Z(n3169) );
  BUFFD0 U3156 ( .I(n3171), .Z(n3170) );
  BUFFD0 U3157 ( .I(n3172), .Z(n3171) );
  BUFFD0 U3158 ( .I(n3173), .Z(n3172) );
  BUFFD0 U3159 ( .I(n3174), .Z(n3173) );
  BUFFD0 U3160 ( .I(n3175), .Z(n3174) );
  BUFFD0 U3161 ( .I(n3176), .Z(n3175) );
  BUFFD0 U3162 ( .I(n3177), .Z(n3176) );
  BUFFD0 U3163 ( .I(n3178), .Z(n3177) );
  BUFFD0 U3164 ( .I(n3179), .Z(n3178) );
  BUFFD0 U3165 ( .I(n3180), .Z(n3179) );
  BUFFD0 U3166 ( .I(n3181), .Z(n3180) );
  BUFFD0 U3167 ( .I(n3182), .Z(n3181) );
  BUFFD0 U3168 ( .I(n3183), .Z(n3182) );
  BUFFD0 U3169 ( .I(n3184), .Z(n3183) );
  BUFFD0 U3170 ( .I(n3185), .Z(n3184) );
  BUFFD0 U3171 ( .I(n3186), .Z(n3185) );
  BUFFD0 U3172 ( .I(n3187), .Z(n3186) );
  BUFFD0 U3173 ( .I(n3188), .Z(n3187) );
  BUFFD0 U3174 ( .I(n3189), .Z(n3188) );
  BUFFD0 U3175 ( .I(n3190), .Z(n3189) );
  BUFFD0 U3176 ( .I(n3191), .Z(n3190) );
  BUFFD0 U3177 ( .I(n3192), .Z(n3191) );
  BUFFD0 U3178 ( .I(n3193), .Z(n3192) );
  BUFFD0 U3179 ( .I(n3194), .Z(n3193) );
  BUFFD0 U3180 ( .I(n3195), .Z(n3194) );
  BUFFD0 U3181 ( .I(n3196), .Z(n3195) );
  BUFFD0 U3182 ( .I(n3197), .Z(n3196) );
  BUFFD0 U3183 ( .I(n3198), .Z(n3197) );
  BUFFD0 U3184 ( .I(n3199), .Z(n3198) );
  BUFFD0 U3185 ( .I(n3200), .Z(n3199) );
  BUFFD0 U3186 ( .I(n3201), .Z(n3200) );
  BUFFD0 U3187 ( .I(n3202), .Z(n3201) );
  BUFFD0 U3188 ( .I(n3203), .Z(n3202) );
  BUFFD0 U3189 ( .I(n3204), .Z(n3203) );
  BUFFD0 U3190 ( .I(n3205), .Z(n3204) );
  BUFFD0 U3191 ( .I(n3206), .Z(n3205) );
  BUFFD0 U3192 ( .I(n3207), .Z(n3206) );
  BUFFD0 U3193 ( .I(n3208), .Z(n3207) );
  BUFFD0 U3194 ( .I(n3209), .Z(n3208) );
  BUFFD0 U3195 ( .I(n3210), .Z(n3209) );
  BUFFD0 U3196 ( .I(n3211), .Z(n3210) );
  BUFFD0 U3197 ( .I(n3212), .Z(n3211) );
  BUFFD0 U3198 ( .I(n3213), .Z(n3212) );
  BUFFD0 U3199 ( .I(n3214), .Z(n3213) );
  BUFFD0 U3200 ( .I(n3215), .Z(n3214) );
  BUFFD0 U3201 ( .I(n3216), .Z(n3215) );
  BUFFD0 U3202 ( .I(n3217), .Z(n3216) );
  BUFFD0 U3203 ( .I(n3218), .Z(n3217) );
  BUFFD0 U3204 ( .I(n3219), .Z(n3218) );
  BUFFD0 U3205 ( .I(n3220), .Z(n3219) );
  BUFFD0 U3206 ( .I(n3221), .Z(n3220) );
  BUFFD0 U3207 ( .I(n3222), .Z(n3221) );
  BUFFD0 U3208 ( .I(n3223), .Z(n3222) );
  BUFFD0 U3209 ( .I(n3224), .Z(n3223) );
  BUFFD0 U3210 ( .I(n3225), .Z(n3224) );
  BUFFD0 U3211 ( .I(n3226), .Z(n3225) );
  BUFFD0 U3212 ( .I(n3227), .Z(n3226) );
  BUFFD0 U3213 ( .I(n3228), .Z(n3227) );
  BUFFD0 U3214 ( .I(n3229), .Z(n3228) );
  BUFFD0 U3215 ( .I(n3230), .Z(n3229) );
  BUFFD0 U3216 ( .I(N72), .Z(n3230) );
  BUFFD0 U3217 ( .I(n3232), .Z(n3231) );
  BUFFD0 U3218 ( .I(n3233), .Z(n3232) );
  BUFFD0 U3219 ( .I(n3234), .Z(n3233) );
  BUFFD0 U3220 ( .I(n3235), .Z(n3234) );
  BUFFD0 U3221 ( .I(n3236), .Z(n3235) );
  BUFFD0 U3222 ( .I(n3237), .Z(n3236) );
  BUFFD0 U3223 ( .I(n3238), .Z(n3237) );
  BUFFD0 U3224 ( .I(n3239), .Z(n3238) );
  BUFFD0 U3225 ( .I(n3240), .Z(n3239) );
  BUFFD0 U3226 ( .I(n3241), .Z(n3240) );
  BUFFD0 U3227 ( .I(n3242), .Z(n3241) );
  BUFFD0 U3228 ( .I(n3243), .Z(n3242) );
  BUFFD0 U3229 ( .I(n3244), .Z(n3243) );
  BUFFD0 U3230 ( .I(n3245), .Z(n3244) );
  BUFFD0 U3231 ( .I(n3246), .Z(n3245) );
  BUFFD0 U3232 ( .I(n3247), .Z(n3246) );
  BUFFD0 U3233 ( .I(n3248), .Z(n3247) );
  BUFFD0 U3234 ( .I(n3249), .Z(n3248) );
  BUFFD0 U3235 ( .I(n3250), .Z(n3249) );
  BUFFD0 U3236 ( .I(n3251), .Z(n3250) );
  BUFFD0 U3237 ( .I(n3252), .Z(n3251) );
  BUFFD0 U3238 ( .I(n3253), .Z(n3252) );
  BUFFD0 U3239 ( .I(n3254), .Z(n3253) );
  BUFFD0 U3240 ( .I(n3255), .Z(n3254) );
  BUFFD0 U3241 ( .I(n3256), .Z(n3255) );
  BUFFD0 U3242 ( .I(n3257), .Z(n3256) );
  BUFFD0 U3243 ( .I(n3258), .Z(n3257) );
  BUFFD0 U3244 ( .I(n3259), .Z(n3258) );
  BUFFD0 U3245 ( .I(n3260), .Z(n3259) );
  BUFFD0 U3246 ( .I(n3261), .Z(n3260) );
  BUFFD0 U3247 ( .I(n3262), .Z(n3261) );
  BUFFD0 U3248 ( .I(n3263), .Z(n3262) );
  BUFFD0 U3249 ( .I(n3264), .Z(n3263) );
  BUFFD0 U3250 ( .I(n3265), .Z(n3264) );
  BUFFD0 U3251 ( .I(n3266), .Z(n3265) );
  BUFFD0 U3252 ( .I(n3267), .Z(n3266) );
  BUFFD0 U3253 ( .I(n3268), .Z(n3267) );
  BUFFD0 U3254 ( .I(n3269), .Z(n3268) );
  BUFFD0 U3255 ( .I(n3270), .Z(n3269) );
  BUFFD0 U3256 ( .I(n3271), .Z(n3270) );
  BUFFD0 U3257 ( .I(n3272), .Z(n3271) );
  BUFFD0 U3258 ( .I(n3273), .Z(n3272) );
  BUFFD0 U3259 ( .I(n3274), .Z(n3273) );
  BUFFD0 U3260 ( .I(n3275), .Z(n3274) );
  BUFFD0 U3261 ( .I(n3276), .Z(n3275) );
  BUFFD0 U3262 ( .I(n3277), .Z(n3276) );
  BUFFD0 U3263 ( .I(n3278), .Z(n3277) );
  BUFFD0 U3264 ( .I(n3279), .Z(n3278) );
  BUFFD0 U3265 ( .I(n3280), .Z(n3279) );
  BUFFD0 U3266 ( .I(n3281), .Z(n3280) );
  BUFFD0 U3267 ( .I(n3282), .Z(n3281) );
  BUFFD0 U3268 ( .I(n3283), .Z(n3282) );
  BUFFD0 U3269 ( .I(n3284), .Z(n3283) );
  BUFFD0 U3270 ( .I(n3285), .Z(n3284) );
  BUFFD0 U3271 ( .I(n3286), .Z(n3285) );
  BUFFD0 U3272 ( .I(n3287), .Z(n3286) );
  BUFFD0 U3273 ( .I(n3288), .Z(n3287) );
  BUFFD0 U3274 ( .I(n3289), .Z(n3288) );
  BUFFD0 U3275 ( .I(n3290), .Z(n3289) );
  BUFFD0 U3276 ( .I(n3291), .Z(n3290) );
  BUFFD0 U3277 ( .I(n3292), .Z(n3291) );
  BUFFD0 U3278 ( .I(n3293), .Z(n3292) );
  BUFFD0 U3279 ( .I(n3294), .Z(n3293) );
  BUFFD0 U3280 ( .I(n3295), .Z(n3294) );
  BUFFD0 U3281 ( .I(n3296), .Z(n3295) );
  BUFFD0 U3282 ( .I(n3297), .Z(n3296) );
  BUFFD0 U3283 ( .I(n3298), .Z(n3297) );
  BUFFD0 U3284 ( .I(n3299), .Z(n3298) );
  BUFFD0 U3285 ( .I(n3300), .Z(n3299) );
  BUFFD0 U3286 ( .I(N73), .Z(n3300) );
  BUFFD0 U3287 ( .I(n3302), .Z(n3301) );
  BUFFD0 U3288 ( .I(n3303), .Z(n3302) );
  BUFFD0 U3289 ( .I(n3304), .Z(n3303) );
  BUFFD0 U3290 ( .I(n3305), .Z(n3304) );
  BUFFD0 U3291 ( .I(n3306), .Z(n3305) );
  BUFFD0 U3292 ( .I(n3307), .Z(n3306) );
  BUFFD0 U3293 ( .I(n3308), .Z(n3307) );
  BUFFD0 U3294 ( .I(n3309), .Z(n3308) );
  BUFFD0 U3295 ( .I(n3310), .Z(n3309) );
  BUFFD0 U3296 ( .I(n3311), .Z(n3310) );
  BUFFD0 U3297 ( .I(n3312), .Z(n3311) );
  BUFFD0 U3298 ( .I(n3313), .Z(n3312) );
  BUFFD0 U3299 ( .I(n3314), .Z(n3313) );
  BUFFD0 U3300 ( .I(n3315), .Z(n3314) );
  BUFFD0 U3301 ( .I(n3316), .Z(n3315) );
  BUFFD0 U3302 ( .I(n3317), .Z(n3316) );
  BUFFD0 U3303 ( .I(n3318), .Z(n3317) );
  BUFFD0 U3304 ( .I(n3319), .Z(n3318) );
  BUFFD0 U3305 ( .I(n3320), .Z(n3319) );
  BUFFD0 U3306 ( .I(n3321), .Z(n3320) );
  BUFFD0 U3307 ( .I(n3322), .Z(n3321) );
  BUFFD0 U3308 ( .I(n3323), .Z(n3322) );
  BUFFD0 U3309 ( .I(n3324), .Z(n3323) );
  BUFFD0 U3310 ( .I(n3325), .Z(n3324) );
  BUFFD0 U3311 ( .I(n3326), .Z(n3325) );
  BUFFD0 U3312 ( .I(n3327), .Z(n3326) );
  BUFFD0 U3313 ( .I(n3328), .Z(n3327) );
  BUFFD0 U3314 ( .I(n3329), .Z(n3328) );
  BUFFD0 U3315 ( .I(n3330), .Z(n3329) );
  BUFFD0 U3316 ( .I(n3331), .Z(n3330) );
  BUFFD0 U3317 ( .I(n3332), .Z(n3331) );
  BUFFD0 U3318 ( .I(n3333), .Z(n3332) );
  BUFFD0 U3319 ( .I(n3334), .Z(n3333) );
  BUFFD0 U3320 ( .I(n3335), .Z(n3334) );
  BUFFD0 U3321 ( .I(n3336), .Z(n3335) );
  BUFFD0 U3322 ( .I(n3337), .Z(n3336) );
  BUFFD0 U3323 ( .I(n3338), .Z(n3337) );
  BUFFD0 U3324 ( .I(n3339), .Z(n3338) );
  BUFFD0 U3325 ( .I(n3340), .Z(n3339) );
  BUFFD0 U3326 ( .I(n3341), .Z(n3340) );
  BUFFD0 U3327 ( .I(n3342), .Z(n3341) );
  BUFFD0 U3328 ( .I(n3343), .Z(n3342) );
  BUFFD0 U3329 ( .I(n3344), .Z(n3343) );
  BUFFD0 U3330 ( .I(n3345), .Z(n3344) );
  BUFFD0 U3331 ( .I(n3346), .Z(n3345) );
  BUFFD0 U3332 ( .I(n3347), .Z(n3346) );
  BUFFD0 U3333 ( .I(n3348), .Z(n3347) );
  BUFFD0 U3334 ( .I(n3349), .Z(n3348) );
  BUFFD0 U3335 ( .I(n3350), .Z(n3349) );
  BUFFD0 U3336 ( .I(n3351), .Z(n3350) );
  BUFFD0 U3337 ( .I(n3352), .Z(n3351) );
  BUFFD0 U3338 ( .I(n3353), .Z(n3352) );
  BUFFD0 U3339 ( .I(n3354), .Z(n3353) );
  BUFFD0 U3340 ( .I(n3355), .Z(n3354) );
  BUFFD0 U3341 ( .I(n3356), .Z(n3355) );
  BUFFD0 U3342 ( .I(n3357), .Z(n3356) );
  BUFFD0 U3343 ( .I(n3358), .Z(n3357) );
  BUFFD0 U3344 ( .I(n3359), .Z(n3358) );
  BUFFD0 U3345 ( .I(n3360), .Z(n3359) );
  BUFFD0 U3346 ( .I(n3361), .Z(n3360) );
  BUFFD0 U3347 ( .I(n3362), .Z(n3361) );
  BUFFD0 U3348 ( .I(n3363), .Z(n3362) );
  BUFFD0 U3349 ( .I(n3364), .Z(n3363) );
  BUFFD0 U3350 ( .I(n3365), .Z(n3364) );
  BUFFD0 U3351 ( .I(n3366), .Z(n3365) );
  BUFFD0 U3352 ( .I(n3367), .Z(n3366) );
  BUFFD0 U3353 ( .I(n3368), .Z(n3367) );
  BUFFD0 U3354 ( .I(n3369), .Z(n3368) );
  BUFFD0 U3355 ( .I(n3370), .Z(n3369) );
  BUFFD0 U3356 ( .I(N74), .Z(n3370) );
  BUFFD0 U3357 ( .I(n3372), .Z(n3371) );
  BUFFD0 U3358 ( .I(n3373), .Z(n3372) );
  BUFFD0 U3359 ( .I(n3374), .Z(n3373) );
  BUFFD0 U3360 ( .I(n3375), .Z(n3374) );
  BUFFD0 U3361 ( .I(n3376), .Z(n3375) );
  BUFFD0 U3362 ( .I(n3377), .Z(n3376) );
  BUFFD0 U3363 ( .I(n3378), .Z(n3377) );
  BUFFD0 U3364 ( .I(n3379), .Z(n3378) );
  BUFFD0 U3365 ( .I(n3380), .Z(n3379) );
  BUFFD0 U3366 ( .I(n3381), .Z(n3380) );
  BUFFD0 U3367 ( .I(n3382), .Z(n3381) );
  BUFFD0 U3368 ( .I(n3383), .Z(n3382) );
  BUFFD0 U3369 ( .I(n3384), .Z(n3383) );
  BUFFD0 U3370 ( .I(n3385), .Z(n3384) );
  BUFFD0 U3371 ( .I(n3386), .Z(n3385) );
  BUFFD0 U3372 ( .I(n3387), .Z(n3386) );
  BUFFD0 U3373 ( .I(n3388), .Z(n3387) );
  BUFFD0 U3374 ( .I(n3389), .Z(n3388) );
  BUFFD0 U3375 ( .I(n3390), .Z(n3389) );
  BUFFD0 U3376 ( .I(n3391), .Z(n3390) );
  BUFFD0 U3377 ( .I(n3392), .Z(n3391) );
  BUFFD0 U3378 ( .I(n3393), .Z(n3392) );
  BUFFD0 U3379 ( .I(n3394), .Z(n3393) );
  BUFFD0 U3380 ( .I(n3395), .Z(n3394) );
  BUFFD0 U3381 ( .I(n3396), .Z(n3395) );
  BUFFD0 U3382 ( .I(n3397), .Z(n3396) );
  BUFFD0 U3383 ( .I(n3398), .Z(n3397) );
  BUFFD0 U3384 ( .I(n3399), .Z(n3398) );
  BUFFD0 U3385 ( .I(n3400), .Z(n3399) );
  BUFFD0 U3386 ( .I(n3401), .Z(n3400) );
  BUFFD0 U3387 ( .I(n3402), .Z(n3401) );
  BUFFD0 U3388 ( .I(n3403), .Z(n3402) );
  BUFFD0 U3389 ( .I(n3404), .Z(n3403) );
  BUFFD0 U3390 ( .I(n3405), .Z(n3404) );
  BUFFD0 U3391 ( .I(n3406), .Z(n3405) );
  BUFFD0 U3392 ( .I(n3407), .Z(n3406) );
  BUFFD0 U3393 ( .I(n3408), .Z(n3407) );
  BUFFD0 U3394 ( .I(n3409), .Z(n3408) );
  BUFFD0 U3395 ( .I(n3410), .Z(n3409) );
  BUFFD0 U3396 ( .I(n3411), .Z(n3410) );
  BUFFD0 U3397 ( .I(n3412), .Z(n3411) );
  BUFFD0 U3398 ( .I(n3413), .Z(n3412) );
  BUFFD0 U3399 ( .I(n3414), .Z(n3413) );
  BUFFD0 U3400 ( .I(n3415), .Z(n3414) );
  BUFFD0 U3401 ( .I(n3416), .Z(n3415) );
  BUFFD0 U3402 ( .I(n3417), .Z(n3416) );
  BUFFD0 U3403 ( .I(n3418), .Z(n3417) );
  BUFFD0 U3404 ( .I(n3419), .Z(n3418) );
  BUFFD0 U3405 ( .I(n3420), .Z(n3419) );
  BUFFD0 U3406 ( .I(n3421), .Z(n3420) );
  BUFFD0 U3407 ( .I(n3422), .Z(n3421) );
  BUFFD0 U3408 ( .I(n3423), .Z(n3422) );
  BUFFD0 U3409 ( .I(n3424), .Z(n3423) );
  BUFFD0 U3410 ( .I(n3425), .Z(n3424) );
  BUFFD0 U3411 ( .I(n3426), .Z(n3425) );
  BUFFD0 U3412 ( .I(n3427), .Z(n3426) );
  BUFFD0 U3413 ( .I(n3428), .Z(n3427) );
  BUFFD0 U3414 ( .I(n3429), .Z(n3428) );
  BUFFD0 U3415 ( .I(n3430), .Z(n3429) );
  BUFFD0 U3416 ( .I(n3431), .Z(n3430) );
  BUFFD0 U3417 ( .I(n3432), .Z(n3431) );
  BUFFD0 U3418 ( .I(n3433), .Z(n3432) );
  BUFFD0 U3419 ( .I(n3434), .Z(n3433) );
  BUFFD0 U3420 ( .I(n3435), .Z(n3434) );
  BUFFD0 U3421 ( .I(n3436), .Z(n3435) );
  BUFFD0 U3422 ( .I(n3437), .Z(n3436) );
  BUFFD0 U3423 ( .I(n3438), .Z(n3437) );
  BUFFD0 U3424 ( .I(n3439), .Z(n3438) );
  BUFFD0 U3425 ( .I(n3440), .Z(n3439) );
  BUFFD0 U3426 ( .I(N75), .Z(n3440) );
  BUFFD0 U3427 ( .I(n3442), .Z(n3441) );
  BUFFD0 U3428 ( .I(n3443), .Z(n3442) );
  BUFFD0 U3429 ( .I(n3446), .Z(n3443) );
  BUFFD0 U3430 ( .I(n4064), .Z(n3444) );
  BUFFD0 U3431 ( .I(n3444), .Z(n3445) );
  BUFFD0 U3432 ( .I(n3447), .Z(n3446) );
  BUFFD0 U3433 ( .I(n3448), .Z(n3447) );
  BUFFD0 U3434 ( .I(n3449), .Z(n3448) );
  BUFFD0 U3435 ( .I(n3450), .Z(n3449) );
  BUFFD0 U3436 ( .I(n3451), .Z(n3450) );
  BUFFD0 U3437 ( .I(n3452), .Z(n3451) );
  BUFFD0 U3438 ( .I(n3453), .Z(n3452) );
  BUFFD0 U3439 ( .I(n3454), .Z(n3453) );
  BUFFD0 U3440 ( .I(n3455), .Z(n3454) );
  BUFFD0 U3441 ( .I(n3456), .Z(n3455) );
  BUFFD0 U3442 ( .I(n3457), .Z(n3456) );
  BUFFD0 U3443 ( .I(n3458), .Z(n3457) );
  BUFFD0 U3444 ( .I(n3459), .Z(n3458) );
  BUFFD0 U3445 ( .I(n3460), .Z(n3459) );
  BUFFD0 U3446 ( .I(n3461), .Z(n3460) );
  BUFFD0 U3447 ( .I(n3462), .Z(n3461) );
  BUFFD0 U3448 ( .I(n3463), .Z(n3462) );
  BUFFD0 U3449 ( .I(n3464), .Z(n3463) );
  BUFFD0 U3450 ( .I(n3465), .Z(n3464) );
  BUFFD0 U3451 ( .I(n3466), .Z(n3465) );
  BUFFD0 U3452 ( .I(n3467), .Z(n3466) );
  BUFFD0 U3453 ( .I(n3468), .Z(n3467) );
  BUFFD0 U3454 ( .I(n3469), .Z(n3468) );
  BUFFD0 U3455 ( .I(n3470), .Z(n3469) );
  BUFFD0 U3456 ( .I(n3471), .Z(n3470) );
  BUFFD0 U3457 ( .I(n3472), .Z(n3471) );
  BUFFD0 U3458 ( .I(n3473), .Z(n3472) );
  BUFFD0 U3459 ( .I(n3474), .Z(n3473) );
  BUFFD0 U3460 ( .I(n3475), .Z(n3474) );
  BUFFD0 U3461 ( .I(n3476), .Z(n3475) );
  BUFFD0 U3462 ( .I(n3477), .Z(n3476) );
  BUFFD0 U3463 ( .I(n3478), .Z(n3477) );
  BUFFD0 U3464 ( .I(n3479), .Z(n3478) );
  BUFFD0 U3465 ( .I(n3480), .Z(n3479) );
  BUFFD0 U3466 ( .I(n3481), .Z(n3480) );
  BUFFD0 U3467 ( .I(n3482), .Z(n3481) );
  BUFFD0 U3468 ( .I(n3483), .Z(n3482) );
  BUFFD0 U3469 ( .I(n3484), .Z(n3483) );
  BUFFD0 U3470 ( .I(n3485), .Z(n3484) );
  BUFFD0 U3471 ( .I(n3486), .Z(n3485) );
  BUFFD0 U3472 ( .I(n3487), .Z(n3486) );
  BUFFD0 U3473 ( .I(n3488), .Z(n3487) );
  BUFFD0 U3474 ( .I(n3489), .Z(n3488) );
  BUFFD0 U3475 ( .I(n3490), .Z(n3489) );
  BUFFD0 U3476 ( .I(n3491), .Z(n3490) );
  BUFFD0 U3477 ( .I(n3492), .Z(n3491) );
  BUFFD0 U3478 ( .I(n3493), .Z(n3492) );
  BUFFD0 U3479 ( .I(n3494), .Z(n3493) );
  BUFFD0 U3480 ( .I(n3495), .Z(n3494) );
  BUFFD0 U3481 ( .I(n3496), .Z(n3495) );
  BUFFD0 U3482 ( .I(n3497), .Z(n3496) );
  BUFFD0 U3483 ( .I(n3498), .Z(n3497) );
  BUFFD0 U3484 ( .I(n3499), .Z(n3498) );
  BUFFD0 U3485 ( .I(n3500), .Z(n3499) );
  BUFFD0 U3486 ( .I(n3501), .Z(n3500) );
  BUFFD0 U3487 ( .I(n3502), .Z(n3501) );
  BUFFD0 U3488 ( .I(n3503), .Z(n3502) );
  BUFFD0 U3489 ( .I(n3504), .Z(n3503) );
  BUFFD0 U3490 ( .I(n3505), .Z(n3504) );
  BUFFD0 U3491 ( .I(n3506), .Z(n3505) );
  BUFFD0 U3492 ( .I(n3508), .Z(n3506) );
  BUFFD0 U3493 ( .I(N76), .Z(n3507) );
  BUFFD0 U3494 ( .I(n3509), .Z(n3508) );
  BUFFD0 U3495 ( .I(n3445), .Z(n3509) );
  BUFFD0 U3496 ( .I(n3511), .Z(n3510) );
  BUFFD0 U3497 ( .I(n3512), .Z(n3511) );
  BUFFD0 U3498 ( .I(n3513), .Z(n3512) );
  BUFFD0 U3499 ( .I(n3514), .Z(n3513) );
  BUFFD0 U3500 ( .I(n3515), .Z(n3514) );
  BUFFD0 U3501 ( .I(n3516), .Z(n3515) );
  BUFFD0 U3502 ( .I(n3517), .Z(n3516) );
  BUFFD0 U3503 ( .I(n3518), .Z(n3517) );
  BUFFD0 U3504 ( .I(n3519), .Z(n3518) );
  BUFFD0 U3505 ( .I(n3520), .Z(n3519) );
  BUFFD0 U3506 ( .I(n3521), .Z(n3520) );
  BUFFD0 U3507 ( .I(n3522), .Z(n3521) );
  BUFFD0 U3508 ( .I(n3523), .Z(n3522) );
  BUFFD0 U3509 ( .I(n3524), .Z(n3523) );
  BUFFD0 U3510 ( .I(n3525), .Z(n3524) );
  BUFFD0 U3511 ( .I(n3526), .Z(n3525) );
  BUFFD0 U3512 ( .I(n3527), .Z(n3526) );
  BUFFD0 U3513 ( .I(n3528), .Z(n3527) );
  BUFFD0 U3514 ( .I(n3529), .Z(n3528) );
  BUFFD0 U3515 ( .I(n3530), .Z(n3529) );
  BUFFD0 U3516 ( .I(n3531), .Z(n3530) );
  BUFFD0 U3517 ( .I(n3532), .Z(n3531) );
  BUFFD0 U3518 ( .I(n3533), .Z(n3532) );
  BUFFD0 U3519 ( .I(n3534), .Z(n3533) );
  BUFFD0 U3520 ( .I(n3535), .Z(n3534) );
  BUFFD0 U3521 ( .I(n3536), .Z(n3535) );
  BUFFD0 U3522 ( .I(n3537), .Z(n3536) );
  BUFFD0 U3523 ( .I(n3538), .Z(n3537) );
  BUFFD0 U3524 ( .I(n3539), .Z(n3538) );
  BUFFD0 U3525 ( .I(n3540), .Z(n3539) );
  BUFFD0 U3526 ( .I(n3541), .Z(n3540) );
  BUFFD0 U3527 ( .I(n3542), .Z(n3541) );
  BUFFD0 U3528 ( .I(n3543), .Z(n3542) );
  BUFFD0 U3529 ( .I(n3544), .Z(n3543) );
  BUFFD0 U3530 ( .I(n3545), .Z(n3544) );
  BUFFD0 U3531 ( .I(n3546), .Z(n3545) );
  BUFFD0 U3532 ( .I(n3547), .Z(n3546) );
  BUFFD0 U3533 ( .I(n3548), .Z(n3547) );
  BUFFD0 U3534 ( .I(n3549), .Z(n3548) );
  BUFFD0 U3535 ( .I(n3550), .Z(n3549) );
  BUFFD0 U3536 ( .I(n3551), .Z(n3550) );
  BUFFD0 U3537 ( .I(n3552), .Z(n3551) );
  BUFFD0 U3538 ( .I(n3553), .Z(n3552) );
  BUFFD0 U3539 ( .I(n3554), .Z(n3553) );
  BUFFD0 U3540 ( .I(n3555), .Z(n3554) );
  BUFFD0 U3541 ( .I(n3556), .Z(n3555) );
  BUFFD0 U3542 ( .I(n3557), .Z(n3556) );
  BUFFD0 U3543 ( .I(n3558), .Z(n3557) );
  BUFFD0 U3544 ( .I(n3559), .Z(n3558) );
  BUFFD0 U3545 ( .I(n3560), .Z(n3559) );
  BUFFD0 U3546 ( .I(n3561), .Z(n3560) );
  BUFFD0 U3547 ( .I(n3562), .Z(n3561) );
  BUFFD0 U3548 ( .I(n3563), .Z(n3562) );
  BUFFD0 U3549 ( .I(n3564), .Z(n3563) );
  BUFFD0 U3550 ( .I(n3565), .Z(n3564) );
  BUFFD0 U3551 ( .I(n3566), .Z(n3565) );
  BUFFD0 U3552 ( .I(n3567), .Z(n3566) );
  BUFFD0 U3553 ( .I(n3568), .Z(n3567) );
  BUFFD0 U3554 ( .I(n3569), .Z(n3568) );
  BUFFD0 U3555 ( .I(n3570), .Z(n3569) );
  BUFFD0 U3556 ( .I(n3571), .Z(n3570) );
  BUFFD0 U3557 ( .I(n3572), .Z(n3571) );
  BUFFD0 U3558 ( .I(n3573), .Z(n3572) );
  BUFFD0 U3559 ( .I(n3574), .Z(n3573) );
  BUFFD0 U3560 ( .I(n3575), .Z(n3574) );
  BUFFD0 U3561 ( .I(n3576), .Z(n3575) );
  BUFFD0 U3562 ( .I(n3577), .Z(n3576) );
  BUFFD0 U3563 ( .I(n3578), .Z(n3577) );
  BUFFD0 U3564 ( .I(n3579), .Z(n3578) );
  BUFFD0 U3565 ( .I(N77), .Z(n3579) );
  BUFFD0 U3566 ( .I(n3581), .Z(n3580) );
  BUFFD0 U3567 ( .I(n3582), .Z(n3581) );
  BUFFD0 U3568 ( .I(n3583), .Z(n3582) );
  BUFFD0 U3569 ( .I(n3584), .Z(n3583) );
  BUFFD0 U3570 ( .I(n3585), .Z(n3584) );
  BUFFD0 U3571 ( .I(n3586), .Z(n3585) );
  BUFFD0 U3572 ( .I(n3587), .Z(n3586) );
  BUFFD0 U3573 ( .I(n3588), .Z(n3587) );
  BUFFD0 U3574 ( .I(n3589), .Z(n3588) );
  BUFFD0 U3575 ( .I(n3590), .Z(n3589) );
  BUFFD0 U3576 ( .I(n3591), .Z(n3590) );
  BUFFD0 U3577 ( .I(n3592), .Z(n3591) );
  BUFFD0 U3578 ( .I(n3593), .Z(n3592) );
  BUFFD0 U3579 ( .I(n3594), .Z(n3593) );
  BUFFD0 U3580 ( .I(n3595), .Z(n3594) );
  BUFFD0 U3581 ( .I(n3596), .Z(n3595) );
  BUFFD0 U3582 ( .I(n3597), .Z(n3596) );
  BUFFD0 U3583 ( .I(n3598), .Z(n3597) );
  BUFFD0 U3584 ( .I(n3599), .Z(n3598) );
  BUFFD0 U3585 ( .I(n3600), .Z(n3599) );
  BUFFD0 U3586 ( .I(n3601), .Z(n3600) );
  BUFFD0 U3587 ( .I(n3602), .Z(n3601) );
  BUFFD0 U3588 ( .I(n3603), .Z(n3602) );
  BUFFD0 U3589 ( .I(n3604), .Z(n3603) );
  BUFFD0 U3590 ( .I(n3605), .Z(n3604) );
  BUFFD0 U3591 ( .I(n3606), .Z(n3605) );
  BUFFD0 U3592 ( .I(n3607), .Z(n3606) );
  BUFFD0 U3593 ( .I(n3608), .Z(n3607) );
  BUFFD0 U3594 ( .I(n3609), .Z(n3608) );
  BUFFD0 U3595 ( .I(n3610), .Z(n3609) );
  BUFFD0 U3596 ( .I(n3611), .Z(n3610) );
  BUFFD0 U3597 ( .I(n3612), .Z(n3611) );
  BUFFD0 U3598 ( .I(n3613), .Z(n3612) );
  BUFFD0 U3599 ( .I(n3614), .Z(n3613) );
  BUFFD0 U3600 ( .I(n3615), .Z(n3614) );
  BUFFD0 U3601 ( .I(n3616), .Z(n3615) );
  BUFFD0 U3602 ( .I(n3617), .Z(n3616) );
  BUFFD0 U3603 ( .I(n3618), .Z(n3617) );
  BUFFD0 U3604 ( .I(n3619), .Z(n3618) );
  BUFFD0 U3605 ( .I(n3620), .Z(n3619) );
  BUFFD0 U3606 ( .I(n3621), .Z(n3620) );
  BUFFD0 U3607 ( .I(n3622), .Z(n3621) );
  BUFFD0 U3608 ( .I(n3623), .Z(n3622) );
  BUFFD0 U3609 ( .I(n3624), .Z(n3623) );
  BUFFD0 U3610 ( .I(n3625), .Z(n3624) );
  BUFFD0 U3611 ( .I(n3626), .Z(n3625) );
  BUFFD0 U3612 ( .I(n3627), .Z(n3626) );
  BUFFD0 U3613 ( .I(n3628), .Z(n3627) );
  BUFFD0 U3614 ( .I(n3629), .Z(n3628) );
  BUFFD0 U3615 ( .I(n3630), .Z(n3629) );
  BUFFD0 U3616 ( .I(n3631), .Z(n3630) );
  BUFFD0 U3617 ( .I(n3632), .Z(n3631) );
  BUFFD0 U3618 ( .I(n3633), .Z(n3632) );
  BUFFD0 U3619 ( .I(n3634), .Z(n3633) );
  BUFFD0 U3620 ( .I(n3635), .Z(n3634) );
  BUFFD0 U3621 ( .I(n3636), .Z(n3635) );
  BUFFD0 U3622 ( .I(n3637), .Z(n3636) );
  BUFFD0 U3623 ( .I(n3638), .Z(n3637) );
  BUFFD0 U3624 ( .I(n3639), .Z(n3638) );
  BUFFD0 U3625 ( .I(n3640), .Z(n3639) );
  BUFFD0 U3626 ( .I(n3641), .Z(n3640) );
  BUFFD0 U3627 ( .I(n3642), .Z(n3641) );
  BUFFD0 U3628 ( .I(n3643), .Z(n3642) );
  BUFFD0 U3629 ( .I(n3644), .Z(n3643) );
  BUFFD0 U3630 ( .I(n3645), .Z(n3644) );
  BUFFD0 U3631 ( .I(n3646), .Z(n3645) );
  BUFFD0 U3632 ( .I(n3647), .Z(n3646) );
  BUFFD0 U3633 ( .I(n3648), .Z(n3647) );
  BUFFD0 U3634 ( .I(n3649), .Z(n3648) );
  BUFFD0 U3635 ( .I(N78), .Z(n3649) );
  BUFFD0 U3636 ( .I(n3651), .Z(n3650) );
  BUFFD0 U3637 ( .I(n3652), .Z(n3651) );
  BUFFD0 U3638 ( .I(n3653), .Z(n3652) );
  BUFFD0 U3639 ( .I(n3654), .Z(n3653) );
  BUFFD0 U3640 ( .I(n3655), .Z(n3654) );
  BUFFD0 U3641 ( .I(n3656), .Z(n3655) );
  BUFFD0 U3642 ( .I(n3657), .Z(n3656) );
  BUFFD0 U3643 ( .I(n3658), .Z(n3657) );
  BUFFD0 U3644 ( .I(n3659), .Z(n3658) );
  BUFFD0 U3645 ( .I(n3660), .Z(n3659) );
  BUFFD0 U3646 ( .I(n3661), .Z(n3660) );
  BUFFD0 U3647 ( .I(n3662), .Z(n3661) );
  BUFFD0 U3648 ( .I(n3663), .Z(n3662) );
  BUFFD0 U3649 ( .I(n3664), .Z(n3663) );
  BUFFD0 U3650 ( .I(n3665), .Z(n3664) );
  BUFFD0 U3651 ( .I(n3666), .Z(n3665) );
  BUFFD0 U3652 ( .I(n3667), .Z(n3666) );
  BUFFD0 U3653 ( .I(n3668), .Z(n3667) );
  BUFFD0 U3654 ( .I(n3669), .Z(n3668) );
  BUFFD0 U3655 ( .I(n3670), .Z(n3669) );
  BUFFD0 U3656 ( .I(n3671), .Z(n3670) );
  BUFFD0 U3657 ( .I(n3672), .Z(n3671) );
  BUFFD0 U3658 ( .I(n3673), .Z(n3672) );
  BUFFD0 U3659 ( .I(n3674), .Z(n3673) );
  BUFFD0 U3660 ( .I(n3675), .Z(n3674) );
  BUFFD0 U3661 ( .I(n3676), .Z(n3675) );
  BUFFD0 U3662 ( .I(n3677), .Z(n3676) );
  BUFFD0 U3663 ( .I(n3678), .Z(n3677) );
  BUFFD0 U3664 ( .I(n3679), .Z(n3678) );
  BUFFD0 U3665 ( .I(n3680), .Z(n3679) );
  BUFFD0 U3666 ( .I(n3681), .Z(n3680) );
  BUFFD0 U3667 ( .I(n3682), .Z(n3681) );
  BUFFD0 U3668 ( .I(n3683), .Z(n3682) );
  BUFFD0 U3669 ( .I(n3684), .Z(n3683) );
  BUFFD0 U3670 ( .I(n3685), .Z(n3684) );
  BUFFD0 U3671 ( .I(n3686), .Z(n3685) );
  BUFFD0 U3672 ( .I(n3687), .Z(n3686) );
  BUFFD0 U3673 ( .I(n3688), .Z(n3687) );
  BUFFD0 U3674 ( .I(n3689), .Z(n3688) );
  BUFFD0 U3675 ( .I(n3690), .Z(n3689) );
  BUFFD0 U3676 ( .I(n3691), .Z(n3690) );
  BUFFD0 U3677 ( .I(n3692), .Z(n3691) );
  BUFFD0 U3678 ( .I(n3693), .Z(n3692) );
  BUFFD0 U3679 ( .I(n3694), .Z(n3693) );
  BUFFD0 U3680 ( .I(n3695), .Z(n3694) );
  BUFFD0 U3681 ( .I(n3696), .Z(n3695) );
  BUFFD0 U3682 ( .I(n3697), .Z(n3696) );
  BUFFD0 U3683 ( .I(n3698), .Z(n3697) );
  BUFFD0 U3684 ( .I(n3699), .Z(n3698) );
  BUFFD0 U3685 ( .I(n3700), .Z(n3699) );
  BUFFD0 U3686 ( .I(n3701), .Z(n3700) );
  BUFFD0 U3687 ( .I(n3702), .Z(n3701) );
  BUFFD0 U3688 ( .I(n3703), .Z(n3702) );
  BUFFD0 U3689 ( .I(n3704), .Z(n3703) );
  BUFFD0 U3690 ( .I(n3705), .Z(n3704) );
  BUFFD0 U3691 ( .I(n3706), .Z(n3705) );
  BUFFD0 U3692 ( .I(n3707), .Z(n3706) );
  BUFFD0 U3693 ( .I(n3708), .Z(n3707) );
  BUFFD0 U3694 ( .I(n3709), .Z(n3708) );
  BUFFD0 U3695 ( .I(n3710), .Z(n3709) );
  BUFFD0 U3696 ( .I(n3711), .Z(n3710) );
  BUFFD0 U3697 ( .I(n3712), .Z(n3711) );
  BUFFD0 U3698 ( .I(n3713), .Z(n3712) );
  BUFFD0 U3699 ( .I(n3714), .Z(n3713) );
  BUFFD0 U3700 ( .I(n3715), .Z(n3714) );
  BUFFD0 U3701 ( .I(n3716), .Z(n3715) );
  BUFFD0 U3702 ( .I(n3717), .Z(n3716) );
  BUFFD0 U3703 ( .I(n3718), .Z(n3717) );
  BUFFD0 U3704 ( .I(n3719), .Z(n3718) );
  BUFFD0 U3705 ( .I(N79), .Z(n3719) );
  BUFFD0 U3706 ( .I(n3721), .Z(n3720) );
  BUFFD0 U3707 ( .I(n3722), .Z(n3721) );
  BUFFD0 U3708 ( .I(n3723), .Z(n3722) );
  BUFFD0 U3709 ( .I(n3724), .Z(n3723) );
  BUFFD0 U3710 ( .I(n3725), .Z(n3724) );
  BUFFD0 U3711 ( .I(n3726), .Z(n3725) );
  BUFFD0 U3712 ( .I(n3727), .Z(n3726) );
  BUFFD0 U3713 ( .I(n3728), .Z(n3727) );
  BUFFD0 U3714 ( .I(n3729), .Z(n3728) );
  BUFFD0 U3715 ( .I(n3730), .Z(n3729) );
  BUFFD0 U3716 ( .I(n3731), .Z(n3730) );
  BUFFD0 U3717 ( .I(n3732), .Z(n3731) );
  BUFFD0 U3718 ( .I(n3733), .Z(n3732) );
  BUFFD0 U3719 ( .I(n3734), .Z(n3733) );
  BUFFD0 U3720 ( .I(n3735), .Z(n3734) );
  BUFFD0 U3721 ( .I(n3736), .Z(n3735) );
  BUFFD0 U3722 ( .I(n3737), .Z(n3736) );
  BUFFD0 U3723 ( .I(n3738), .Z(n3737) );
  BUFFD0 U3724 ( .I(n3739), .Z(n3738) );
  BUFFD0 U3725 ( .I(n3740), .Z(n3739) );
  BUFFD0 U3726 ( .I(n3741), .Z(n3740) );
  BUFFD0 U3727 ( .I(n3742), .Z(n3741) );
  BUFFD0 U3728 ( .I(n3743), .Z(n3742) );
  BUFFD0 U3729 ( .I(n3744), .Z(n3743) );
  BUFFD0 U3730 ( .I(n3745), .Z(n3744) );
  BUFFD0 U3731 ( .I(n3746), .Z(n3745) );
  BUFFD0 U3732 ( .I(n3747), .Z(n3746) );
  BUFFD0 U3733 ( .I(n3748), .Z(n3747) );
  BUFFD0 U3734 ( .I(n3749), .Z(n3748) );
  BUFFD0 U3735 ( .I(n3750), .Z(n3749) );
  BUFFD0 U3736 ( .I(n3751), .Z(n3750) );
  BUFFD0 U3737 ( .I(n3752), .Z(n3751) );
  BUFFD0 U3738 ( .I(n3753), .Z(n3752) );
  BUFFD0 U3739 ( .I(n3754), .Z(n3753) );
  BUFFD0 U3740 ( .I(n3755), .Z(n3754) );
  BUFFD0 U3741 ( .I(n3756), .Z(n3755) );
  BUFFD0 U3742 ( .I(n3757), .Z(n3756) );
  BUFFD0 U3743 ( .I(n3758), .Z(n3757) );
  BUFFD0 U3744 ( .I(n3759), .Z(n3758) );
  BUFFD0 U3745 ( .I(n3760), .Z(n3759) );
  BUFFD0 U3746 ( .I(n3761), .Z(n3760) );
  BUFFD0 U3747 ( .I(n3762), .Z(n3761) );
  BUFFD0 U3748 ( .I(n3763), .Z(n3762) );
  BUFFD0 U3749 ( .I(n3764), .Z(n3763) );
  BUFFD0 U3750 ( .I(n3765), .Z(n3764) );
  BUFFD0 U3751 ( .I(n3766), .Z(n3765) );
  BUFFD0 U3752 ( .I(n3767), .Z(n3766) );
  BUFFD0 U3753 ( .I(n3768), .Z(n3767) );
  BUFFD0 U3754 ( .I(n3769), .Z(n3768) );
  BUFFD0 U3755 ( .I(n3770), .Z(n3769) );
  BUFFD0 U3756 ( .I(n3771), .Z(n3770) );
  BUFFD0 U3757 ( .I(n3772), .Z(n3771) );
  BUFFD0 U3758 ( .I(n3773), .Z(n3772) );
  BUFFD0 U3759 ( .I(n3774), .Z(n3773) );
  BUFFD0 U3760 ( .I(n3775), .Z(n3774) );
  BUFFD0 U3761 ( .I(n3776), .Z(n3775) );
  BUFFD0 U3762 ( .I(n3777), .Z(n3776) );
  BUFFD0 U3763 ( .I(n3778), .Z(n3777) );
  BUFFD0 U3764 ( .I(n3779), .Z(n3778) );
  BUFFD0 U3765 ( .I(n3780), .Z(n3779) );
  BUFFD0 U3766 ( .I(n3781), .Z(n3780) );
  BUFFD0 U3767 ( .I(n3782), .Z(n3781) );
  BUFFD0 U3768 ( .I(n3783), .Z(n3782) );
  BUFFD0 U3769 ( .I(n3784), .Z(n3783) );
  BUFFD0 U3770 ( .I(n3785), .Z(n3784) );
  BUFFD0 U3771 ( .I(n3786), .Z(n3785) );
  BUFFD0 U3772 ( .I(n3787), .Z(n3786) );
  BUFFD0 U3773 ( .I(n3788), .Z(n3787) );
  BUFFD0 U3774 ( .I(N80), .Z(n3788) );
  CKBD0 U3775 ( .CLK(n3790), .C(n3854) );
  BUFFD0 U3776 ( .I(n3793), .Z(n3789) );
  BUFFD0 U3777 ( .I(N81), .Z(n3790) );
  BUFFD0 U3778 ( .I(n4065), .Z(n3791) );
  BUFFD0 U3779 ( .I(n3791), .Z(n3792) );
  BUFFD0 U3780 ( .I(n3794), .Z(n3793) );
  BUFFD0 U3781 ( .I(n3795), .Z(n3794) );
  BUFFD0 U3782 ( .I(n3796), .Z(n3795) );
  BUFFD0 U3783 ( .I(n3797), .Z(n3796) );
  BUFFD0 U3784 ( .I(n3798), .Z(n3797) );
  BUFFD0 U3785 ( .I(n3799), .Z(n3798) );
  BUFFD0 U3786 ( .I(n3800), .Z(n3799) );
  BUFFD0 U3787 ( .I(n3801), .Z(n3800) );
  BUFFD0 U3788 ( .I(n3802), .Z(n3801) );
  BUFFD0 U3789 ( .I(n3803), .Z(n3802) );
  BUFFD0 U3790 ( .I(n3804), .Z(n3803) );
  BUFFD0 U3791 ( .I(n3805), .Z(n3804) );
  BUFFD0 U3792 ( .I(n3806), .Z(n3805) );
  BUFFD0 U3793 ( .I(n3807), .Z(n3806) );
  BUFFD0 U3794 ( .I(n3808), .Z(n3807) );
  BUFFD0 U3795 ( .I(n3809), .Z(n3808) );
  BUFFD0 U3796 ( .I(n3810), .Z(n3809) );
  BUFFD0 U3797 ( .I(n3811), .Z(n3810) );
  BUFFD0 U3798 ( .I(n3812), .Z(n3811) );
  BUFFD0 U3799 ( .I(n3813), .Z(n3812) );
  BUFFD0 U3800 ( .I(n3814), .Z(n3813) );
  BUFFD0 U3801 ( .I(n3815), .Z(n3814) );
  BUFFD0 U3802 ( .I(n3816), .Z(n3815) );
  BUFFD0 U3803 ( .I(n3817), .Z(n3816) );
  BUFFD0 U3804 ( .I(n3818), .Z(n3817) );
  BUFFD0 U3805 ( .I(n3819), .Z(n3818) );
  BUFFD0 U3806 ( .I(n3820), .Z(n3819) );
  BUFFD0 U3807 ( .I(n3821), .Z(n3820) );
  BUFFD0 U3808 ( .I(n3822), .Z(n3821) );
  BUFFD0 U3809 ( .I(n3823), .Z(n3822) );
  BUFFD0 U3810 ( .I(n3824), .Z(n3823) );
  BUFFD0 U3811 ( .I(n3825), .Z(n3824) );
  BUFFD0 U3812 ( .I(n3826), .Z(n3825) );
  BUFFD0 U3813 ( .I(n3827), .Z(n3826) );
  BUFFD0 U3814 ( .I(n3828), .Z(n3827) );
  BUFFD0 U3815 ( .I(n3829), .Z(n3828) );
  BUFFD0 U3816 ( .I(n3830), .Z(n3829) );
  BUFFD0 U3817 ( .I(n3831), .Z(n3830) );
  BUFFD0 U3818 ( .I(n3832), .Z(n3831) );
  BUFFD0 U3819 ( .I(n3833), .Z(n3832) );
  BUFFD0 U3820 ( .I(n3834), .Z(n3833) );
  BUFFD0 U3821 ( .I(n3835), .Z(n3834) );
  BUFFD0 U3822 ( .I(n3836), .Z(n3835) );
  BUFFD0 U3823 ( .I(n3837), .Z(n3836) );
  BUFFD0 U3824 ( .I(n3838), .Z(n3837) );
  BUFFD0 U3825 ( .I(n3839), .Z(n3838) );
  BUFFD0 U3826 ( .I(n3840), .Z(n3839) );
  BUFFD0 U3827 ( .I(n3841), .Z(n3840) );
  BUFFD0 U3828 ( .I(n3842), .Z(n3841) );
  BUFFD0 U3829 ( .I(n3843), .Z(n3842) );
  BUFFD0 U3830 ( .I(n3844), .Z(n3843) );
  BUFFD0 U3831 ( .I(n3845), .Z(n3844) );
  BUFFD0 U3832 ( .I(n3846), .Z(n3845) );
  BUFFD0 U3833 ( .I(n3847), .Z(n3846) );
  BUFFD0 U3834 ( .I(n3848), .Z(n3847) );
  BUFFD0 U3835 ( .I(n3849), .Z(n3848) );
  BUFFD0 U3836 ( .I(n3850), .Z(n3849) );
  BUFFD0 U3837 ( .I(n3851), .Z(n3850) );
  BUFFD0 U3838 ( .I(n3852), .Z(n3851) );
  BUFFD0 U3839 ( .I(n3853), .Z(n3852) );
  BUFFD0 U3840 ( .I(n3855), .Z(n3853) );
  BUFFD0 U3841 ( .I(n3856), .Z(n3855) );
  BUFFD0 U3842 ( .I(n3792), .Z(n3856) );
  BUFFD0 U3843 ( .I(n3858), .Z(n3857) );
  BUFFD0 U3844 ( .I(n3859), .Z(n3858) );
  BUFFD0 U3845 ( .I(n3860), .Z(n3859) );
  BUFFD0 U3846 ( .I(n3861), .Z(n3860) );
  BUFFD0 U3847 ( .I(n3862), .Z(n3861) );
  BUFFD0 U3848 ( .I(n3863), .Z(n3862) );
  BUFFD0 U3849 ( .I(n3864), .Z(n3863) );
  BUFFD0 U3850 ( .I(n3865), .Z(n3864) );
  BUFFD0 U3851 ( .I(n3866), .Z(n3865) );
  BUFFD0 U3852 ( .I(n3867), .Z(n3866) );
  BUFFD0 U3853 ( .I(n3868), .Z(n3867) );
  BUFFD0 U3854 ( .I(n3869), .Z(n3868) );
  BUFFD0 U3855 ( .I(n3870), .Z(n3869) );
  BUFFD0 U3856 ( .I(n3871), .Z(n3870) );
  BUFFD0 U3857 ( .I(n3872), .Z(n3871) );
  BUFFD0 U3858 ( .I(n3873), .Z(n3872) );
  BUFFD0 U3859 ( .I(n3874), .Z(n3873) );
  BUFFD0 U3860 ( .I(n3875), .Z(n3874) );
  BUFFD0 U3861 ( .I(n3876), .Z(n3875) );
  BUFFD0 U3862 ( .I(n3877), .Z(n3876) );
  BUFFD0 U3863 ( .I(n3878), .Z(n3877) );
  BUFFD0 U3864 ( .I(n3879), .Z(n3878) );
  BUFFD0 U3865 ( .I(n3880), .Z(n3879) );
  BUFFD0 U3866 ( .I(n3881), .Z(n3880) );
  BUFFD0 U3867 ( .I(n3882), .Z(n3881) );
  BUFFD0 U3868 ( .I(n3883), .Z(n3882) );
  BUFFD0 U3869 ( .I(n3884), .Z(n3883) );
  BUFFD0 U3870 ( .I(n3885), .Z(n3884) );
  BUFFD0 U3871 ( .I(n3886), .Z(n3885) );
  BUFFD0 U3872 ( .I(n3887), .Z(n3886) );
  BUFFD0 U3873 ( .I(n3888), .Z(n3887) );
  BUFFD0 U3874 ( .I(n3889), .Z(n3888) );
  BUFFD0 U3875 ( .I(n3890), .Z(n3889) );
  BUFFD0 U3876 ( .I(n3891), .Z(n3890) );
  BUFFD0 U3877 ( .I(n3892), .Z(n3891) );
  BUFFD0 U3878 ( .I(n3893), .Z(n3892) );
  BUFFD0 U3879 ( .I(n3894), .Z(n3893) );
  BUFFD0 U3880 ( .I(n3895), .Z(n3894) );
  BUFFD0 U3881 ( .I(n3896), .Z(n3895) );
  BUFFD0 U3882 ( .I(n3897), .Z(n3896) );
  BUFFD0 U3883 ( .I(n3898), .Z(n3897) );
  BUFFD0 U3884 ( .I(n3899), .Z(n3898) );
  BUFFD0 U3885 ( .I(n3900), .Z(n3899) );
  BUFFD0 U3886 ( .I(n3901), .Z(n3900) );
  BUFFD0 U3887 ( .I(n3902), .Z(n3901) );
  BUFFD0 U3888 ( .I(n3903), .Z(n3902) );
  BUFFD0 U3889 ( .I(n3904), .Z(n3903) );
  BUFFD0 U3890 ( .I(n3905), .Z(n3904) );
  BUFFD0 U3891 ( .I(n3906), .Z(n3905) );
  BUFFD0 U3892 ( .I(n3907), .Z(n3906) );
  BUFFD0 U3893 ( .I(n3908), .Z(n3907) );
  BUFFD0 U3894 ( .I(n3909), .Z(n3908) );
  BUFFD0 U3895 ( .I(n3910), .Z(n3909) );
  BUFFD0 U3896 ( .I(n3911), .Z(n3910) );
  BUFFD0 U3897 ( .I(n3912), .Z(n3911) );
  BUFFD0 U3898 ( .I(n3913), .Z(n3912) );
  BUFFD0 U3899 ( .I(n3914), .Z(n3913) );
  BUFFD0 U3900 ( .I(n3915), .Z(n3914) );
  BUFFD0 U3901 ( .I(n3916), .Z(n3915) );
  BUFFD0 U3902 ( .I(n3917), .Z(n3916) );
  BUFFD0 U3903 ( .I(n3918), .Z(n3917) );
  BUFFD0 U3904 ( .I(n3919), .Z(n3918) );
  BUFFD0 U3905 ( .I(n3920), .Z(n3919) );
  BUFFD0 U3906 ( .I(n3921), .Z(n3920) );
  BUFFD0 U3907 ( .I(n3922), .Z(n3921) );
  BUFFD0 U3908 ( .I(n3923), .Z(n3922) );
  BUFFD0 U3909 ( .I(n3924), .Z(n3923) );
  BUFFD0 U3910 ( .I(n3925), .Z(n3924) );
  BUFFD0 U3911 ( .I(N82), .Z(n3925) );
  BUFFD0 U3912 ( .I(n3927), .Z(n3926) );
  BUFFD0 U3913 ( .I(n3928), .Z(n3927) );
  BUFFD0 U3914 ( .I(n3929), .Z(n3928) );
  BUFFD0 U3915 ( .I(n3930), .Z(n3929) );
  BUFFD0 U3916 ( .I(n3931), .Z(n3930) );
  BUFFD0 U3917 ( .I(n3932), .Z(n3931) );
  BUFFD0 U3918 ( .I(n3933), .Z(n3932) );
  BUFFD0 U3919 ( .I(n3934), .Z(n3933) );
  BUFFD0 U3920 ( .I(n3935), .Z(n3934) );
  BUFFD0 U3921 ( .I(n3936), .Z(n3935) );
  BUFFD0 U3922 ( .I(n3937), .Z(n3936) );
  BUFFD0 U3923 ( .I(n3938), .Z(n3937) );
  BUFFD0 U3924 ( .I(n3939), .Z(n3938) );
  BUFFD0 U3925 ( .I(n3940), .Z(n3939) );
  BUFFD0 U3926 ( .I(n3941), .Z(n3940) );
  BUFFD0 U3927 ( .I(n3942), .Z(n3941) );
  BUFFD0 U3928 ( .I(n3943), .Z(n3942) );
  BUFFD0 U3929 ( .I(n3944), .Z(n3943) );
  BUFFD0 U3930 ( .I(n3945), .Z(n3944) );
  BUFFD0 U3931 ( .I(n3946), .Z(n3945) );
  BUFFD0 U3932 ( .I(n3947), .Z(n3946) );
  BUFFD0 U3933 ( .I(n3948), .Z(n3947) );
  BUFFD0 U3934 ( .I(n3949), .Z(n3948) );
  BUFFD0 U3935 ( .I(n3950), .Z(n3949) );
  BUFFD0 U3936 ( .I(n3951), .Z(n3950) );
  BUFFD0 U3937 ( .I(n3952), .Z(n3951) );
  BUFFD0 U3938 ( .I(n3953), .Z(n3952) );
  BUFFD0 U3939 ( .I(n3954), .Z(n3953) );
  BUFFD0 U3940 ( .I(n3955), .Z(n3954) );
  BUFFD0 U3941 ( .I(n3956), .Z(n3955) );
  BUFFD0 U3942 ( .I(n3957), .Z(n3956) );
  BUFFD0 U3943 ( .I(n3958), .Z(n3957) );
  BUFFD0 U3944 ( .I(n3959), .Z(n3958) );
  BUFFD0 U3945 ( .I(n3960), .Z(n3959) );
  BUFFD0 U3946 ( .I(n3961), .Z(n3960) );
  BUFFD0 U3947 ( .I(n3962), .Z(n3961) );
  BUFFD0 U3948 ( .I(n3963), .Z(n3962) );
  BUFFD0 U3949 ( .I(n3964), .Z(n3963) );
  BUFFD0 U3950 ( .I(n3965), .Z(n3964) );
  BUFFD0 U3951 ( .I(n3966), .Z(n3965) );
  BUFFD0 U3952 ( .I(n3967), .Z(n3966) );
  BUFFD0 U3953 ( .I(n3968), .Z(n3967) );
  BUFFD0 U3954 ( .I(n3969), .Z(n3968) );
  BUFFD0 U3955 ( .I(n3970), .Z(n3969) );
  BUFFD0 U3956 ( .I(n3971), .Z(n3970) );
  BUFFD0 U3957 ( .I(n3972), .Z(n3971) );
  BUFFD0 U3958 ( .I(n3973), .Z(n3972) );
  BUFFD0 U3959 ( .I(n3974), .Z(n3973) );
  BUFFD0 U3960 ( .I(n3975), .Z(n3974) );
  BUFFD0 U3961 ( .I(n3976), .Z(n3975) );
  BUFFD0 U3962 ( .I(n3977), .Z(n3976) );
  BUFFD0 U3963 ( .I(n3978), .Z(n3977) );
  BUFFD0 U3964 ( .I(n3979), .Z(n3978) );
  BUFFD0 U3965 ( .I(n3980), .Z(n3979) );
  BUFFD0 U3966 ( .I(n3981), .Z(n3980) );
  BUFFD0 U3967 ( .I(n3982), .Z(n3981) );
  BUFFD0 U3968 ( .I(n3983), .Z(n3982) );
  BUFFD0 U3969 ( .I(n3984), .Z(n3983) );
  BUFFD0 U3970 ( .I(n3985), .Z(n3984) );
  BUFFD0 U3971 ( .I(n3986), .Z(n3985) );
  BUFFD0 U3972 ( .I(n3987), .Z(n3986) );
  BUFFD0 U3973 ( .I(n3988), .Z(n3987) );
  BUFFD0 U3974 ( .I(n3989), .Z(n3988) );
  BUFFD0 U3975 ( .I(n3990), .Z(n3989) );
  BUFFD0 U3976 ( .I(n3991), .Z(n3990) );
  BUFFD0 U3977 ( .I(n3992), .Z(n3991) );
  BUFFD0 U3978 ( .I(n3993), .Z(n3992) );
  BUFFD0 U3979 ( .I(n3994), .Z(n3993) );
  BUFFD0 U3980 ( .I(N83), .Z(n3994) );
  BUFFD0 U3981 ( .I(n3996), .Z(n3995) );
  BUFFD0 U3982 ( .I(n3997), .Z(n3996) );
  BUFFD0 U3983 ( .I(n3998), .Z(n3997) );
  BUFFD0 U3984 ( .I(n3999), .Z(n3998) );
  BUFFD0 U3985 ( .I(n4000), .Z(n3999) );
  BUFFD0 U3986 ( .I(n4001), .Z(n4000) );
  BUFFD0 U3987 ( .I(n4002), .Z(n4001) );
  BUFFD0 U3988 ( .I(n4003), .Z(n4002) );
  BUFFD0 U3989 ( .I(n4004), .Z(n4003) );
  BUFFD0 U3990 ( .I(n4005), .Z(n4004) );
  BUFFD0 U3991 ( .I(n4006), .Z(n4005) );
  BUFFD0 U3992 ( .I(n4007), .Z(n4006) );
  BUFFD0 U3993 ( .I(n4008), .Z(n4007) );
  BUFFD0 U3994 ( .I(n4009), .Z(n4008) );
  BUFFD0 U3995 ( .I(n4010), .Z(n4009) );
  BUFFD0 U3996 ( .I(n4011), .Z(n4010) );
  BUFFD0 U3997 ( .I(n4012), .Z(n4011) );
  BUFFD0 U3998 ( .I(n4013), .Z(n4012) );
  BUFFD0 U3999 ( .I(n4014), .Z(n4013) );
  BUFFD0 U4000 ( .I(n4015), .Z(n4014) );
  BUFFD0 U4001 ( .I(n4016), .Z(n4015) );
  BUFFD0 U4002 ( .I(n4017), .Z(n4016) );
  BUFFD0 U4003 ( .I(n4018), .Z(n4017) );
  BUFFD0 U4004 ( .I(n4019), .Z(n4018) );
  BUFFD0 U4005 ( .I(n4020), .Z(n4019) );
  BUFFD0 U4006 ( .I(n4021), .Z(n4020) );
  BUFFD0 U4007 ( .I(n4022), .Z(n4021) );
  BUFFD0 U4008 ( .I(n4023), .Z(n4022) );
  BUFFD0 U4009 ( .I(n4024), .Z(n4023) );
  BUFFD0 U4010 ( .I(n4025), .Z(n4024) );
  BUFFD0 U4011 ( .I(n4026), .Z(n4025) );
  BUFFD0 U4012 ( .I(n4027), .Z(n4026) );
  BUFFD0 U4013 ( .I(n4028), .Z(n4027) );
  BUFFD0 U4014 ( .I(n4029), .Z(n4028) );
  BUFFD0 U4015 ( .I(n4030), .Z(n4029) );
  BUFFD0 U4016 ( .I(n4031), .Z(n4030) );
  BUFFD0 U4017 ( .I(n4032), .Z(n4031) );
  BUFFD0 U4018 ( .I(n4033), .Z(n4032) );
  BUFFD0 U4019 ( .I(n4034), .Z(n4033) );
  BUFFD0 U4020 ( .I(n4035), .Z(n4034) );
  BUFFD0 U4021 ( .I(n4036), .Z(n4035) );
  BUFFD0 U4022 ( .I(n4037), .Z(n4036) );
  BUFFD0 U4023 ( .I(n4038), .Z(n4037) );
  BUFFD0 U4024 ( .I(n4039), .Z(n4038) );
  BUFFD0 U4025 ( .I(n4040), .Z(n4039) );
  BUFFD0 U4026 ( .I(n4041), .Z(n4040) );
  BUFFD0 U4027 ( .I(n4042), .Z(n4041) );
  BUFFD0 U4028 ( .I(n4043), .Z(n4042) );
  BUFFD0 U4029 ( .I(n4044), .Z(n4043) );
  BUFFD0 U4030 ( .I(n4045), .Z(n4044) );
  BUFFD0 U4031 ( .I(n4046), .Z(n4045) );
  BUFFD0 U4032 ( .I(n4047), .Z(n4046) );
  BUFFD0 U4033 ( .I(n4048), .Z(n4047) );
  BUFFD0 U4034 ( .I(n4049), .Z(n4048) );
  BUFFD0 U4035 ( .I(n4050), .Z(n4049) );
  BUFFD0 U4036 ( .I(n4051), .Z(n4050) );
  BUFFD0 U4037 ( .I(n4052), .Z(n4051) );
  BUFFD0 U4038 ( .I(n4053), .Z(n4052) );
  BUFFD0 U4039 ( .I(n4054), .Z(n4053) );
  BUFFD0 U4040 ( .I(n4055), .Z(n4054) );
  BUFFD0 U4041 ( .I(n4056), .Z(n4055) );
  BUFFD0 U4042 ( .I(n4057), .Z(n4056) );
  BUFFD0 U4043 ( .I(n4058), .Z(n4057) );
  BUFFD0 U4044 ( .I(n4059), .Z(n4058) );
  BUFFD0 U4045 ( .I(n4060), .Z(n4059) );
  BUFFD0 U4046 ( .I(n4061), .Z(n4060) );
  BUFFD0 U4047 ( .I(n4062), .Z(n4061) );
  BUFFD0 U4048 ( .I(n4063), .Z(n4062) );
  BUFFD0 U4049 ( .I(N84), .Z(n4063) );
  BUFFD0 U4050 ( .I(n3507), .Z(n4064) );
  BUFFD0 U4051 ( .I(n3854), .Z(n4065) );
  BUFFD0 U4052 ( .I(n4067), .Z(n4066) );
  BUFFD0 U4053 ( .I(n4068), .Z(n4067) );
  BUFFD0 U4054 ( .I(n4069), .Z(n4068) );
  BUFFD0 U4055 ( .I(n4070), .Z(n4069) );
  BUFFD0 U4056 ( .I(n4071), .Z(n4070) );
  BUFFD0 U4057 ( .I(n4072), .Z(n4071) );
  BUFFD0 U4058 ( .I(n4073), .Z(n4072) );
  BUFFD0 U4059 ( .I(n4074), .Z(n4073) );
  BUFFD0 U4060 ( .I(n4075), .Z(n4074) );
  BUFFD0 U4061 ( .I(n4076), .Z(n4075) );
  BUFFD0 U4062 ( .I(n4077), .Z(n4076) );
  BUFFD0 U4063 ( .I(n4078), .Z(n4077) );
  BUFFD0 U4064 ( .I(n4079), .Z(n4078) );
  BUFFD0 U4065 ( .I(n4080), .Z(n4079) );
  BUFFD0 U4066 ( .I(n4081), .Z(n4080) );
  BUFFD0 U4067 ( .I(n4082), .Z(n4081) );
  BUFFD0 U4068 ( .I(n4083), .Z(n4082) );
  BUFFD0 U4069 ( .I(n4084), .Z(n4083) );
  BUFFD0 U4070 ( .I(n4085), .Z(n4084) );
  BUFFD0 U4071 ( .I(n4086), .Z(n4085) );
  BUFFD0 U4072 ( .I(n4087), .Z(n4086) );
  BUFFD0 U4073 ( .I(n4088), .Z(n4087) );
  BUFFD0 U4074 ( .I(n4089), .Z(n4088) );
  BUFFD0 U4075 ( .I(n4090), .Z(n4089) );
  BUFFD0 U4076 ( .I(n4091), .Z(n4090) );
  BUFFD0 U4077 ( .I(n4092), .Z(n4091) );
  BUFFD0 U4078 ( .I(n4093), .Z(n4092) );
  BUFFD0 U4079 ( .I(n4094), .Z(n4093) );
  BUFFD0 U4080 ( .I(n4095), .Z(n4094) );
  BUFFD0 U4081 ( .I(n4096), .Z(n4095) );
  BUFFD0 U4082 ( .I(n4097), .Z(n4096) );
  BUFFD0 U4083 ( .I(n4098), .Z(n4097) );
  BUFFD0 U4084 ( .I(n4099), .Z(n4098) );
  BUFFD0 U4085 ( .I(n4100), .Z(n4099) );
  BUFFD0 U4086 ( .I(n4101), .Z(n4100) );
  BUFFD0 U4087 ( .I(n4102), .Z(n4101) );
  BUFFD0 U4088 ( .I(n4103), .Z(n4102) );
  BUFFD0 U4089 ( .I(n4104), .Z(n4103) );
  BUFFD0 U4090 ( .I(n4105), .Z(n4104) );
  BUFFD0 U4091 ( .I(n4106), .Z(n4105) );
  BUFFD0 U4092 ( .I(n4107), .Z(n4106) );
  BUFFD0 U4093 ( .I(n4108), .Z(n4107) );
  BUFFD0 U4094 ( .I(n4109), .Z(n4108) );
  BUFFD0 U4095 ( .I(n4110), .Z(n4109) );
  BUFFD0 U4096 ( .I(n4111), .Z(n4110) );
  BUFFD0 U4097 ( .I(n4112), .Z(n4111) );
  BUFFD0 U4098 ( .I(n4113), .Z(n4112) );
  BUFFD0 U4099 ( .I(n4114), .Z(n4113) );
  BUFFD0 U4100 ( .I(n4115), .Z(n4114) );
  BUFFD0 U4101 ( .I(n4116), .Z(n4115) );
  BUFFD0 U4102 ( .I(n4117), .Z(n4116) );
  BUFFD0 U4103 ( .I(n4118), .Z(n4117) );
  BUFFD0 U4104 ( .I(n4119), .Z(n4118) );
  BUFFD0 U4105 ( .I(n4120), .Z(n4119) );
  BUFFD0 U4106 ( .I(n4121), .Z(n4120) );
  BUFFD0 U4107 ( .I(n4122), .Z(n4121) );
  BUFFD0 U4108 ( .I(n4123), .Z(n4122) );
  BUFFD0 U4109 ( .I(n4124), .Z(n4123) );
  BUFFD0 U4110 ( .I(n4125), .Z(n4124) );
  BUFFD0 U4111 ( .I(n4126), .Z(n4125) );
  BUFFD0 U4112 ( .I(n4127), .Z(n4126) );
  BUFFD0 U4113 ( .I(n4128), .Z(n4127) );
  BUFFD0 U4114 ( .I(n4129), .Z(n4128) );
  BUFFD0 U4115 ( .I(n4130), .Z(n4129) );
  BUFFD0 U4116 ( .I(n4131), .Z(n4130) );
  BUFFD0 U4117 ( .I(N85), .Z(n4131) );
  BUFFD0 U4118 ( .I(n4133), .Z(n4132) );
  BUFFD0 U4119 ( .I(n4134), .Z(n4133) );
  BUFFD0 U4120 ( .I(n4135), .Z(n4134) );
  BUFFD0 U4121 ( .I(n4136), .Z(n4135) );
  BUFFD0 U4122 ( .I(n4137), .Z(n4136) );
  BUFFD0 U4123 ( .I(n4138), .Z(n4137) );
  BUFFD0 U4124 ( .I(n4139), .Z(n4138) );
  BUFFD0 U4125 ( .I(n4140), .Z(n4139) );
  BUFFD0 U4126 ( .I(n4141), .Z(n4140) );
  BUFFD0 U4127 ( .I(n4142), .Z(n4141) );
  BUFFD0 U4128 ( .I(n4143), .Z(n4142) );
  BUFFD0 U4129 ( .I(n4144), .Z(n4143) );
  BUFFD0 U4130 ( .I(n4145), .Z(n4144) );
  BUFFD0 U4131 ( .I(n4146), .Z(n4145) );
  BUFFD0 U4132 ( .I(n4147), .Z(n4146) );
  BUFFD0 U4133 ( .I(n4148), .Z(n4147) );
  BUFFD0 U4134 ( .I(n4149), .Z(n4148) );
  BUFFD0 U4135 ( .I(n4150), .Z(n4149) );
  BUFFD0 U4136 ( .I(n4151), .Z(n4150) );
  BUFFD0 U4137 ( .I(n4152), .Z(n4151) );
  BUFFD0 U4138 ( .I(n4153), .Z(n4152) );
  BUFFD0 U4139 ( .I(n4154), .Z(n4153) );
  BUFFD0 U4140 ( .I(n4155), .Z(n4154) );
  BUFFD0 U4141 ( .I(n4156), .Z(n4155) );
  BUFFD0 U4142 ( .I(n4157), .Z(n4156) );
  BUFFD0 U4143 ( .I(n4158), .Z(n4157) );
  BUFFD0 U4144 ( .I(n4159), .Z(n4158) );
  BUFFD0 U4145 ( .I(n4160), .Z(n4159) );
  BUFFD0 U4146 ( .I(n4161), .Z(n4160) );
  BUFFD0 U4147 ( .I(n4162), .Z(n4161) );
  BUFFD0 U4148 ( .I(n4163), .Z(n4162) );
  BUFFD0 U4149 ( .I(n4164), .Z(n4163) );
  BUFFD0 U4150 ( .I(n4165), .Z(n4164) );
  BUFFD0 U4151 ( .I(n4166), .Z(n4165) );
  BUFFD0 U4152 ( .I(n4167), .Z(n4166) );
  BUFFD0 U4153 ( .I(n4168), .Z(n4167) );
  BUFFD0 U4154 ( .I(n4169), .Z(n4168) );
  BUFFD0 U4155 ( .I(n4170), .Z(n4169) );
  BUFFD0 U4156 ( .I(n4171), .Z(n4170) );
  BUFFD0 U4157 ( .I(n4172), .Z(n4171) );
  BUFFD0 U4158 ( .I(n4173), .Z(n4172) );
  BUFFD0 U4159 ( .I(n4174), .Z(n4173) );
  BUFFD0 U4160 ( .I(n4175), .Z(n4174) );
  BUFFD0 U4161 ( .I(n4176), .Z(n4175) );
  BUFFD0 U4162 ( .I(n4177), .Z(n4176) );
  BUFFD0 U4163 ( .I(n4178), .Z(n4177) );
  BUFFD0 U4164 ( .I(n4179), .Z(n4178) );
  BUFFD0 U4165 ( .I(n4327), .Z(n4179) );
  CKAN2D0 U4166 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U4167 ( .I(N50), .ZN(n4280) );
  BUFFD1 U4168 ( .I(n4342), .Z(n4330) );
  BUFFD1 U4169 ( .I(n4344), .Z(n4331) );
  BUFFD1 U4170 ( .I(n4343), .Z(n4332) );
  BUFFD1 U4171 ( .I(n4339), .Z(n4333) );
  BUFFD1 U4172 ( .I(n4341), .Z(n4334) );
  BUFFD1 U4173 ( .I(n4341), .Z(n4335) );
  BUFFD1 U4174 ( .I(n4340), .Z(n4336) );
  BUFFD1 U4175 ( .I(n4340), .Z(n4337) );
  BUFFD1 U4176 ( .I(n4339), .Z(n4338) );
  BUFFD1 U4177 ( .I(n4343), .Z(n4342) );
  BUFFD1 U4178 ( .I(n4343), .Z(n4341) );
  BUFFD1 U4179 ( .I(n4344), .Z(n4340) );
  BUFFD1 U4180 ( .I(n4344), .Z(n4339) );
  BUFFD1 U4181 ( .I(n4345), .Z(n4343) );
  BUFFD1 U4182 ( .I(n4345), .Z(n4344) );
  INVD1 U4183 ( .I(Reset), .ZN(n4345) );
  BUFFD1 U4184 ( .I(ClockW), .Z(n4314) );
  BUFFD1 U4185 ( .I(n4319), .Z(n4313) );
  BUFFD1 U4186 ( .I(n4314), .Z(n4312) );
  INVD1 U4187 ( .I(n4303), .ZN(n4304) );
  INVD1 U4188 ( .I(n4301), .ZN(n4300) );
  INVD1 U4189 ( .I(n4301), .ZN(n4299) );
  INVD1 U4190 ( .I(n3), .ZN(n4293) );
  INVD1 U4191 ( .I(n3), .ZN(n4292) );
  INVD1 U4192 ( .I(n4291), .ZN(n4290) );
  INVD1 U4193 ( .I(n4291), .ZN(n4289) );
  BUFFD1 U4194 ( .I(n4321), .Z(n4318) );
  BUFFD1 U4195 ( .I(n4321), .Z(n4317) );
  BUFFD1 U4196 ( .I(n4322), .Z(n4316) );
  BUFFD1 U4197 ( .I(n4322), .Z(n4315) );
  BUFFD1 U4198 ( .I(n4320), .Z(n4319) );
  INVD1 U4199 ( .I(N227), .ZN(n4301) );
  INVD1 U4200 ( .I(N359), .ZN(n4291) );
  INVD1 U4201 ( .I(n4309), .ZN(n4308) );
  INVD1 U4202 ( .I(n4309), .ZN(n4307) );
  INVD1 U4203 ( .I(n5), .ZN(n4306) );
  INVD1 U4204 ( .I(n5), .ZN(n4305) );
  INVD1 U4205 ( .I(n6), .ZN(n4298) );
  INVD1 U4206 ( .I(n4294), .ZN(n4296) );
  INVD1 U4207 ( .I(n4294), .ZN(n4295) );
  BUFFD1 U4208 ( .I(n4310), .Z(n4320) );
  BUFFD1 U4209 ( .I(n4310), .Z(n4321) );
  BUFFD1 U4210 ( .I(n4310), .Z(n4322) );
  INVD1 U4211 ( .I(n4), .ZN(n4324) );
  INVD1 U4212 ( .I(n4), .ZN(n4323) );
  XOR3D1 U4213 ( .A1(N69), .A2(N68), .A3(n4354), .Z(n4356) );
  XOR3D1 U4214 ( .A1(N67), .A2(n4353), .A3(n4352), .Z(n4354) );
  XOR3D1 U4215 ( .A1(N62), .A2(N61), .A3(n4351), .Z(n4352) );
  XOR3D1 U4216 ( .A1(n4350), .A2(N60), .A3(n4349), .Z(n4351) );
  XOR3D1 U4217 ( .A1(n4065), .A2(n4064), .A3(n4360), .Z(N85) );
  XOR3D1 U4218 ( .A1(N75), .A2(n4359), .A3(n4358), .Z(n4360) );
  XOR3D1 U4219 ( .A1(N79), .A2(N78), .A3(n4357), .Z(n4358) );
  BUFFD1 U4220 ( .I(n4328), .Z(n4286) );
  BUFFD1 U4221 ( .I(n4328), .Z(n4287) );
  BUFFD1 U4222 ( .I(n4285), .Z(n4288) );
  BUFFD1 U4223 ( .I(n4328), .Z(n4285) );
  BUFFD1 U4224 ( .I(n4329), .Z(n4284) );
  BUFFD1 U4225 ( .I(n4329), .Z(n4283) );
  INVD1 U4226 ( .I(n4280), .ZN(n4281) );
  INVD1 U4227 ( .I(n4280), .ZN(n4282) );
  INVD1 U4228 ( .I(AddrW[0]), .ZN(n4346) );
  INVD1 U4229 ( .I(N99), .ZN(n4309) );
  INVD1 U4230 ( .I(n4303), .ZN(n4302) );
  INVD1 U4231 ( .I(N194), .ZN(n4303) );
  NR3D0 U4232 ( .A1(n4348), .A2(AddrW[0]), .A3(n4373), .ZN(N194) );
  NR3D0 U4233 ( .A1(n4348), .A2(n4373), .A3(n4346), .ZN(N227) );
  NR3D0 U4234 ( .A1(n4348), .A2(n4347), .A3(n4346), .ZN(N359) );
  INVD1 U4235 ( .I(n2), .ZN(n4325) );
  INVD1 U4236 ( .I(n2), .ZN(n4326) );
  BUFFD1 U4237 ( .I(n4311), .Z(n4310) );
  BUFFD1 U4238 ( .I(ClockW), .Z(n4311) );
  XOR3D1 U4239 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n4372), .Z(N87) );
  XOR3D1 U4240 ( .A1(DataI[0]), .A2(n4371), .A3(n4370), .Z(n4372) );
  XOR3D1 U4241 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n4369), .Z(n4370) );
  XOR3D1 U4242 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n4363), .Z(n4364) );
  XOR3D1 U4243 ( .A1(n4362), .A2(DataI[17]), .A3(n4361), .Z(n4363) );
  XOR3D1 U4244 ( .A1(n4368), .A2(DataI[3]), .A3(n4367), .Z(n4369) );
  XOR3D1 U4245 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n4366), .Z(n4367) );
  XOR3D1 U4246 ( .A1(n4365), .A2(DataI[10]), .A3(n4364), .Z(n4366) );
  MUX4ND0 U4247 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n4286), .S1(n4283), .ZN(
        n4261) );
  MUX4ND0 U4248 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n4288), .S1(n4283), .ZN(
        n4264) );
  MUX4ND0 U4249 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n4286), .S1(n4283), .ZN(
        n4258) );
  MUX4ND0 U4250 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n4288), .S1(n4283), .ZN(
        n4267) );
  BUFFD1 U4251 ( .I(N48), .Z(n4328) );
  MUX4ND0 U4252 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n4288), .S1(N49), .ZN(
        n4186) );
  MUX4ND0 U4253 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n4288), .S1(N49), .ZN(
        n4189) );
  MUX4ND0 U4254 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n4288), .S1(n4283), .ZN(
        n4204) );
  MUX4ND0 U4255 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(N48), .S1(n4283), .ZN(
        n4219) );
  MUX4ND0 U4256 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n4286), .S1(n4283), .ZN(
        n4222) );
  MUX4ND0 U4257 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n4286), .S1(n4284), .ZN(
        n4240) );
  MUX4ND0 U4258 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(N48), .S1(N49), .ZN(
        n4243) );
  MUX4ND0 U4259 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n4288), .S1(n4283), .ZN(
        n4273) );
  MUX4ND0 U4260 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n4288), .S1(n4283), .ZN(
        n4276) );
  MUX4ND0 U4261 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n4328), .S1(n4283), .ZN(
        n4201) );
  MUX4ND0 U4262 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n4285), .S1(n4329), .ZN(
        n4207) );
  MUX4ND0 U4263 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(N48), .S1(n4283), .ZN(
        n4231) );
  MUX4ND0 U4264 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n4286), .S1(n4284), .ZN(
        n4252) );
  MUX4ND0 U4265 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n4288), .S1(n4283), .ZN(
        n4255) );
  MUX4ND0 U4266 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n4288), .S1(N49), .ZN(
        n4183) );
  MUX4ND0 U4267 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n4285), .S1(N49), .ZN(
        n4195) );
  MUX4ND0 U4268 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(N48), .S1(n4329), .ZN(
        n4213) );
  MUX4ND0 U4269 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n4285), .S1(n4283), .ZN(
        n4216) );
  MUX4ND0 U4270 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(N48), .S1(n4283), .ZN(
        n4225) );
  MUX4ND0 U4271 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n4286), .S1(n4283), .ZN(
        n4237) );
  MUX4ND0 U4272 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n4286), .S1(n4283), .ZN(
        n4246) );
  MUX4ND0 U4273 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n4288), .S1(n4284), .ZN(
        n4270) );
  MUX4ND0 U4274 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n4288), .S1(N49), .ZN(
        n4192) );
  MUX4ND0 U4275 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n4288), .S1(N49), .ZN(
        n4198) );
  MUX4ND0 U4276 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n4328), .S1(N49), .ZN(
        n4210) );
  MUX4ND0 U4277 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(N48), .S1(n4283), .ZN(
        n4228) );
  MUX4ND0 U4278 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n4286), .S1(n4283), .ZN(
        n4234) );
  MUX4ND0 U4279 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(N48), .S1(n4329), .ZN(
        n4249) );
  MUX4ND0 U4280 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n4288), .S1(n4283), .ZN(
        n4279) );
  BUFFD1 U4281 ( .I(N49), .Z(n4329) );
  INVD1 U4282 ( .I(n6), .ZN(n4297) );
  NR3D0 U4283 ( .A1(n4373), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N99) );
  INVD1 U4284 ( .I(N293), .ZN(n4294) );
  NR3D0 U4285 ( .A1(n4346), .A2(AddrW[1]), .A3(n4347), .ZN(N293) );
  INVD1 U4286 ( .I(AddrW[1]), .ZN(n4348) );
  ND2D1 U4287 ( .A1(AddrW[2]), .A2(Write), .ZN(n4347) );
  IND2D1 U4288 ( .A1(AddrW[2]), .B1(Write), .ZN(n4373) );
  INVD1 U4289 ( .I(Read), .ZN(n4327) );
  CKAN2D0 U4290 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  MUX3ND0 U4291 ( .I0(n4181), .I1(n4182), .I2(n4183), .S0(n4284), .S1(n4281), 
        .ZN(N84) );
  MUX3ND0 U4292 ( .I0(n4184), .I1(n4185), .I2(n4186), .S0(n4284), .S1(n4281), 
        .ZN(N83) );
  MUX3ND0 U4293 ( .I0(n4187), .I1(n4188), .I2(n4189), .S0(n4284), .S1(n4281), 
        .ZN(N82) );
  MUX3ND0 U4294 ( .I0(n4190), .I1(n4191), .I2(n4192), .S0(n4284), .S1(n4281), 
        .ZN(N81) );
  MUX3ND0 U4295 ( .I0(n4193), .I1(n4194), .I2(n4195), .S0(n4284), .S1(n4281), 
        .ZN(N80) );
  MUX3ND0 U4296 ( .I0(n4196), .I1(n4197), .I2(n4198), .S0(n4284), .S1(n4281), 
        .ZN(N79) );
  MUX3ND0 U4297 ( .I0(n4199), .I1(n4200), .I2(n4201), .S0(n4284), .S1(n4281), 
        .ZN(N78) );
  MUX3ND0 U4298 ( .I0(n4202), .I1(n4203), .I2(n4204), .S0(n4284), .S1(n4281), 
        .ZN(N77) );
  MUX3ND0 U4299 ( .I0(n4205), .I1(n4206), .I2(n4207), .S0(n4284), .S1(n4281), 
        .ZN(N76) );
  MUX3ND0 U4300 ( .I0(n4208), .I1(n4209), .I2(n4210), .S0(n4284), .S1(n4281), 
        .ZN(N75) );
  MUX3ND0 U4301 ( .I0(n4211), .I1(n4212), .I2(n4213), .S0(n4284), .S1(n4281), 
        .ZN(N74) );
  MUX3ND0 U4302 ( .I0(n4214), .I1(n4215), .I2(n4216), .S0(n4284), .S1(n4281), 
        .ZN(N73) );
  MUX3ND0 U4303 ( .I0(n4217), .I1(n4218), .I2(n4219), .S0(n4284), .S1(n4281), 
        .ZN(N72) );
  MUX3ND0 U4304 ( .I0(n4220), .I1(n4221), .I2(n4222), .S0(n4329), .S1(n4281), 
        .ZN(N71) );
  MUX3ND0 U4305 ( .I0(n4223), .I1(n4224), .I2(n4225), .S0(n4329), .S1(n4281), 
        .ZN(N70) );
  MUX3ND0 U4306 ( .I0(n4226), .I1(n4227), .I2(n4228), .S0(n4329), .S1(n4281), 
        .ZN(N69) );
  MUX3ND0 U4307 ( .I0(n4229), .I1(n4230), .I2(n4231), .S0(n4329), .S1(n4281), 
        .ZN(N68) );
  MUX3ND0 U4308 ( .I0(n4232), .I1(n4233), .I2(n4234), .S0(n4329), .S1(n4281), 
        .ZN(N67) );
  MUX3ND0 U4309 ( .I0(n4235), .I1(n4236), .I2(n4237), .S0(n4329), .S1(n4281), 
        .ZN(N66) );
  MUX3ND0 U4310 ( .I0(n4238), .I1(n4239), .I2(n4240), .S0(n4329), .S1(n4281), 
        .ZN(N65) );
  MUX3ND0 U4311 ( .I0(n4241), .I1(n4242), .I2(n4243), .S0(n4329), .S1(n4282), 
        .ZN(N64) );
  MUX3ND0 U4312 ( .I0(n4244), .I1(n4245), .I2(n4246), .S0(n4329), .S1(n4282), 
        .ZN(N63) );
  MUX3ND0 U4313 ( .I0(n4247), .I1(n4248), .I2(n4249), .S0(n4329), .S1(n4282), 
        .ZN(N62) );
  MUX3ND0 U4314 ( .I0(n4250), .I1(n4251), .I2(n4252), .S0(n4329), .S1(n4282), 
        .ZN(N61) );
  MUX3ND0 U4315 ( .I0(n4253), .I1(n4254), .I2(n4255), .S0(n4329), .S1(n4282), 
        .ZN(N60) );
  MUX3ND0 U4316 ( .I0(n4256), .I1(n4257), .I2(n4258), .S0(n4284), .S1(n4282), 
        .ZN(N59) );
  MUX3ND0 U4317 ( .I0(n4259), .I1(n4260), .I2(n4261), .S0(n4284), .S1(n4282), 
        .ZN(N58) );
  MUX3ND0 U4318 ( .I0(n4262), .I1(n4263), .I2(n4264), .S0(n4284), .S1(n4282), 
        .ZN(N57) );
  MUX3ND0 U4319 ( .I0(n4265), .I1(n4266), .I2(n4267), .S0(n4329), .S1(n4282), 
        .ZN(N56) );
  MUX3ND0 U4320 ( .I0(n4268), .I1(n4269), .I2(n4270), .S0(N49), .S1(n4282), 
        .ZN(N55) );
  MUX3ND0 U4321 ( .I0(n4271), .I1(n4272), .I2(n4273), .S0(N49), .S1(n4282), 
        .ZN(N54) );
  MUX3ND0 U4322 ( .I0(n4274), .I1(n4275), .I2(n4276), .S0(N49), .S1(n4282), 
        .ZN(N53) );
  MUX3ND0 U4323 ( .I0(n4277), .I1(n4278), .I2(n4279), .S0(N49), .S1(n4282), 
        .ZN(N52) );
  MUX2ND0 U4324 ( .I0(\Storage[2][0] ), .I1(\Storage[3][0] ), .S(n4285), .ZN(
        n4182) );
  MUX2ND0 U4325 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .S(n4285), .ZN(
        n4181) );
  MUX2ND0 U4326 ( .I0(\Storage[2][1] ), .I1(\Storage[3][1] ), .S(N48), .ZN(
        n4185) );
  MUX2ND0 U4327 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .S(n4328), .ZN(
        n4184) );
  MUX2ND0 U4328 ( .I0(\Storage[2][2] ), .I1(\Storage[3][2] ), .S(n4328), .ZN(
        n4188) );
  MUX2ND0 U4329 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .S(n4286), .ZN(
        n4187) );
  MUX2ND0 U4330 ( .I0(\Storage[2][3] ), .I1(\Storage[3][3] ), .S(n4328), .ZN(
        n4191) );
  MUX2ND0 U4331 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .S(n4328), .ZN(
        n4190) );
  MUX2ND0 U4332 ( .I0(\Storage[2][4] ), .I1(\Storage[3][4] ), .S(n4286), .ZN(
        n4194) );
  MUX2ND0 U4333 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .S(n4328), .ZN(
        n4193) );
  MUX2ND0 U4334 ( .I0(\Storage[2][5] ), .I1(\Storage[3][5] ), .S(n4286), .ZN(
        n4197) );
  MUX2ND0 U4335 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .S(n4285), .ZN(
        n4196) );
  MUX2ND0 U4336 ( .I0(\Storage[2][6] ), .I1(\Storage[3][6] ), .S(n4328), .ZN(
        n4200) );
  MUX2ND0 U4337 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .S(n4286), .ZN(
        n4199) );
  MUX2ND0 U4338 ( .I0(\Storage[2][7] ), .I1(\Storage[3][7] ), .S(n4328), .ZN(
        n4203) );
  MUX2ND0 U4339 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .S(n4328), .ZN(
        n4202) );
  MUX2ND0 U4340 ( .I0(\Storage[2][8] ), .I1(\Storage[3][8] ), .S(n4286), .ZN(
        n4206) );
  MUX2ND0 U4341 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .S(n4286), .ZN(
        n4205) );
  MUX2ND0 U4342 ( .I0(\Storage[2][9] ), .I1(\Storage[3][9] ), .S(n4285), .ZN(
        n4209) );
  MUX2ND0 U4343 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .S(n4285), .ZN(
        n4208) );
  MUX2ND0 U4344 ( .I0(\Storage[2][10] ), .I1(\Storage[3][10] ), .S(n4328), 
        .ZN(n4212) );
  MUX2ND0 U4345 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .S(n4328), 
        .ZN(n4211) );
  MUX2ND0 U4346 ( .I0(\Storage[2][11] ), .I1(\Storage[3][11] ), .S(n4328), 
        .ZN(n4215) );
  MUX2ND0 U4347 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .S(n4285), 
        .ZN(n4214) );
  MUX2ND0 U4348 ( .I0(\Storage[2][12] ), .I1(\Storage[3][12] ), .S(n4328), 
        .ZN(n4218) );
  MUX2ND0 U4349 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .S(n4286), 
        .ZN(n4217) );
  MUX2ND0 U4350 ( .I0(\Storage[2][13] ), .I1(\Storage[3][13] ), .S(n4287), 
        .ZN(n4221) );
  MUX2ND0 U4351 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .S(n4285), 
        .ZN(n4220) );
  MUX2ND0 U4352 ( .I0(\Storage[2][14] ), .I1(\Storage[3][14] ), .S(n4328), 
        .ZN(n4224) );
  MUX2ND0 U4353 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .S(n4285), 
        .ZN(n4223) );
  MUX2ND0 U4354 ( .I0(\Storage[2][15] ), .I1(\Storage[3][15] ), .S(N48), .ZN(
        n4227) );
  MUX2ND0 U4355 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .S(N48), .ZN(
        n4226) );
  MUX2ND0 U4356 ( .I0(\Storage[2][16] ), .I1(\Storage[3][16] ), .S(N48), .ZN(
        n4230) );
  MUX2ND0 U4357 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .S(n4328), 
        .ZN(n4229) );
  MUX2ND0 U4358 ( .I0(\Storage[2][17] ), .I1(\Storage[3][17] ), .S(n4286), 
        .ZN(n4233) );
  MUX2ND0 U4359 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .S(n4285), 
        .ZN(n4232) );
  MUX2ND0 U4360 ( .I0(\Storage[2][18] ), .I1(\Storage[3][18] ), .S(n4286), 
        .ZN(n4236) );
  MUX2ND0 U4361 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .S(n4285), 
        .ZN(n4235) );
  MUX2ND0 U4362 ( .I0(\Storage[2][19] ), .I1(\Storage[3][19] ), .S(N48), .ZN(
        n4239) );
  MUX2ND0 U4363 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .S(n4285), 
        .ZN(n4238) );
  MUX2ND0 U4364 ( .I0(\Storage[2][20] ), .I1(\Storage[3][20] ), .S(n4285), 
        .ZN(n4242) );
  MUX2ND0 U4365 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .S(N48), .ZN(
        n4241) );
  MUX2ND0 U4366 ( .I0(\Storage[2][21] ), .I1(\Storage[3][21] ), .S(N48), .ZN(
        n4245) );
  MUX2ND0 U4367 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .S(n4287), 
        .ZN(n4244) );
  MUX2ND0 U4368 ( .I0(\Storage[2][22] ), .I1(\Storage[3][22] ), .S(n4286), 
        .ZN(n4248) );
  MUX2ND0 U4369 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .S(n4287), 
        .ZN(n4247) );
  MUX2ND0 U4370 ( .I0(\Storage[2][23] ), .I1(\Storage[3][23] ), .S(n4287), 
        .ZN(n4251) );
  MUX2ND0 U4371 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .S(n4287), 
        .ZN(n4250) );
  MUX2ND0 U4372 ( .I0(\Storage[2][24] ), .I1(\Storage[3][24] ), .S(n4287), 
        .ZN(n4254) );
  MUX2ND0 U4373 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .S(n4287), 
        .ZN(n4253) );
  MUX2ND0 U4374 ( .I0(\Storage[2][25] ), .I1(\Storage[3][25] ), .S(n4287), 
        .ZN(n4257) );
  MUX2ND0 U4375 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .S(n4287), 
        .ZN(n4256) );
  MUX2ND0 U4376 ( .I0(\Storage[2][26] ), .I1(\Storage[3][26] ), .S(n4287), 
        .ZN(n4260) );
  MUX2ND0 U4377 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .S(n4287), 
        .ZN(n4259) );
  MUX2ND0 U4378 ( .I0(\Storage[2][27] ), .I1(\Storage[3][27] ), .S(n4287), 
        .ZN(n4263) );
  MUX2ND0 U4379 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .S(n4287), 
        .ZN(n4262) );
  MUX2ND0 U4380 ( .I0(\Storage[2][28] ), .I1(\Storage[3][28] ), .S(n4287), 
        .ZN(n4266) );
  MUX2ND0 U4381 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .S(n4287), 
        .ZN(n4265) );
  MUX2ND0 U4382 ( .I0(\Storage[2][29] ), .I1(\Storage[3][29] ), .S(n4287), 
        .ZN(n4269) );
  MUX2ND0 U4383 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .S(n4287), 
        .ZN(n4268) );
  MUX2ND0 U4384 ( .I0(\Storage[2][30] ), .I1(\Storage[3][30] ), .S(n4287), 
        .ZN(n4272) );
  MUX2ND0 U4385 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .S(n4287), 
        .ZN(n4271) );
  MUX2ND0 U4386 ( .I0(\Storage[2][31] ), .I1(\Storage[3][31] ), .S(n4287), 
        .ZN(n4275) );
  MUX2ND0 U4387 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .S(n4286), 
        .ZN(n4274) );
  MUX2ND0 U4388 ( .I0(\Storage[2][32] ), .I1(\Storage[3][32] ), .S(n4286), 
        .ZN(n4278) );
  MUX2ND0 U4389 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .S(n4328), 
        .ZN(n4277) );
endmodule


module PLLTop_1 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_1 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_1 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_1 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module PLLTop_2 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_2 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_2 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_2 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module PLLTop_3 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_3 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_3 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_3 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module FIFOStateM_AWid4_1 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [3:0] ReadAddr;
  output [3:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n1799, n1800, n1801, StateClockRaw, StateClock, N47, N48, N49, N50,
         N51, N67, N68, N69, N70, N71, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n69, n88, n89, n93,
         n133, n134, n135, n136, n137, n138, n139, n140, n142, n145, n146,
         n161, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1746, n1747, n1748, n1749,
         n1750, n1751, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798;
  wire   [2:0] NextState;
  wire   [3:0] OldReadAr;
  wire   [3:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n191), .CPN(StateClock), .Q(n1799) );
  DFND1 EmptyFIFOr_reg ( .D(n6), .CPN(StateClock), .Q(EmptyFIFO), .QN(n1705)
         );
  OA21D1 U11 ( .A1(n1677), .A2(n1679), .B(n1798), .Z(n1789) );
  IAO21D1 U31 ( .A1(n1761), .A2(n1760), .B(n1778), .ZN(n1762) );
  OA21D1 U34 ( .A1(ReadAddr[2]), .A2(n1758), .B(n1759), .Z(n1753) );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n252), .CPN(StateClock), .CDN(n1675), .QN(
        n1792) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n310), .CPN(StateClock), .CDN(n1675), .QN(
        n1794) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n368), .CPN(StateClock), .CDN(n1674), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n426), .CPN(StateClock), .CDN(n1674), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n488), .CPN(StateClock), .CDN(n1675), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n550), .CPN(StateClock), .CDN(n1675), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n611), .CPN(StateClock), .CDN(n1675), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n672), .CPN(StateClock), .CDN(n1675), .Q(
        OldReadAr[1]) );
  DFNCND1 \NextState_reg[0]  ( .D(n786), .CPN(StateClock), .CDN(n1674), .Q(
        NextState[0]), .QN(n1702) );
  DFNCND1 \NextState_reg[1]  ( .D(n848), .CPN(StateClock), .CDN(n1674), .Q(
        NextState[1]), .QN(n1703) );
  DFNCND1 \NextState_reg[2]  ( .D(n910), .CPN(StateClock), .CDN(n1674), .Q(
        NextState[2]), .QN(n1704) );
  DFNCND1 WriteCmdr_reg ( .D(n976), .CPN(StateClock), .CDN(n1674), .Q(n1801)
         );
  DFNCND1 ReadCmdr_reg ( .D(n1036), .CPN(StateClock), .CDN(n1674), .Q(n1800)
         );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n1674), 
        .QN(n1679) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n1674), 
        .Q(n1781), .QN(n1677) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n1674), 
        .Q(n5), .QN(n1678) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(n1105), .E(n3), .CP(StateClock), .CDN(n1675), 
        .Q(WriteAddr[1]) );
  EDFCND1 \ReadAr_reg[3]  ( .D(n1167), .E(n1387), .CP(StateClock), .CDN(n1674), 
        .Q(ReadAddr[3]), .QN(n1686) );
  EDFCND1 \ReadAr_reg[2]  ( .D(n1221), .E(n1387), .CP(StateClock), .CDN(n1675), 
        .Q(ReadAddr[2]), .QN(n1685) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n1279), .E(n1387), .CP(StateClock), .CDN(n1675), 
        .Q(ReadAddr[1]), .QN(n1684) );
  EDFCND1 \ReadAr_reg[0]  ( .D(n1333), .E(n1387), .CP(StateClock), .CDN(n1675), 
        .Q(ReadAddr[0]), .QN(n1683) );
  EDFCND1 \WriteAr_reg[3]  ( .D(n1434), .E(n3), .CP(StateClock), .CDN(n1675), 
        .Q(WriteAddr[3]), .QN(n1682) );
  EDFCND1 \WriteAr_reg[2]  ( .D(n1494), .E(n3), .CP(StateClock), .CDN(n1674), 
        .Q(WriteAddr[2]), .QN(n1681) );
  EDFCND1 \WriteAr_reg[0]  ( .D(n1554), .E(n3), .CP(StateClock), .CDN(n1675), 
        .Q(WriteAddr[0]), .QN(n1680) );
  CKBD0 U3 ( .CLK(n1798), .C(n1416) );
  BUFFD0 U4 ( .I(n1664), .Z(n1) );
  BUFFD0 U5 ( .I(n1), .Z(n2) );
  BUFFD0 U6 ( .I(n1616), .Z(n3) );
  AN3D1 U7 ( .A1(n1791), .A2(n1664), .A3(n1777), .Z(n4) );
  INVD1 U8 ( .I(n4), .ZN(N71) );
  BUFFD0 U9 ( .I(n8), .Z(n6) );
  BUFFD0 U10 ( .I(n1701), .Z(n7) );
  BUFFD0 U12 ( .I(n9), .Z(n8) );
  BUFFD0 U13 ( .I(n10), .Z(n9) );
  BUFFD0 U14 ( .I(n14), .Z(n10) );
  BUFFD0 U15 ( .I(n12), .Z(n11) );
  BUFFD0 U16 ( .I(n13), .Z(n12) );
  BUFFD0 U17 ( .I(n1705), .Z(n13) );
  BUFFD0 U18 ( .I(n15), .Z(n14) );
  BUFFD0 U19 ( .I(n16), .Z(n15) );
  BUFFD0 U20 ( .I(n17), .Z(n16) );
  BUFFD0 U21 ( .I(n18), .Z(n17) );
  BUFFD0 U22 ( .I(n19), .Z(n18) );
  BUFFD0 U23 ( .I(n20), .Z(n19) );
  BUFFD0 U24 ( .I(n21), .Z(n20) );
  BUFFD0 U25 ( .I(n22), .Z(n21) );
  BUFFD0 U26 ( .I(n23), .Z(n22) );
  BUFFD0 U27 ( .I(n24), .Z(n23) );
  BUFFD0 U28 ( .I(n25), .Z(n24) );
  BUFFD0 U29 ( .I(n26), .Z(n25) );
  BUFFD0 U30 ( .I(n27), .Z(n26) );
  BUFFD0 U32 ( .I(n28), .Z(n27) );
  BUFFD0 U33 ( .I(n29), .Z(n28) );
  BUFFD0 U35 ( .I(n30), .Z(n29) );
  BUFFD0 U36 ( .I(n31), .Z(n30) );
  BUFFD0 U37 ( .I(n32), .Z(n31) );
  BUFFD0 U38 ( .I(n33), .Z(n32) );
  BUFFD0 U39 ( .I(n34), .Z(n33) );
  BUFFD0 U40 ( .I(n69), .Z(n34) );
  BUFFD0 U41 ( .I(n88), .Z(n69) );
  BUFFD0 U42 ( .I(n89), .Z(n88) );
  BUFFD0 U43 ( .I(n93), .Z(n89) );
  BUFFD0 U44 ( .I(n133), .Z(n93) );
  BUFFD0 U45 ( .I(n134), .Z(n133) );
  BUFFD0 U46 ( .I(n135), .Z(n134) );
  BUFFD0 U47 ( .I(n136), .Z(n135) );
  BUFFD0 U48 ( .I(n137), .Z(n136) );
  BUFFD0 U49 ( .I(n138), .Z(n137) );
  BUFFD0 U50 ( .I(n139), .Z(n138) );
  BUFFD0 U51 ( .I(n140), .Z(n139) );
  BUFFD0 U52 ( .I(n142), .Z(n140) );
  BUFFD0 U53 ( .I(n145), .Z(n142) );
  BUFFD0 U54 ( .I(n146), .Z(n145) );
  BUFFD0 U55 ( .I(n161), .Z(n146) );
  BUFFD0 U56 ( .I(n173), .Z(n161) );
  BUFFD0 U57 ( .I(n174), .Z(n173) );
  BUFFD0 U58 ( .I(n175), .Z(n174) );
  BUFFD0 U59 ( .I(n176), .Z(n175) );
  BUFFD0 U60 ( .I(n177), .Z(n176) );
  BUFFD0 U61 ( .I(n178), .Z(n177) );
  BUFFD0 U62 ( .I(n179), .Z(n178) );
  BUFFD0 U63 ( .I(n180), .Z(n179) );
  BUFFD0 U64 ( .I(n181), .Z(n180) );
  BUFFD0 U65 ( .I(n182), .Z(n181) );
  BUFFD0 U66 ( .I(n183), .Z(n182) );
  BUFFD0 U67 ( .I(n184), .Z(n183) );
  BUFFD0 U68 ( .I(n185), .Z(n184) );
  BUFFD0 U69 ( .I(n186), .Z(n185) );
  BUFFD0 U70 ( .I(n187), .Z(n186) );
  BUFFD0 U71 ( .I(n188), .Z(n187) );
  BUFFD0 U72 ( .I(n189), .Z(n188) );
  BUFFD0 U73 ( .I(n190), .Z(n189) );
  BUFFD0 U74 ( .I(n7), .Z(n190) );
  BUFFD0 U75 ( .I(n217), .Z(n191) );
  BUFFD0 U76 ( .I(n193), .Z(n192) );
  BUFFD0 U77 ( .I(n194), .Z(n193) );
  BUFFD0 U78 ( .I(n195), .Z(n194) );
  BUFFD0 U79 ( .I(n196), .Z(n195) );
  BUFFD0 U80 ( .I(n197), .Z(n196) );
  BUFFD0 U81 ( .I(n198), .Z(n197) );
  BUFFD0 U82 ( .I(n199), .Z(n198) );
  BUFFD0 U83 ( .I(n200), .Z(n199) );
  BUFFD0 U84 ( .I(n201), .Z(n200) );
  BUFFD0 U85 ( .I(n202), .Z(n201) );
  BUFFD0 U86 ( .I(n203), .Z(n202) );
  BUFFD0 U87 ( .I(n204), .Z(n203) );
  BUFFD0 U88 ( .I(n205), .Z(n204) );
  BUFFD0 U89 ( .I(n206), .Z(n205) );
  BUFFD0 U90 ( .I(n207), .Z(n206) );
  BUFFD0 U91 ( .I(n208), .Z(n207) );
  BUFFD0 U92 ( .I(n209), .Z(n208) );
  BUFFD0 U93 ( .I(n210), .Z(n209) );
  BUFFD0 U94 ( .I(n211), .Z(n210) );
  BUFFD0 U95 ( .I(n212), .Z(n211) );
  BUFFD0 U96 ( .I(n213), .Z(n212) );
  BUFFD0 U97 ( .I(n214), .Z(n213) );
  BUFFD0 U98 ( .I(n215), .Z(n214) );
  BUFFD0 U99 ( .I(n225), .Z(n215) );
  BUFFD0 U100 ( .I(n1799), .Z(FullFIFO) );
  BUFFD0 U101 ( .I(n218), .Z(n217) );
  BUFFD0 U102 ( .I(n219), .Z(n218) );
  BUFFD0 U103 ( .I(n220), .Z(n219) );
  BUFFD0 U104 ( .I(n221), .Z(n220) );
  BUFFD0 U105 ( .I(n222), .Z(n221) );
  BUFFD0 U106 ( .I(n223), .Z(n222) );
  BUFFD0 U107 ( .I(n224), .Z(n223) );
  BUFFD0 U108 ( .I(n226), .Z(n224) );
  BUFFD0 U109 ( .I(n1790), .Z(n225) );
  BUFFD0 U110 ( .I(n227), .Z(n226) );
  BUFFD0 U111 ( .I(n228), .Z(n227) );
  BUFFD0 U112 ( .I(n229), .Z(n228) );
  BUFFD0 U113 ( .I(n230), .Z(n229) );
  BUFFD0 U114 ( .I(n231), .Z(n230) );
  BUFFD0 U115 ( .I(n232), .Z(n231) );
  BUFFD0 U116 ( .I(n233), .Z(n232) );
  BUFFD0 U117 ( .I(n234), .Z(n233) );
  BUFFD0 U118 ( .I(n235), .Z(n234) );
  BUFFD0 U119 ( .I(n236), .Z(n235) );
  BUFFD0 U120 ( .I(n237), .Z(n236) );
  BUFFD0 U121 ( .I(n238), .Z(n237) );
  BUFFD0 U122 ( .I(n239), .Z(n238) );
  BUFFD0 U123 ( .I(n240), .Z(n239) );
  BUFFD0 U124 ( .I(n241), .Z(n240) );
  BUFFD0 U125 ( .I(n242), .Z(n241) );
  BUFFD0 U126 ( .I(n243), .Z(n242) );
  BUFFD0 U127 ( .I(n244), .Z(n243) );
  BUFFD0 U128 ( .I(n245), .Z(n244) );
  BUFFD0 U129 ( .I(n246), .Z(n245) );
  BUFFD0 U130 ( .I(n247), .Z(n246) );
  BUFFD0 U131 ( .I(n248), .Z(n247) );
  BUFFD0 U132 ( .I(n249), .Z(n248) );
  BUFFD0 U133 ( .I(n250), .Z(n249) );
  BUFFD0 U134 ( .I(n1697), .Z(n250) );
  CKBD0 U135 ( .CLK(n1801), .C(n251) );
  BUFFD0 U136 ( .I(n254), .Z(n252) );
  BUFFD0 U137 ( .I(n1792), .Z(n253) );
  BUFFD0 U138 ( .I(n256), .Z(n254) );
  BUFFD0 U139 ( .I(n253), .Z(n255) );
  BUFFD0 U140 ( .I(n258), .Z(n256) );
  BUFFD0 U141 ( .I(n255), .Z(n257) );
  BUFFD0 U142 ( .I(n260), .Z(n258) );
  BUFFD0 U143 ( .I(n257), .Z(n259) );
  BUFFD0 U144 ( .I(n262), .Z(n260) );
  BUFFD0 U145 ( .I(n259), .Z(n261) );
  BUFFD0 U146 ( .I(n264), .Z(n262) );
  BUFFD0 U147 ( .I(n261), .Z(n263) );
  BUFFD0 U148 ( .I(n266), .Z(n264) );
  BUFFD0 U149 ( .I(n263), .Z(n265) );
  BUFFD0 U150 ( .I(n268), .Z(n266) );
  BUFFD0 U151 ( .I(n265), .Z(n267) );
  BUFFD0 U152 ( .I(n270), .Z(n268) );
  BUFFD0 U153 ( .I(n267), .Z(n269) );
  BUFFD0 U154 ( .I(n272), .Z(n270) );
  BUFFD0 U155 ( .I(n269), .Z(n271) );
  BUFFD0 U156 ( .I(n274), .Z(n272) );
  BUFFD0 U157 ( .I(n271), .Z(n273) );
  BUFFD0 U158 ( .I(n276), .Z(n274) );
  BUFFD0 U159 ( .I(n273), .Z(n275) );
  BUFFD0 U160 ( .I(n278), .Z(n276) );
  BUFFD0 U161 ( .I(n275), .Z(n277) );
  BUFFD0 U162 ( .I(n280), .Z(n278) );
  BUFFD0 U163 ( .I(n277), .Z(n279) );
  BUFFD0 U164 ( .I(n282), .Z(n280) );
  BUFFD0 U165 ( .I(n279), .Z(n281) );
  BUFFD0 U166 ( .I(n284), .Z(n282) );
  BUFFD0 U167 ( .I(n281), .Z(n283) );
  BUFFD0 U168 ( .I(n286), .Z(n284) );
  BUFFD0 U169 ( .I(n283), .Z(n285) );
  BUFFD0 U170 ( .I(n288), .Z(n286) );
  BUFFD0 U171 ( .I(n285), .Z(n287) );
  BUFFD0 U172 ( .I(n290), .Z(n288) );
  BUFFD0 U173 ( .I(n287), .Z(n289) );
  BUFFD0 U174 ( .I(n292), .Z(n290) );
  BUFFD0 U175 ( .I(n289), .Z(n291) );
  BUFFD0 U176 ( .I(n294), .Z(n292) );
  BUFFD0 U177 ( .I(n291), .Z(n293) );
  BUFFD0 U178 ( .I(n296), .Z(n294) );
  BUFFD0 U179 ( .I(n293), .Z(n295) );
  BUFFD0 U180 ( .I(n298), .Z(n296) );
  BUFFD0 U181 ( .I(n295), .Z(n297) );
  BUFFD0 U182 ( .I(n300), .Z(n298) );
  BUFFD0 U183 ( .I(n297), .Z(n299) );
  BUFFD0 U184 ( .I(n302), .Z(n300) );
  BUFFD0 U185 ( .I(n299), .Z(n301) );
  BUFFD0 U186 ( .I(n304), .Z(n302) );
  BUFFD0 U187 ( .I(n301), .Z(n303) );
  BUFFD0 U188 ( .I(n306), .Z(n304) );
  BUFFD0 U189 ( .I(n303), .Z(n305) );
  BUFFD0 U190 ( .I(n308), .Z(n306) );
  BUFFD0 U191 ( .I(n305), .Z(n307) );
  BUFFD0 U192 ( .I(n309), .Z(n308) );
  BUFFD0 U193 ( .I(n1698), .Z(n309) );
  BUFFD0 U194 ( .I(n312), .Z(n310) );
  BUFFD0 U195 ( .I(n1794), .Z(n311) );
  BUFFD0 U196 ( .I(n314), .Z(n312) );
  BUFFD0 U197 ( .I(n311), .Z(n313) );
  BUFFD0 U198 ( .I(n316), .Z(n314) );
  BUFFD0 U199 ( .I(n313), .Z(n315) );
  BUFFD0 U200 ( .I(n318), .Z(n316) );
  BUFFD0 U201 ( .I(n315), .Z(n317) );
  BUFFD0 U202 ( .I(n320), .Z(n318) );
  BUFFD0 U203 ( .I(n317), .Z(n319) );
  BUFFD0 U204 ( .I(n322), .Z(n320) );
  BUFFD0 U205 ( .I(n319), .Z(n321) );
  BUFFD0 U206 ( .I(n324), .Z(n322) );
  BUFFD0 U207 ( .I(n321), .Z(n323) );
  BUFFD0 U208 ( .I(n326), .Z(n324) );
  BUFFD0 U209 ( .I(n323), .Z(n325) );
  BUFFD0 U210 ( .I(n328), .Z(n326) );
  BUFFD0 U211 ( .I(n325), .Z(n327) );
  BUFFD0 U212 ( .I(n330), .Z(n328) );
  BUFFD0 U213 ( .I(n327), .Z(n329) );
  BUFFD0 U214 ( .I(n332), .Z(n330) );
  BUFFD0 U215 ( .I(n329), .Z(n331) );
  BUFFD0 U216 ( .I(n334), .Z(n332) );
  BUFFD0 U217 ( .I(n331), .Z(n333) );
  BUFFD0 U218 ( .I(n336), .Z(n334) );
  BUFFD0 U219 ( .I(n333), .Z(n335) );
  BUFFD0 U220 ( .I(n338), .Z(n336) );
  BUFFD0 U221 ( .I(n335), .Z(n337) );
  BUFFD0 U222 ( .I(n340), .Z(n338) );
  BUFFD0 U223 ( .I(n337), .Z(n339) );
  BUFFD0 U224 ( .I(n342), .Z(n340) );
  BUFFD0 U225 ( .I(n339), .Z(n341) );
  BUFFD0 U226 ( .I(n344), .Z(n342) );
  BUFFD0 U227 ( .I(n341), .Z(n343) );
  BUFFD0 U228 ( .I(n346), .Z(n344) );
  BUFFD0 U229 ( .I(n343), .Z(n345) );
  BUFFD0 U230 ( .I(n348), .Z(n346) );
  BUFFD0 U231 ( .I(n345), .Z(n347) );
  BUFFD0 U232 ( .I(n350), .Z(n348) );
  BUFFD0 U233 ( .I(n347), .Z(n349) );
  BUFFD0 U234 ( .I(n352), .Z(n350) );
  BUFFD0 U235 ( .I(n349), .Z(n351) );
  BUFFD0 U236 ( .I(n354), .Z(n352) );
  BUFFD0 U237 ( .I(n351), .Z(n353) );
  BUFFD0 U238 ( .I(n356), .Z(n354) );
  BUFFD0 U239 ( .I(n353), .Z(n355) );
  BUFFD0 U240 ( .I(n358), .Z(n356) );
  BUFFD0 U241 ( .I(n355), .Z(n357) );
  BUFFD0 U242 ( .I(n360), .Z(n358) );
  BUFFD0 U243 ( .I(n357), .Z(n359) );
  BUFFD0 U244 ( .I(n362), .Z(n360) );
  BUFFD0 U245 ( .I(n359), .Z(n361) );
  BUFFD0 U246 ( .I(n364), .Z(n362) );
  BUFFD0 U247 ( .I(n361), .Z(n363) );
  BUFFD0 U248 ( .I(n366), .Z(n364) );
  BUFFD0 U249 ( .I(n363), .Z(n365) );
  BUFFD0 U250 ( .I(n367), .Z(n366) );
  BUFFD0 U251 ( .I(n1700), .Z(n367) );
  MOAI22D0 U252 ( .A1(n1683), .A2(n1793), .B1(n1793), .B2(n371), .ZN(n1687) );
  BUFFD0 U253 ( .I(n369), .Z(n368) );
  BUFFD0 U254 ( .I(n370), .Z(n369) );
  BUFFD0 U255 ( .I(n372), .Z(n370) );
  BUFFD0 U256 ( .I(n421), .Z(n371) );
  BUFFD0 U257 ( .I(n373), .Z(n372) );
  BUFFD0 U258 ( .I(n374), .Z(n373) );
  BUFFD0 U259 ( .I(n375), .Z(n374) );
  BUFFD0 U260 ( .I(n376), .Z(n375) );
  BUFFD0 U261 ( .I(n377), .Z(n376) );
  BUFFD0 U262 ( .I(n378), .Z(n377) );
  BUFFD0 U263 ( .I(n379), .Z(n378) );
  BUFFD0 U264 ( .I(n380), .Z(n379) );
  BUFFD0 U265 ( .I(n381), .Z(n380) );
  BUFFD0 U266 ( .I(n382), .Z(n381) );
  BUFFD0 U267 ( .I(n383), .Z(n382) );
  BUFFD0 U268 ( .I(n384), .Z(n383) );
  BUFFD0 U269 ( .I(n385), .Z(n384) );
  BUFFD0 U270 ( .I(n386), .Z(n385) );
  BUFFD0 U271 ( .I(n387), .Z(n386) );
  BUFFD0 U272 ( .I(n388), .Z(n387) );
  BUFFD0 U273 ( .I(n389), .Z(n388) );
  BUFFD0 U274 ( .I(n390), .Z(n389) );
  BUFFD0 U275 ( .I(n391), .Z(n390) );
  BUFFD0 U276 ( .I(n392), .Z(n391) );
  BUFFD0 U277 ( .I(n393), .Z(n392) );
  BUFFD0 U278 ( .I(n394), .Z(n393) );
  BUFFD0 U279 ( .I(n395), .Z(n394) );
  BUFFD0 U280 ( .I(n396), .Z(n395) );
  BUFFD0 U281 ( .I(n397), .Z(n396) );
  BUFFD0 U282 ( .I(n398), .Z(n397) );
  BUFFD0 U283 ( .I(n399), .Z(n398) );
  BUFFD0 U284 ( .I(n400), .Z(n399) );
  BUFFD0 U285 ( .I(n401), .Z(n400) );
  BUFFD0 U286 ( .I(n402), .Z(n401) );
  BUFFD0 U287 ( .I(n403), .Z(n402) );
  BUFFD0 U288 ( .I(n404), .Z(n403) );
  BUFFD0 U289 ( .I(n405), .Z(n404) );
  BUFFD0 U290 ( .I(n406), .Z(n405) );
  BUFFD0 U291 ( .I(n407), .Z(n406) );
  BUFFD0 U292 ( .I(n408), .Z(n407) );
  BUFFD0 U293 ( .I(n409), .Z(n408) );
  BUFFD0 U294 ( .I(n410), .Z(n409) );
  BUFFD0 U295 ( .I(n411), .Z(n410) );
  BUFFD0 U296 ( .I(n412), .Z(n411) );
  BUFFD0 U297 ( .I(n413), .Z(n412) );
  BUFFD0 U298 ( .I(n414), .Z(n413) );
  BUFFD0 U299 ( .I(n415), .Z(n414) );
  BUFFD0 U300 ( .I(n416), .Z(n415) );
  BUFFD0 U301 ( .I(n417), .Z(n416) );
  BUFFD0 U302 ( .I(n418), .Z(n417) );
  BUFFD0 U303 ( .I(n419), .Z(n418) );
  BUFFD0 U304 ( .I(n420), .Z(n419) );
  BUFFD0 U305 ( .I(n422), .Z(n420) );
  BUFFD0 U306 ( .I(n423), .Z(n421) );
  BUFFD0 U307 ( .I(n424), .Z(n422) );
  BUFFD0 U308 ( .I(n425), .Z(n423) );
  BUFFD0 U309 ( .I(n1687), .Z(n424) );
  BUFFD0 U310 ( .I(n1089), .Z(n425) );
  BUFFD0 U311 ( .I(n429), .Z(n426) );
  BUFFD0 U312 ( .I(n1693), .Z(n427) );
  BUFFD0 U313 ( .I(n427), .Z(n428) );
  BUFFD0 U314 ( .I(n430), .Z(n429) );
  BUFFD0 U315 ( .I(n431), .Z(n430) );
  BUFFD0 U316 ( .I(n432), .Z(n431) );
  BUFFD0 U317 ( .I(n433), .Z(n432) );
  BUFFD0 U318 ( .I(n434), .Z(n433) );
  BUFFD0 U319 ( .I(n435), .Z(n434) );
  BUFFD0 U320 ( .I(n436), .Z(n435) );
  BUFFD0 U321 ( .I(n437), .Z(n436) );
  BUFFD0 U322 ( .I(n438), .Z(n437) );
  BUFFD0 U323 ( .I(n439), .Z(n438) );
  BUFFD0 U324 ( .I(n440), .Z(n439) );
  BUFFD0 U325 ( .I(n441), .Z(n440) );
  BUFFD0 U326 ( .I(n442), .Z(n441) );
  BUFFD0 U327 ( .I(n443), .Z(n442) );
  BUFFD0 U328 ( .I(n444), .Z(n443) );
  BUFFD0 U329 ( .I(n445), .Z(n444) );
  BUFFD0 U330 ( .I(n446), .Z(n445) );
  BUFFD0 U331 ( .I(n447), .Z(n446) );
  BUFFD0 U332 ( .I(n448), .Z(n447) );
  BUFFD0 U333 ( .I(n449), .Z(n448) );
  BUFFD0 U334 ( .I(n450), .Z(n449) );
  BUFFD0 U335 ( .I(n451), .Z(n450) );
  BUFFD0 U336 ( .I(n452), .Z(n451) );
  BUFFD0 U337 ( .I(n453), .Z(n452) );
  BUFFD0 U338 ( .I(n454), .Z(n453) );
  BUFFD0 U339 ( .I(n455), .Z(n454) );
  BUFFD0 U340 ( .I(n456), .Z(n455) );
  BUFFD0 U341 ( .I(n457), .Z(n456) );
  BUFFD0 U342 ( .I(n458), .Z(n457) );
  BUFFD0 U343 ( .I(n459), .Z(n458) );
  BUFFD0 U344 ( .I(n460), .Z(n459) );
  BUFFD0 U345 ( .I(n461), .Z(n460) );
  BUFFD0 U346 ( .I(n462), .Z(n461) );
  BUFFD0 U347 ( .I(n463), .Z(n462) );
  BUFFD0 U348 ( .I(n464), .Z(n463) );
  BUFFD0 U349 ( .I(n465), .Z(n464) );
  BUFFD0 U350 ( .I(n466), .Z(n465) );
  BUFFD0 U351 ( .I(n467), .Z(n466) );
  BUFFD0 U352 ( .I(n468), .Z(n467) );
  BUFFD0 U353 ( .I(n469), .Z(n468) );
  BUFFD0 U354 ( .I(n470), .Z(n469) );
  BUFFD0 U355 ( .I(n471), .Z(n470) );
  BUFFD0 U356 ( .I(n472), .Z(n471) );
  BUFFD0 U357 ( .I(n473), .Z(n472) );
  BUFFD0 U358 ( .I(n474), .Z(n473) );
  BUFFD0 U359 ( .I(n475), .Z(n474) );
  BUFFD0 U360 ( .I(n476), .Z(n475) );
  BUFFD0 U361 ( .I(n477), .Z(n476) );
  BUFFD0 U362 ( .I(n478), .Z(n477) );
  BUFFD0 U363 ( .I(n479), .Z(n478) );
  BUFFD0 U364 ( .I(n480), .Z(n479) );
  BUFFD0 U365 ( .I(n481), .Z(n480) );
  BUFFD0 U366 ( .I(n482), .Z(n481) );
  BUFFD0 U367 ( .I(n483), .Z(n482) );
  BUFFD0 U368 ( .I(n484), .Z(n483) );
  BUFFD0 U369 ( .I(n485), .Z(n484) );
  IOA22D0 U370 ( .B1(n1682), .B2(n1788), .A1(n1788), .A2(OldWriteAr[3]), .ZN(
        n1693) );
  BUFFD0 U371 ( .I(n486), .Z(n485) );
  BUFFD0 U372 ( .I(n487), .Z(n486) );
  BUFFD0 U373 ( .I(n428), .Z(n487) );
  BUFFD0 U374 ( .I(n490), .Z(n488) );
  BUFFD0 U375 ( .I(OldWriteAr[1]), .Z(n489) );
  BUFFD0 U376 ( .I(n491), .Z(n490) );
  BUFFD0 U377 ( .I(n492), .Z(n491) );
  BUFFD0 U378 ( .I(n493), .Z(n492) );
  BUFFD0 U379 ( .I(n494), .Z(n493) );
  BUFFD0 U380 ( .I(n497), .Z(n494) );
  BUFFD0 U381 ( .I(n496), .Z(n495) );
  BUFFD0 U382 ( .I(n489), .Z(n496) );
  BUFFD0 U383 ( .I(n498), .Z(n497) );
  BUFFD0 U384 ( .I(n499), .Z(n498) );
  BUFFD0 U385 ( .I(n500), .Z(n499) );
  BUFFD0 U386 ( .I(n501), .Z(n500) );
  BUFFD0 U387 ( .I(n502), .Z(n501) );
  BUFFD0 U388 ( .I(n503), .Z(n502) );
  BUFFD0 U389 ( .I(n504), .Z(n503) );
  BUFFD0 U390 ( .I(n505), .Z(n504) );
  BUFFD0 U391 ( .I(n506), .Z(n505) );
  BUFFD0 U392 ( .I(n507), .Z(n506) );
  BUFFD0 U393 ( .I(n508), .Z(n507) );
  BUFFD0 U394 ( .I(n509), .Z(n508) );
  BUFFD0 U395 ( .I(n510), .Z(n509) );
  BUFFD0 U396 ( .I(n511), .Z(n510) );
  BUFFD0 U397 ( .I(n512), .Z(n511) );
  BUFFD0 U398 ( .I(n513), .Z(n512) );
  BUFFD0 U399 ( .I(n514), .Z(n513) );
  BUFFD0 U400 ( .I(n515), .Z(n514) );
  BUFFD0 U401 ( .I(n516), .Z(n515) );
  BUFFD0 U402 ( .I(n517), .Z(n516) );
  BUFFD0 U403 ( .I(n518), .Z(n517) );
  BUFFD0 U404 ( .I(n519), .Z(n518) );
  BUFFD0 U405 ( .I(n520), .Z(n519) );
  BUFFD0 U406 ( .I(n521), .Z(n520) );
  BUFFD0 U407 ( .I(n522), .Z(n521) );
  BUFFD0 U408 ( .I(n523), .Z(n522) );
  BUFFD0 U409 ( .I(n524), .Z(n523) );
  BUFFD0 U410 ( .I(n525), .Z(n524) );
  BUFFD0 U411 ( .I(n526), .Z(n525) );
  BUFFD0 U412 ( .I(n527), .Z(n526) );
  BUFFD0 U413 ( .I(n528), .Z(n527) );
  BUFFD0 U414 ( .I(n529), .Z(n528) );
  BUFFD0 U415 ( .I(n530), .Z(n529) );
  BUFFD0 U416 ( .I(n531), .Z(n530) );
  BUFFD0 U417 ( .I(n532), .Z(n531) );
  BUFFD0 U418 ( .I(n533), .Z(n532) );
  BUFFD0 U419 ( .I(n534), .Z(n533) );
  BUFFD0 U420 ( .I(n535), .Z(n534) );
  BUFFD0 U421 ( .I(n536), .Z(n535) );
  BUFFD0 U422 ( .I(n537), .Z(n536) );
  BUFFD0 U423 ( .I(n538), .Z(n537) );
  BUFFD0 U424 ( .I(n539), .Z(n538) );
  BUFFD0 U425 ( .I(n540), .Z(n539) );
  BUFFD0 U426 ( .I(n541), .Z(n540) );
  BUFFD0 U427 ( .I(n542), .Z(n541) );
  BUFFD0 U428 ( .I(n543), .Z(n542) );
  BUFFD0 U429 ( .I(n544), .Z(n543) );
  BUFFD0 U430 ( .I(n545), .Z(n544) );
  BUFFD0 U431 ( .I(n546), .Z(n545) );
  BUFFD0 U432 ( .I(n547), .Z(n546) );
  BUFFD0 U433 ( .I(n548), .Z(n547) );
  BUFFD0 U434 ( .I(n549), .Z(n548) );
  MOAI22D0 U435 ( .A1(n1788), .A2(n1787), .B1(n1788), .B2(n495), .ZN(n1694) );
  BUFFD0 U436 ( .I(n1694), .Z(n549) );
  BUFFD0 U437 ( .I(n551), .Z(n550) );
  BUFFD0 U438 ( .I(n552), .Z(n551) );
  BUFFD0 U439 ( .I(n553), .Z(n552) );
  BUFFD0 U440 ( .I(n554), .Z(n553) );
  BUFFD0 U441 ( .I(n555), .Z(n554) );
  BUFFD0 U442 ( .I(n556), .Z(n555) );
  BUFFD0 U443 ( .I(n557), .Z(n556) );
  BUFFD0 U444 ( .I(n558), .Z(n557) );
  BUFFD0 U445 ( .I(n559), .Z(n558) );
  BUFFD0 U446 ( .I(n560), .Z(n559) );
  BUFFD0 U447 ( .I(n561), .Z(n560) );
  BUFFD0 U448 ( .I(n562), .Z(n561) );
  BUFFD0 U449 ( .I(n563), .Z(n562) );
  BUFFD0 U450 ( .I(n564), .Z(n563) );
  BUFFD0 U451 ( .I(n565), .Z(n564) );
  BUFFD0 U452 ( .I(n566), .Z(n565) );
  BUFFD0 U453 ( .I(n567), .Z(n566) );
  BUFFD0 U454 ( .I(n568), .Z(n567) );
  BUFFD0 U455 ( .I(n569), .Z(n568) );
  BUFFD0 U456 ( .I(n570), .Z(n569) );
  BUFFD0 U457 ( .I(n571), .Z(n570) );
  BUFFD0 U458 ( .I(n572), .Z(n571) );
  BUFFD0 U459 ( .I(n573), .Z(n572) );
  BUFFD0 U460 ( .I(n574), .Z(n573) );
  BUFFD0 U461 ( .I(n575), .Z(n574) );
  BUFFD0 U462 ( .I(n576), .Z(n575) );
  BUFFD0 U463 ( .I(n577), .Z(n576) );
  BUFFD0 U464 ( .I(n578), .Z(n577) );
  BUFFD0 U465 ( .I(n579), .Z(n578) );
  BUFFD0 U466 ( .I(n580), .Z(n579) );
  BUFFD0 U467 ( .I(n581), .Z(n580) );
  BUFFD0 U468 ( .I(n582), .Z(n581) );
  BUFFD0 U469 ( .I(n583), .Z(n582) );
  BUFFD0 U470 ( .I(n584), .Z(n583) );
  BUFFD0 U471 ( .I(n585), .Z(n584) );
  BUFFD0 U472 ( .I(n586), .Z(n585) );
  BUFFD0 U473 ( .I(n587), .Z(n586) );
  BUFFD0 U474 ( .I(n588), .Z(n587) );
  BUFFD0 U475 ( .I(n589), .Z(n588) );
  BUFFD0 U476 ( .I(n590), .Z(n589) );
  BUFFD0 U477 ( .I(n591), .Z(n590) );
  BUFFD0 U478 ( .I(n592), .Z(n591) );
  BUFFD0 U479 ( .I(n593), .Z(n592) );
  BUFFD0 U480 ( .I(n594), .Z(n593) );
  BUFFD0 U481 ( .I(n595), .Z(n594) );
  BUFFD0 U482 ( .I(n596), .Z(n595) );
  BUFFD0 U483 ( .I(n597), .Z(n596) );
  BUFFD0 U484 ( .I(n598), .Z(n597) );
  BUFFD0 U485 ( .I(n599), .Z(n598) );
  BUFFD0 U486 ( .I(n600), .Z(n599) );
  BUFFD0 U487 ( .I(n601), .Z(n600) );
  BUFFD0 U488 ( .I(n602), .Z(n601) );
  BUFFD0 U489 ( .I(n603), .Z(n602) );
  BUFFD0 U490 ( .I(n604), .Z(n603) );
  BUFFD0 U491 ( .I(n605), .Z(n604) );
  BUFFD0 U492 ( .I(n606), .Z(n605) );
  BUFFD0 U493 ( .I(n607), .Z(n606) );
  BUFFD0 U494 ( .I(n608), .Z(n607) );
  BUFFD0 U495 ( .I(n609), .Z(n608) );
  BUFFD0 U496 ( .I(n610), .Z(n609) );
  BUFFD0 U497 ( .I(n1695), .Z(n610) );
  IOA22D0 U498 ( .B1(n1680), .B2(n1788), .A1(n1788), .A2(n973), .ZN(n1695) );
  BUFFD0 U499 ( .I(n612), .Z(n611) );
  BUFFD0 U500 ( .I(n613), .Z(n612) );
  BUFFD0 U501 ( .I(n614), .Z(n613) );
  BUFFD0 U502 ( .I(n615), .Z(n614) );
  BUFFD0 U503 ( .I(n616), .Z(n615) );
  BUFFD0 U504 ( .I(n617), .Z(n616) );
  BUFFD0 U505 ( .I(n618), .Z(n617) );
  BUFFD0 U506 ( .I(n619), .Z(n618) );
  BUFFD0 U507 ( .I(n620), .Z(n619) );
  BUFFD0 U508 ( .I(n621), .Z(n620) );
  BUFFD0 U509 ( .I(n622), .Z(n621) );
  BUFFD0 U510 ( .I(n623), .Z(n622) );
  BUFFD0 U511 ( .I(n624), .Z(n623) );
  BUFFD0 U512 ( .I(n625), .Z(n624) );
  BUFFD0 U513 ( .I(n626), .Z(n625) );
  BUFFD0 U514 ( .I(n627), .Z(n626) );
  BUFFD0 U515 ( .I(n628), .Z(n627) );
  BUFFD0 U516 ( .I(n629), .Z(n628) );
  BUFFD0 U517 ( .I(n630), .Z(n629) );
  BUFFD0 U518 ( .I(n631), .Z(n630) );
  BUFFD0 U519 ( .I(n632), .Z(n631) );
  BUFFD0 U520 ( .I(n633), .Z(n632) );
  BUFFD0 U521 ( .I(n634), .Z(n633) );
  BUFFD0 U522 ( .I(n635), .Z(n634) );
  BUFFD0 U523 ( .I(n636), .Z(n635) );
  BUFFD0 U524 ( .I(n637), .Z(n636) );
  BUFFD0 U525 ( .I(n638), .Z(n637) );
  BUFFD0 U526 ( .I(n639), .Z(n638) );
  BUFFD0 U527 ( .I(n640), .Z(n639) );
  BUFFD0 U528 ( .I(n641), .Z(n640) );
  BUFFD0 U529 ( .I(n642), .Z(n641) );
  BUFFD0 U530 ( .I(n643), .Z(n642) );
  BUFFD0 U531 ( .I(n644), .Z(n643) );
  BUFFD0 U532 ( .I(n645), .Z(n644) );
  BUFFD0 U533 ( .I(n646), .Z(n645) );
  BUFFD0 U534 ( .I(n647), .Z(n646) );
  BUFFD0 U535 ( .I(n648), .Z(n647) );
  BUFFD0 U536 ( .I(n649), .Z(n648) );
  BUFFD0 U537 ( .I(n650), .Z(n649) );
  BUFFD0 U538 ( .I(n651), .Z(n650) );
  BUFFD0 U539 ( .I(n652), .Z(n651) );
  BUFFD0 U540 ( .I(n653), .Z(n652) );
  BUFFD0 U541 ( .I(n654), .Z(n653) );
  BUFFD0 U542 ( .I(n655), .Z(n654) );
  BUFFD0 U543 ( .I(n656), .Z(n655) );
  BUFFD0 U544 ( .I(n657), .Z(n656) );
  BUFFD0 U545 ( .I(n658), .Z(n657) );
  BUFFD0 U546 ( .I(n659), .Z(n658) );
  BUFFD0 U547 ( .I(n660), .Z(n659) );
  BUFFD0 U548 ( .I(n661), .Z(n660) );
  BUFFD0 U549 ( .I(n662), .Z(n661) );
  BUFFD0 U550 ( .I(n663), .Z(n662) );
  BUFFD0 U551 ( .I(n664), .Z(n663) );
  BUFFD0 U552 ( .I(n665), .Z(n664) );
  BUFFD0 U553 ( .I(n666), .Z(n665) );
  BUFFD0 U554 ( .I(n667), .Z(n666) );
  BUFFD0 U555 ( .I(n668), .Z(n667) );
  BUFFD0 U556 ( .I(n669), .Z(n668) );
  BUFFD0 U557 ( .I(n670), .Z(n669) );
  BUFFD0 U558 ( .I(n671), .Z(n670) );
  BUFFD0 U559 ( .I(n1696), .Z(n671) );
  IOA22D0 U560 ( .B1(n1681), .B2(n1788), .A1(n1788), .A2(n972), .ZN(n1696) );
  MOAI22D0 U561 ( .A1(n1684), .A2(n1793), .B1(n1793), .B2(n675), .ZN(n1699) );
  BUFFD0 U562 ( .I(n673), .Z(n672) );
  BUFFD0 U563 ( .I(n674), .Z(n673) );
  BUFFD0 U564 ( .I(n676), .Z(n674) );
  BUFFD0 U565 ( .I(n725), .Z(n675) );
  BUFFD0 U566 ( .I(n677), .Z(n676) );
  BUFFD0 U567 ( .I(n678), .Z(n677) );
  BUFFD0 U568 ( .I(n679), .Z(n678) );
  BUFFD0 U569 ( .I(n680), .Z(n679) );
  BUFFD0 U570 ( .I(n681), .Z(n680) );
  BUFFD0 U571 ( .I(n682), .Z(n681) );
  BUFFD0 U572 ( .I(n683), .Z(n682) );
  BUFFD0 U573 ( .I(n684), .Z(n683) );
  BUFFD0 U574 ( .I(n685), .Z(n684) );
  BUFFD0 U575 ( .I(n686), .Z(n685) );
  BUFFD0 U576 ( .I(n687), .Z(n686) );
  BUFFD0 U577 ( .I(n688), .Z(n687) );
  BUFFD0 U578 ( .I(n689), .Z(n688) );
  BUFFD0 U579 ( .I(n690), .Z(n689) );
  BUFFD0 U580 ( .I(n691), .Z(n690) );
  BUFFD0 U581 ( .I(n692), .Z(n691) );
  BUFFD0 U582 ( .I(n693), .Z(n692) );
  BUFFD0 U583 ( .I(n694), .Z(n693) );
  BUFFD0 U584 ( .I(n695), .Z(n694) );
  BUFFD0 U585 ( .I(n696), .Z(n695) );
  BUFFD0 U586 ( .I(n697), .Z(n696) );
  BUFFD0 U587 ( .I(n698), .Z(n697) );
  BUFFD0 U588 ( .I(n699), .Z(n698) );
  BUFFD0 U589 ( .I(n700), .Z(n699) );
  BUFFD0 U590 ( .I(n701), .Z(n700) );
  BUFFD0 U591 ( .I(n702), .Z(n701) );
  BUFFD0 U592 ( .I(n703), .Z(n702) );
  BUFFD0 U593 ( .I(n704), .Z(n703) );
  BUFFD0 U594 ( .I(n705), .Z(n704) );
  BUFFD0 U595 ( .I(n706), .Z(n705) );
  BUFFD0 U596 ( .I(n707), .Z(n706) );
  BUFFD0 U597 ( .I(n708), .Z(n707) );
  BUFFD0 U598 ( .I(n709), .Z(n708) );
  BUFFD0 U599 ( .I(n710), .Z(n709) );
  BUFFD0 U600 ( .I(n711), .Z(n710) );
  BUFFD0 U601 ( .I(n712), .Z(n711) );
  BUFFD0 U602 ( .I(n713), .Z(n712) );
  BUFFD0 U603 ( .I(n714), .Z(n713) );
  BUFFD0 U604 ( .I(n715), .Z(n714) );
  BUFFD0 U605 ( .I(n716), .Z(n715) );
  BUFFD0 U606 ( .I(n717), .Z(n716) );
  BUFFD0 U607 ( .I(n718), .Z(n717) );
  BUFFD0 U608 ( .I(n719), .Z(n718) );
  BUFFD0 U609 ( .I(n720), .Z(n719) );
  BUFFD0 U610 ( .I(n721), .Z(n720) );
  BUFFD0 U611 ( .I(n722), .Z(n721) );
  BUFFD0 U612 ( .I(n723), .Z(n722) );
  BUFFD0 U613 ( .I(n724), .Z(n723) );
  BUFFD0 U614 ( .I(n726), .Z(n724) );
  BUFFD0 U615 ( .I(n727), .Z(n725) );
  BUFFD0 U616 ( .I(n728), .Z(n726) );
  BUFFD0 U617 ( .I(n729), .Z(n727) );
  BUFFD0 U618 ( .I(n1699), .Z(n728) );
  BUFFD0 U619 ( .I(n1088), .Z(n729) );
  BUFFD0 U620 ( .I(n251), .Z(n730) );
  BUFFD0 U621 ( .I(n730), .Z(n731) );
  BUFFD0 U622 ( .I(n731), .Z(n732) );
  BUFFD0 U623 ( .I(n732), .Z(n733) );
  BUFFD0 U624 ( .I(n733), .Z(n734) );
  BUFFD0 U625 ( .I(n734), .Z(n735) );
  BUFFD0 U626 ( .I(n735), .Z(n736) );
  BUFFD0 U627 ( .I(n736), .Z(n737) );
  BUFFD0 U628 ( .I(n737), .Z(n738) );
  BUFFD0 U629 ( .I(n738), .Z(n739) );
  BUFFD0 U630 ( .I(n739), .Z(n740) );
  BUFFD0 U631 ( .I(n740), .Z(n741) );
  BUFFD0 U632 ( .I(n741), .Z(n742) );
  BUFFD0 U633 ( .I(n742), .Z(n743) );
  BUFFD0 U634 ( .I(n743), .Z(n744) );
  BUFFD0 U635 ( .I(n744), .Z(n745) );
  BUFFD0 U636 ( .I(n745), .Z(n746) );
  BUFFD0 U637 ( .I(n746), .Z(n747) );
  BUFFD0 U638 ( .I(n747), .Z(n748) );
  BUFFD0 U639 ( .I(n748), .Z(n749) );
  BUFFD0 U640 ( .I(n749), .Z(n750) );
  BUFFD0 U641 ( .I(n750), .Z(n751) );
  BUFFD0 U642 ( .I(n751), .Z(n752) );
  BUFFD0 U643 ( .I(n752), .Z(n753) );
  BUFFD0 U644 ( .I(n753), .Z(n754) );
  BUFFD0 U645 ( .I(n754), .Z(n755) );
  BUFFD0 U646 ( .I(n755), .Z(n756) );
  BUFFD0 U647 ( .I(n756), .Z(n757) );
  BUFFD0 U648 ( .I(n757), .Z(n758) );
  BUFFD0 U649 ( .I(n758), .Z(n759) );
  BUFFD0 U650 ( .I(n759), .Z(n760) );
  BUFFD0 U651 ( .I(n760), .Z(n761) );
  BUFFD0 U652 ( .I(n761), .Z(n762) );
  BUFFD0 U653 ( .I(n762), .Z(n763) );
  BUFFD0 U654 ( .I(n763), .Z(n764) );
  BUFFD0 U655 ( .I(n764), .Z(n765) );
  BUFFD0 U656 ( .I(n765), .Z(n766) );
  BUFFD0 U657 ( .I(n766), .Z(n767) );
  BUFFD0 U658 ( .I(n767), .Z(n768) );
  BUFFD0 U659 ( .I(n768), .Z(n769) );
  BUFFD0 U660 ( .I(n769), .Z(n770) );
  BUFFD0 U661 ( .I(n770), .Z(n771) );
  BUFFD0 U662 ( .I(n771), .Z(n772) );
  BUFFD0 U663 ( .I(n772), .Z(n773) );
  BUFFD0 U664 ( .I(n773), .Z(n774) );
  BUFFD0 U665 ( .I(n774), .Z(n775) );
  BUFFD0 U666 ( .I(n775), .Z(n776) );
  BUFFD0 U667 ( .I(n776), .Z(n777) );
  BUFFD0 U668 ( .I(n777), .Z(n778) );
  BUFFD0 U669 ( .I(n778), .Z(n779) );
  BUFFD0 U670 ( .I(n779), .Z(n780) );
  BUFFD0 U671 ( .I(n780), .Z(n781) );
  BUFFD0 U672 ( .I(n781), .Z(n782) );
  BUFFD0 U673 ( .I(n782), .Z(n783) );
  BUFFD0 U674 ( .I(n783), .Z(n784) );
  BUFFD0 U675 ( .I(n784), .Z(n785) );
  BUFFD0 U676 ( .I(n789), .Z(n786) );
  BUFFD0 U677 ( .I(n1689), .Z(n787) );
  BUFFD0 U678 ( .I(n787), .Z(n788) );
  BUFFD0 U679 ( .I(n790), .Z(n789) );
  BUFFD0 U680 ( .I(n796), .Z(n790) );
  BUFFD0 U681 ( .I(n792), .Z(n791) );
  BUFFD0 U682 ( .I(n793), .Z(n792) );
  BUFFD0 U683 ( .I(n794), .Z(n793) );
  BUFFD0 U684 ( .I(n795), .Z(n794) );
  BUFFD0 U685 ( .I(n1702), .Z(n795) );
  BUFFD0 U686 ( .I(n797), .Z(n796) );
  BUFFD0 U687 ( .I(n798), .Z(n797) );
  BUFFD0 U688 ( .I(n799), .Z(n798) );
  BUFFD0 U689 ( .I(n800), .Z(n799) );
  BUFFD0 U690 ( .I(n801), .Z(n800) );
  BUFFD0 U691 ( .I(n802), .Z(n801) );
  BUFFD0 U692 ( .I(n803), .Z(n802) );
  BUFFD0 U693 ( .I(n804), .Z(n803) );
  BUFFD0 U694 ( .I(n805), .Z(n804) );
  BUFFD0 U695 ( .I(n806), .Z(n805) );
  BUFFD0 U696 ( .I(n807), .Z(n806) );
  BUFFD0 U697 ( .I(n808), .Z(n807) );
  BUFFD0 U698 ( .I(n809), .Z(n808) );
  BUFFD0 U699 ( .I(n810), .Z(n809) );
  BUFFD0 U700 ( .I(n811), .Z(n810) );
  BUFFD0 U701 ( .I(n812), .Z(n811) );
  BUFFD0 U702 ( .I(n813), .Z(n812) );
  BUFFD0 U703 ( .I(n814), .Z(n813) );
  BUFFD0 U704 ( .I(n815), .Z(n814) );
  BUFFD0 U705 ( .I(n816), .Z(n815) );
  BUFFD0 U706 ( .I(n817), .Z(n816) );
  BUFFD0 U707 ( .I(n818), .Z(n817) );
  BUFFD0 U708 ( .I(n819), .Z(n818) );
  BUFFD0 U709 ( .I(n820), .Z(n819) );
  BUFFD0 U710 ( .I(n821), .Z(n820) );
  BUFFD0 U711 ( .I(n822), .Z(n821) );
  BUFFD0 U712 ( .I(n823), .Z(n822) );
  BUFFD0 U713 ( .I(n824), .Z(n823) );
  BUFFD0 U714 ( .I(n825), .Z(n824) );
  BUFFD0 U715 ( .I(n826), .Z(n825) );
  BUFFD0 U716 ( .I(n827), .Z(n826) );
  BUFFD0 U717 ( .I(n828), .Z(n827) );
  BUFFD0 U718 ( .I(n829), .Z(n828) );
  BUFFD0 U719 ( .I(n830), .Z(n829) );
  BUFFD0 U720 ( .I(n831), .Z(n830) );
  BUFFD0 U721 ( .I(n832), .Z(n831) );
  BUFFD0 U722 ( .I(n833), .Z(n832) );
  BUFFD0 U723 ( .I(n834), .Z(n833) );
  BUFFD0 U724 ( .I(n835), .Z(n834) );
  BUFFD0 U725 ( .I(n836), .Z(n835) );
  BUFFD0 U726 ( .I(n837), .Z(n836) );
  BUFFD0 U727 ( .I(n838), .Z(n837) );
  BUFFD0 U728 ( .I(n839), .Z(n838) );
  BUFFD0 U729 ( .I(n840), .Z(n839) );
  BUFFD0 U730 ( .I(n841), .Z(n840) );
  BUFFD0 U731 ( .I(n842), .Z(n841) );
  BUFFD0 U732 ( .I(n843), .Z(n842) );
  BUFFD0 U733 ( .I(n844), .Z(n843) );
  BUFFD0 U734 ( .I(n845), .Z(n844) );
  BUFFD0 U735 ( .I(n846), .Z(n845) );
  BUFFD0 U736 ( .I(n847), .Z(n846) );
  BUFFD0 U737 ( .I(n788), .Z(n847) );
  BUFFD0 U738 ( .I(n851), .Z(n848) );
  BUFFD0 U739 ( .I(n1690), .Z(n849) );
  BUFFD0 U740 ( .I(n849), .Z(n850) );
  BUFFD0 U741 ( .I(n852), .Z(n851) );
  BUFFD0 U742 ( .I(n858), .Z(n852) );
  BUFFD0 U743 ( .I(n854), .Z(n853) );
  BUFFD0 U744 ( .I(n855), .Z(n854) );
  BUFFD0 U745 ( .I(n856), .Z(n855) );
  BUFFD0 U746 ( .I(n857), .Z(n856) );
  BUFFD0 U747 ( .I(n1703), .Z(n857) );
  BUFFD0 U748 ( .I(n859), .Z(n858) );
  BUFFD0 U749 ( .I(n860), .Z(n859) );
  BUFFD0 U750 ( .I(n861), .Z(n860) );
  BUFFD0 U751 ( .I(n862), .Z(n861) );
  BUFFD0 U752 ( .I(n863), .Z(n862) );
  BUFFD0 U753 ( .I(n864), .Z(n863) );
  BUFFD0 U754 ( .I(n865), .Z(n864) );
  BUFFD0 U755 ( .I(n866), .Z(n865) );
  BUFFD0 U756 ( .I(n867), .Z(n866) );
  BUFFD0 U757 ( .I(n868), .Z(n867) );
  BUFFD0 U758 ( .I(n869), .Z(n868) );
  BUFFD0 U759 ( .I(n870), .Z(n869) );
  BUFFD0 U760 ( .I(n871), .Z(n870) );
  BUFFD0 U761 ( .I(n872), .Z(n871) );
  BUFFD0 U762 ( .I(n873), .Z(n872) );
  BUFFD0 U763 ( .I(n874), .Z(n873) );
  BUFFD0 U764 ( .I(n875), .Z(n874) );
  BUFFD0 U765 ( .I(n876), .Z(n875) );
  BUFFD0 U766 ( .I(n877), .Z(n876) );
  BUFFD0 U767 ( .I(n878), .Z(n877) );
  BUFFD0 U768 ( .I(n879), .Z(n878) );
  BUFFD0 U769 ( .I(n880), .Z(n879) );
  BUFFD0 U770 ( .I(n881), .Z(n880) );
  BUFFD0 U771 ( .I(n882), .Z(n881) );
  BUFFD0 U772 ( .I(n883), .Z(n882) );
  BUFFD0 U773 ( .I(n884), .Z(n883) );
  BUFFD0 U774 ( .I(n885), .Z(n884) );
  BUFFD0 U775 ( .I(n886), .Z(n885) );
  BUFFD0 U776 ( .I(n887), .Z(n886) );
  BUFFD0 U777 ( .I(n888), .Z(n887) );
  BUFFD0 U778 ( .I(n889), .Z(n888) );
  BUFFD0 U779 ( .I(n890), .Z(n889) );
  BUFFD0 U780 ( .I(n891), .Z(n890) );
  BUFFD0 U781 ( .I(n892), .Z(n891) );
  BUFFD0 U782 ( .I(n893), .Z(n892) );
  BUFFD0 U783 ( .I(n894), .Z(n893) );
  BUFFD0 U784 ( .I(n895), .Z(n894) );
  BUFFD0 U785 ( .I(n896), .Z(n895) );
  BUFFD0 U786 ( .I(n897), .Z(n896) );
  BUFFD0 U787 ( .I(n898), .Z(n897) );
  BUFFD0 U788 ( .I(n899), .Z(n898) );
  BUFFD0 U789 ( .I(n900), .Z(n899) );
  BUFFD0 U790 ( .I(n901), .Z(n900) );
  BUFFD0 U791 ( .I(n902), .Z(n901) );
  BUFFD0 U792 ( .I(n903), .Z(n902) );
  BUFFD0 U793 ( .I(n904), .Z(n903) );
  BUFFD0 U794 ( .I(n905), .Z(n904) );
  BUFFD0 U795 ( .I(n906), .Z(n905) );
  BUFFD0 U796 ( .I(n907), .Z(n906) );
  BUFFD0 U797 ( .I(n908), .Z(n907) );
  BUFFD0 U798 ( .I(n909), .Z(n908) );
  BUFFD0 U799 ( .I(n850), .Z(n909) );
  BUFFD0 U800 ( .I(n913), .Z(n910) );
  BUFFD0 U801 ( .I(n1692), .Z(n911) );
  BUFFD0 U802 ( .I(n911), .Z(n912) );
  BUFFD0 U803 ( .I(n914), .Z(n913) );
  BUFFD0 U804 ( .I(n920), .Z(n914) );
  BUFFD0 U805 ( .I(n916), .Z(n915) );
  BUFFD0 U806 ( .I(n917), .Z(n916) );
  BUFFD0 U807 ( .I(n918), .Z(n917) );
  BUFFD0 U808 ( .I(n919), .Z(n918) );
  BUFFD0 U809 ( .I(n1704), .Z(n919) );
  BUFFD0 U810 ( .I(n921), .Z(n920) );
  BUFFD0 U811 ( .I(n922), .Z(n921) );
  BUFFD0 U812 ( .I(n923), .Z(n922) );
  BUFFD0 U813 ( .I(n924), .Z(n923) );
  BUFFD0 U814 ( .I(n925), .Z(n924) );
  BUFFD0 U815 ( .I(n926), .Z(n925) );
  BUFFD0 U816 ( .I(n927), .Z(n926) );
  BUFFD0 U817 ( .I(n928), .Z(n927) );
  BUFFD0 U818 ( .I(n929), .Z(n928) );
  BUFFD0 U819 ( .I(n930), .Z(n929) );
  BUFFD0 U820 ( .I(n931), .Z(n930) );
  BUFFD0 U821 ( .I(n932), .Z(n931) );
  BUFFD0 U822 ( .I(n933), .Z(n932) );
  BUFFD0 U823 ( .I(n934), .Z(n933) );
  BUFFD0 U824 ( .I(n935), .Z(n934) );
  BUFFD0 U825 ( .I(n936), .Z(n935) );
  BUFFD0 U826 ( .I(n937), .Z(n936) );
  BUFFD0 U827 ( .I(n938), .Z(n937) );
  BUFFD0 U828 ( .I(n939), .Z(n938) );
  BUFFD0 U829 ( .I(n940), .Z(n939) );
  BUFFD0 U830 ( .I(n941), .Z(n940) );
  BUFFD0 U831 ( .I(n942), .Z(n941) );
  BUFFD0 U832 ( .I(n943), .Z(n942) );
  BUFFD0 U833 ( .I(n944), .Z(n943) );
  BUFFD0 U834 ( .I(n945), .Z(n944) );
  BUFFD0 U835 ( .I(n946), .Z(n945) );
  BUFFD0 U836 ( .I(n947), .Z(n946) );
  BUFFD0 U837 ( .I(n948), .Z(n947) );
  BUFFD0 U838 ( .I(n949), .Z(n948) );
  BUFFD0 U839 ( .I(n950), .Z(n949) );
  BUFFD0 U840 ( .I(n951), .Z(n950) );
  BUFFD0 U841 ( .I(n952), .Z(n951) );
  BUFFD0 U842 ( .I(n953), .Z(n952) );
  BUFFD0 U843 ( .I(n954), .Z(n953) );
  BUFFD0 U844 ( .I(n955), .Z(n954) );
  BUFFD0 U845 ( .I(n956), .Z(n955) );
  BUFFD0 U846 ( .I(n957), .Z(n956) );
  BUFFD0 U847 ( .I(n958), .Z(n957) );
  BUFFD0 U848 ( .I(n959), .Z(n958) );
  BUFFD0 U849 ( .I(n960), .Z(n959) );
  BUFFD0 U850 ( .I(n961), .Z(n960) );
  BUFFD0 U851 ( .I(n962), .Z(n961) );
  BUFFD0 U852 ( .I(n963), .Z(n962) );
  BUFFD0 U853 ( .I(n964), .Z(n963) );
  BUFFD0 U854 ( .I(n965), .Z(n964) );
  BUFFD0 U855 ( .I(n966), .Z(n965) );
  BUFFD0 U856 ( .I(n967), .Z(n966) );
  BUFFD0 U857 ( .I(n968), .Z(n967) );
  BUFFD0 U858 ( .I(n969), .Z(n968) );
  BUFFD0 U859 ( .I(n970), .Z(n969) );
  BUFFD0 U860 ( .I(n971), .Z(n970) );
  BUFFD0 U861 ( .I(n912), .Z(n971) );
  BUFFD0 U862 ( .I(OldWriteAr[2]), .Z(n972) );
  BUFFD0 U863 ( .I(OldWriteAr[0]), .Z(n973) );
  BUFFD0 U864 ( .I(n1691), .Z(n974) );
  BUFFD0 U865 ( .I(n974), .Z(n975) );
  BUFFD0 U866 ( .I(n977), .Z(n976) );
  BUFFD0 U867 ( .I(n978), .Z(n977) );
  BUFFD0 U868 ( .I(n979), .Z(n978) );
  BUFFD0 U869 ( .I(n980), .Z(n979) );
  BUFFD0 U870 ( .I(n981), .Z(n980) );
  BUFFD0 U871 ( .I(n982), .Z(n981) );
  BUFFD0 U872 ( .I(n983), .Z(n982) );
  BUFFD0 U873 ( .I(n984), .Z(n983) );
  BUFFD0 U874 ( .I(n985), .Z(n984) );
  BUFFD0 U875 ( .I(n986), .Z(n985) );
  BUFFD0 U876 ( .I(n987), .Z(n986) );
  BUFFD0 U877 ( .I(n988), .Z(n987) );
  BUFFD0 U878 ( .I(n989), .Z(n988) );
  BUFFD0 U879 ( .I(n990), .Z(n989) );
  BUFFD0 U880 ( .I(n991), .Z(n990) );
  BUFFD0 U881 ( .I(n992), .Z(n991) );
  BUFFD0 U882 ( .I(n993), .Z(n992) );
  BUFFD0 U883 ( .I(n994), .Z(n993) );
  BUFFD0 U884 ( .I(n995), .Z(n994) );
  BUFFD0 U885 ( .I(n996), .Z(n995) );
  BUFFD0 U886 ( .I(n997), .Z(n996) );
  BUFFD0 U887 ( .I(n998), .Z(n997) );
  BUFFD0 U888 ( .I(n999), .Z(n998) );
  BUFFD0 U889 ( .I(n1000), .Z(n999) );
  BUFFD0 U890 ( .I(n1001), .Z(n1000) );
  BUFFD0 U891 ( .I(n1002), .Z(n1001) );
  BUFFD0 U892 ( .I(n1003), .Z(n1002) );
  BUFFD0 U893 ( .I(n1004), .Z(n1003) );
  BUFFD0 U894 ( .I(n1005), .Z(n1004) );
  BUFFD0 U895 ( .I(n1006), .Z(n1005) );
  BUFFD0 U896 ( .I(n1007), .Z(n1006) );
  BUFFD0 U897 ( .I(n1008), .Z(n1007) );
  BUFFD0 U898 ( .I(n1009), .Z(n1008) );
  BUFFD0 U899 ( .I(n1010), .Z(n1009) );
  BUFFD0 U900 ( .I(n1011), .Z(n1010) );
  BUFFD0 U901 ( .I(n1012), .Z(n1011) );
  BUFFD0 U902 ( .I(n1013), .Z(n1012) );
  BUFFD0 U903 ( .I(n1014), .Z(n1013) );
  BUFFD0 U904 ( .I(n1015), .Z(n1014) );
  BUFFD0 U905 ( .I(n1016), .Z(n1015) );
  BUFFD0 U906 ( .I(n1017), .Z(n1016) );
  BUFFD0 U907 ( .I(n1018), .Z(n1017) );
  BUFFD0 U908 ( .I(n1019), .Z(n1018) );
  BUFFD0 U909 ( .I(n1020), .Z(n1019) );
  BUFFD0 U910 ( .I(n1021), .Z(n1020) );
  BUFFD0 U911 ( .I(n1022), .Z(n1021) );
  BUFFD0 U912 ( .I(n1025), .Z(n1022) );
  BUFFD0 U913 ( .I(n785), .Z(n1023) );
  BUFFD0 U914 ( .I(n1026), .Z(n1024) );
  BUFFD0 U915 ( .I(n1028), .Z(n1025) );
  BUFFD0 U916 ( .I(n1035), .Z(n1026) );
  CKBXD0 U917 ( .I(n1023), .Z(WriteCmd) );
  BUFFD0 U918 ( .I(n1029), .Z(n1028) );
  BUFFD0 U919 ( .I(n1030), .Z(n1029) );
  BUFFD0 U920 ( .I(n1031), .Z(n1030) );
  BUFFD0 U921 ( .I(n1032), .Z(n1031) );
  BUFFD0 U922 ( .I(n1033), .Z(n1032) );
  BUFFD0 U923 ( .I(n1034), .Z(n1033) );
  BUFFD0 U924 ( .I(n975), .Z(n1034) );
  BUFFD0 U925 ( .I(n1776), .Z(n1035) );
  BUFFD0 U926 ( .I(n1041), .Z(n1036) );
  BUFFD0 U927 ( .I(n1688), .Z(n1037) );
  BUFFD0 U928 ( .I(n1037), .Z(n1038) );
  BUFFD0 U929 ( .I(n1038), .Z(n1039) );
  BUFFD0 U930 ( .I(n1039), .Z(n1040) );
  BUFFD0 U931 ( .I(n1042), .Z(n1041) );
  BUFFD0 U932 ( .I(n1043), .Z(n1042) );
  BUFFD0 U933 ( .I(n1044), .Z(n1043) );
  BUFFD0 U934 ( .I(n1045), .Z(n1044) );
  BUFFD0 U935 ( .I(n1046), .Z(n1045) );
  BUFFD0 U936 ( .I(n1047), .Z(n1046) );
  BUFFD0 U937 ( .I(n1048), .Z(n1047) );
  BUFFD0 U938 ( .I(n1049), .Z(n1048) );
  BUFFD0 U939 ( .I(n1050), .Z(n1049) );
  BUFFD0 U940 ( .I(n1051), .Z(n1050) );
  BUFFD0 U941 ( .I(n1052), .Z(n1051) );
  BUFFD0 U942 ( .I(n1053), .Z(n1052) );
  BUFFD0 U943 ( .I(n1054), .Z(n1053) );
  BUFFD0 U944 ( .I(n1055), .Z(n1054) );
  BUFFD0 U945 ( .I(n1056), .Z(n1055) );
  BUFFD0 U946 ( .I(n1057), .Z(n1056) );
  BUFFD0 U947 ( .I(n1058), .Z(n1057) );
  BUFFD0 U948 ( .I(n1059), .Z(n1058) );
  BUFFD0 U949 ( .I(n1060), .Z(n1059) );
  BUFFD0 U950 ( .I(n1061), .Z(n1060) );
  BUFFD0 U951 ( .I(n1062), .Z(n1061) );
  BUFFD0 U952 ( .I(n1063), .Z(n1062) );
  BUFFD0 U953 ( .I(n1064), .Z(n1063) );
  BUFFD0 U954 ( .I(n1065), .Z(n1064) );
  BUFFD0 U955 ( .I(n1066), .Z(n1065) );
  BUFFD0 U956 ( .I(n1067), .Z(n1066) );
  BUFFD0 U957 ( .I(n1068), .Z(n1067) );
  BUFFD0 U958 ( .I(n1069), .Z(n1068) );
  BUFFD0 U959 ( .I(n1070), .Z(n1069) );
  BUFFD0 U960 ( .I(n1071), .Z(n1070) );
  BUFFD0 U961 ( .I(n1072), .Z(n1071) );
  BUFFD0 U962 ( .I(n1073), .Z(n1072) );
  BUFFD0 U963 ( .I(n1074), .Z(n1073) );
  BUFFD0 U964 ( .I(n1075), .Z(n1074) );
  BUFFD0 U965 ( .I(n1076), .Z(n1075) );
  BUFFD0 U966 ( .I(n1077), .Z(n1076) );
  BUFFD0 U967 ( .I(n1078), .Z(n1077) );
  BUFFD0 U968 ( .I(n1079), .Z(n1078) );
  BUFFD0 U969 ( .I(n1080), .Z(n1079) );
  BUFFD0 U970 ( .I(n1081), .Z(n1080) );
  BUFFD0 U971 ( .I(n1082), .Z(n1081) );
  BUFFD0 U972 ( .I(n1083), .Z(n1082) );
  BUFFD0 U973 ( .I(n1084), .Z(n1083) );
  BUFFD0 U974 ( .I(n1085), .Z(n1084) );
  BUFFD0 U975 ( .I(n1086), .Z(n1085) );
  BUFFD0 U976 ( .I(n1087), .Z(n1086) );
  BUFFD0 U977 ( .I(n1098), .Z(n1087) );
  BUFFD0 U978 ( .I(n1092), .Z(n1088) );
  BUFFD0 U979 ( .I(n1093), .Z(n1089) );
  BUFFD0 U980 ( .I(n1094), .Z(n1090) );
  BUFFD0 U981 ( .I(n1095), .Z(n1091) );
  BUFFD0 U982 ( .I(n1096), .Z(n1092) );
  BUFFD0 U983 ( .I(n1097), .Z(n1093) );
  CKND2D0 U984 ( .A1(ReadCmd), .A2(n1388), .ZN(n1719) );
  BUFFD0 U985 ( .I(n307), .Z(n1094) );
  BUFFD0 U986 ( .I(n365), .Z(n1095) );
  BUFFD0 U987 ( .I(n1099), .Z(n1096) );
  BUFFD0 U988 ( .I(n1100), .Z(n1097) );
  BUFFD0 U989 ( .I(n1101), .Z(n1098) );
  BUFFD0 U990 ( .I(OldReadAr[1]), .Z(n1099) );
  BUFFD0 U991 ( .I(OldReadAr[0]), .Z(n1100) );
  BUFFD0 U992 ( .I(n1102), .Z(n1101) );
  BUFFD0 U993 ( .I(n1104), .Z(n1102) );
  BUFFD0 U994 ( .I(n1717), .Z(n1103) );
  BUFFD0 U995 ( .I(n1040), .Z(n1104) );
  BUFFD0 U996 ( .I(n1110), .Z(n1105) );
  BUFFD0 U997 ( .I(N68), .Z(n1106) );
  BUFFD0 U998 ( .I(n1106), .Z(n1107) );
  BUFFD0 U999 ( .I(n1107), .Z(n1108) );
  BUFFD0 U1000 ( .I(n1108), .Z(n1109) );
  BUFFD0 U1001 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1002 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1003 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1004 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1005 ( .I(n1115), .Z(n1114) );
  BUFFD0 U1006 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1007 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1008 ( .I(n1118), .Z(n1117) );
  BUFFD0 U1009 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1010 ( .I(n1120), .Z(n1119) );
  BUFFD0 U1011 ( .I(n1121), .Z(n1120) );
  BUFFD0 U1012 ( .I(n1122), .Z(n1121) );
  BUFFD0 U1013 ( .I(n1123), .Z(n1122) );
  BUFFD0 U1014 ( .I(n1124), .Z(n1123) );
  BUFFD0 U1015 ( .I(n1125), .Z(n1124) );
  BUFFD0 U1016 ( .I(n1126), .Z(n1125) );
  BUFFD0 U1017 ( .I(n1127), .Z(n1126) );
  BUFFD0 U1018 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1019 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1020 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1021 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1022 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1023 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1024 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1025 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1026 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1027 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1028 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1029 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1030 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1031 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1032 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1033 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1034 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1035 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1036 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1037 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1038 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1039 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1040 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1041 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1042 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1043 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1044 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1045 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1046 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1047 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1048 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1049 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1050 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1051 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1052 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1053 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1054 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1055 ( .I(n1109), .Z(n1164) );
  BUFFD0 U1056 ( .I(n1800), .Z(n1165) );
  CKBD0 U1057 ( .CLK(n1165), .C(ReadCmd) );
  CKBD0 U1058 ( .CLK(n1725), .C(n1220) );
  BUFFD0 U1059 ( .I(n1169), .Z(n1167) );
  BUFFD0 U1060 ( .I(n1170), .Z(n1168) );
  BUFFD0 U1061 ( .I(n1171), .Z(n1169) );
  BUFFD0 U1062 ( .I(n1172), .Z(n1170) );
  BUFFD0 U1063 ( .I(n1173), .Z(n1171) );
  BUFFD0 U1064 ( .I(n1174), .Z(n1172) );
  BUFFD0 U1065 ( .I(n1175), .Z(n1173) );
  BUFFD0 U1066 ( .I(n1176), .Z(n1174) );
  BUFFD0 U1067 ( .I(n1177), .Z(n1175) );
  BUFFD0 U1068 ( .I(n1178), .Z(n1176) );
  BUFFD0 U1069 ( .I(n1179), .Z(n1177) );
  BUFFD0 U1070 ( .I(n1180), .Z(n1178) );
  BUFFD0 U1071 ( .I(n1181), .Z(n1179) );
  BUFFD0 U1072 ( .I(n1182), .Z(n1180) );
  BUFFD0 U1073 ( .I(n1183), .Z(n1181) );
  BUFFD0 U1074 ( .I(n1184), .Z(n1182) );
  BUFFD0 U1075 ( .I(n1185), .Z(n1183) );
  BUFFD0 U1076 ( .I(n1186), .Z(n1184) );
  BUFFD0 U1077 ( .I(n1187), .Z(n1185) );
  BUFFD0 U1078 ( .I(n1188), .Z(n1186) );
  BUFFD0 U1079 ( .I(n1189), .Z(n1187) );
  BUFFD0 U1080 ( .I(n1190), .Z(n1188) );
  BUFFD0 U1081 ( .I(n1191), .Z(n1189) );
  BUFFD0 U1082 ( .I(n1192), .Z(n1190) );
  BUFFD0 U1083 ( .I(n1198), .Z(n1191) );
  BUFFD0 U1084 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1085 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1086 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1087 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1088 ( .I(n1197), .Z(n1196) );
  CKBD0 U1089 ( .CLK(n1686), .C(n1493) );
  BUFFD0 U1090 ( .I(n1199), .Z(n1197) );
  BUFFD0 U1091 ( .I(N51), .Z(n1198) );
  BUFFD0 U1092 ( .I(n1200), .Z(n1199) );
  BUFFD0 U1093 ( .I(n1201), .Z(n1200) );
  BUFFD0 U1094 ( .I(n1202), .Z(n1201) );
  BUFFD0 U1095 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1096 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1097 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1098 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1099 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1100 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1101 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1102 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1103 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1104 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1105 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1106 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1107 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1108 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1109 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1110 ( .I(n1218), .Z(n1217) );
  BUFFD0 U1111 ( .I(n1219), .Z(n1218) );
  BUFFD0 U1112 ( .I(n1220), .Z(n1219) );
  XNR2D0 U1113 ( .A1(n1493), .A2(n1708), .ZN(n1725) );
  BUFFD0 U1114 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1115 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1116 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1117 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1118 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1119 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1120 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1121 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1122 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1123 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1124 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1125 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1126 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1127 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1128 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1129 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1130 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1131 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1132 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1133 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1134 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1135 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1136 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1137 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1138 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1139 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1140 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1141 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1142 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1143 ( .I(n1251), .Z(n1250) );
  BUFFD0 U1144 ( .I(n1252), .Z(n1251) );
  BUFFD0 U1145 ( .I(n1253), .Z(n1252) );
  BUFFD0 U1146 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1147 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1148 ( .I(n1256), .Z(n1255) );
  BUFFD0 U1149 ( .I(n1257), .Z(n1256) );
  BUFFD0 U1150 ( .I(n1258), .Z(n1257) );
  BUFFD0 U1151 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1152 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1153 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1154 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1155 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1156 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1157 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1158 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1159 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1160 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1161 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1162 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1163 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1164 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1165 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1166 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1167 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1168 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1169 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1170 ( .I(N49), .Z(n1277) );
  CKBD0 U1171 ( .CLK(ReadAddr[2]), .C(n1278) );
  OAI21D0 U1172 ( .A1(n1707), .A2(n1278), .B(n1708), .ZN(n1723) );
  BUFFD0 U1173 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1174 ( .I(n1282), .Z(n1280) );
  BUFFD0 U1175 ( .I(n1283), .Z(n1281) );
  BUFFD0 U1176 ( .I(n1284), .Z(n1282) );
  BUFFD0 U1177 ( .I(n1285), .Z(n1283) );
  BUFFD0 U1178 ( .I(n1286), .Z(n1284) );
  BUFFD0 U1179 ( .I(n1287), .Z(n1285) );
  BUFFD0 U1180 ( .I(n1288), .Z(n1286) );
  BUFFD0 U1181 ( .I(n1289), .Z(n1287) );
  BUFFD0 U1182 ( .I(n1290), .Z(n1288) );
  BUFFD0 U1183 ( .I(n1291), .Z(n1289) );
  BUFFD0 U1184 ( .I(n1292), .Z(n1290) );
  BUFFD0 U1185 ( .I(n1293), .Z(n1291) );
  BUFFD0 U1186 ( .I(n1294), .Z(n1292) );
  BUFFD0 U1187 ( .I(n1295), .Z(n1293) );
  BUFFD0 U1188 ( .I(n1296), .Z(n1294) );
  BUFFD0 U1189 ( .I(n1297), .Z(n1295) );
  BUFFD0 U1190 ( .I(n1298), .Z(n1296) );
  BUFFD0 U1191 ( .I(n1299), .Z(n1297) );
  BUFFD0 U1192 ( .I(n1300), .Z(n1298) );
  BUFFD0 U1193 ( .I(n1301), .Z(n1299) );
  BUFFD0 U1194 ( .I(n1302), .Z(n1300) );
  BUFFD0 U1195 ( .I(n1303), .Z(n1301) );
  BUFFD0 U1196 ( .I(n1304), .Z(n1302) );
  BUFFD0 U1197 ( .I(n1305), .Z(n1303) );
  BUFFD0 U1198 ( .I(n1306), .Z(n1304) );
  BUFFD0 U1199 ( .I(n1307), .Z(n1305) );
  BUFFD0 U1200 ( .I(n1308), .Z(n1306) );
  BUFFD0 U1201 ( .I(n1309), .Z(n1307) );
  BUFFD0 U1202 ( .I(N48), .Z(n1308) );
  BUFFD0 U1203 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1204 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1205 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1206 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1207 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1208 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1209 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1210 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1211 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1212 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1213 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1214 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1215 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1216 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1217 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1218 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1219 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1220 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1221 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1222 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1223 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1224 ( .I(n1706), .Z(n1330) );
  BUFFD0 U1225 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1226 ( .I(ReadAddr[1]), .Z(n1332) );
  XNR2D0 U1227 ( .A1(n1331), .A2(n1334), .ZN(n1706) );
  BUFFD0 U1228 ( .I(n1335), .Z(n1333) );
  BUFFD0 U1229 ( .I(n1336), .Z(n1334) );
  BUFFD0 U1230 ( .I(n1337), .Z(n1335) );
  BUFFD0 U1231 ( .I(n1338), .Z(n1336) );
  BUFFD0 U1232 ( .I(n1339), .Z(n1337) );
  BUFFD0 U1233 ( .I(n1340), .Z(n1338) );
  BUFFD0 U1234 ( .I(n1341), .Z(n1339) );
  BUFFD0 U1235 ( .I(n1342), .Z(n1340) );
  BUFFD0 U1236 ( .I(n1343), .Z(n1341) );
  BUFFD0 U1237 ( .I(n1344), .Z(n1342) );
  BUFFD0 U1238 ( .I(n1345), .Z(n1343) );
  BUFFD0 U1239 ( .I(n1346), .Z(n1344) );
  BUFFD0 U1240 ( .I(n1347), .Z(n1345) );
  BUFFD0 U1241 ( .I(n1348), .Z(n1346) );
  BUFFD0 U1242 ( .I(n1349), .Z(n1347) );
  BUFFD0 U1243 ( .I(n1350), .Z(n1348) );
  BUFFD0 U1244 ( .I(n1351), .Z(n1349) );
  BUFFD0 U1245 ( .I(n1352), .Z(n1350) );
  BUFFD0 U1246 ( .I(n1353), .Z(n1351) );
  BUFFD0 U1247 ( .I(n1354), .Z(n1352) );
  BUFFD0 U1248 ( .I(n1355), .Z(n1353) );
  BUFFD0 U1249 ( .I(n1356), .Z(n1354) );
  BUFFD0 U1250 ( .I(n1357), .Z(n1355) );
  BUFFD0 U1251 ( .I(n1358), .Z(n1356) );
  BUFFD0 U1252 ( .I(n1359), .Z(n1357) );
  BUFFD0 U1253 ( .I(n1360), .Z(n1358) );
  BUFFD0 U1254 ( .I(n1361), .Z(n1359) );
  BUFFD0 U1255 ( .I(n1362), .Z(n1360) );
  BUFFD0 U1256 ( .I(n1363), .Z(n1361) );
  BUFFD0 U1257 ( .I(n1364), .Z(n1362) );
  BUFFD0 U1258 ( .I(n1365), .Z(n1363) );
  BUFFD0 U1259 ( .I(n1366), .Z(n1364) );
  BUFFD0 U1260 ( .I(n1367), .Z(n1365) );
  BUFFD0 U1261 ( .I(n1368), .Z(n1366) );
  BUFFD0 U1262 ( .I(n1369), .Z(n1367) );
  BUFFD0 U1263 ( .I(n1370), .Z(n1368) );
  BUFFD0 U1264 ( .I(N47), .Z(n1369) );
  BUFFD0 U1265 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1266 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1267 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1268 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1269 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1270 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1271 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1272 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1273 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1274 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1275 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1276 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1277 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1278 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1279 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1280 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1281 ( .I(ReadAddr[0]), .Z(n1386) );
  BUFFD0 U1282 ( .I(n1389), .Z(n1387) );
  BUFFD0 U1283 ( .I(n1390), .Z(n1388) );
  BUFFD0 U1284 ( .I(n1391), .Z(n1389) );
  BUFFD0 U1285 ( .I(n1392), .Z(n1390) );
  BUFFD0 U1286 ( .I(n1393), .Z(n1391) );
  BUFFD0 U1287 ( .I(n1394), .Z(n1392) );
  BUFFD0 U1288 ( .I(n1395), .Z(n1393) );
  BUFFD0 U1289 ( .I(n1396), .Z(n1394) );
  BUFFD0 U1290 ( .I(n1397), .Z(n1395) );
  BUFFD0 U1291 ( .I(n1398), .Z(n1396) );
  BUFFD0 U1292 ( .I(n1415), .Z(n1397) );
  BUFFD0 U1293 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1294 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1295 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1296 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1297 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1298 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1299 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1300 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1301 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1302 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1303 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1304 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1305 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1306 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1307 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1308 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1309 ( .I(n2), .Z(n1414) );
  BUFFD0 U1310 ( .I(N50), .Z(n1415) );
  BUFFD0 U1311 ( .I(n1416), .Z(n1417) );
  BUFFD0 U1312 ( .I(n1417), .Z(n1418) );
  BUFFD0 U1313 ( .I(n1418), .Z(n1419) );
  BUFFD0 U1314 ( .I(n1419), .Z(n1420) );
  BUFFD0 U1315 ( .I(n1420), .Z(n1421) );
  BUFFD0 U1316 ( .I(n1421), .Z(n1422) );
  BUFFD0 U1317 ( .I(n1422), .Z(n1423) );
  BUFFD0 U1318 ( .I(n1423), .Z(n1424) );
  BUFFD0 U1319 ( .I(n1424), .Z(n1425) );
  BUFFD0 U1320 ( .I(n1425), .Z(n1426) );
  BUFFD0 U1321 ( .I(n1426), .Z(n1427) );
  BUFFD0 U1322 ( .I(n1427), .Z(n1428) );
  BUFFD0 U1323 ( .I(n1428), .Z(n1429) );
  BUFFD0 U1324 ( .I(n1429), .Z(n1430) );
  BUFFD0 U1325 ( .I(n1430), .Z(n1431) );
  BUFFD0 U1326 ( .I(n1431), .Z(n1432) );
  BUFFD0 U1327 ( .I(n1432), .Z(n1433) );
  BUFFD0 U1328 ( .I(n1439), .Z(n1434) );
  BUFFD0 U1329 ( .I(N70), .Z(n1435) );
  BUFFD0 U1330 ( .I(n1435), .Z(n1436) );
  BUFFD0 U1331 ( .I(n1436), .Z(n1437) );
  BUFFD0 U1332 ( .I(n1437), .Z(n1438) );
  BUFFD0 U1333 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1334 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1335 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1336 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1337 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1338 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1339 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1340 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1341 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1342 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1343 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1344 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1345 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1346 ( .I(n1453), .Z(n1452) );
  BUFFD0 U1347 ( .I(n1454), .Z(n1453) );
  BUFFD0 U1348 ( .I(n1455), .Z(n1454) );
  BUFFD0 U1349 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1350 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1351 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1352 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1353 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1354 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1355 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1356 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1357 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1358 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1359 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1360 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1361 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1362 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1363 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1364 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1365 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1366 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1367 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1368 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1369 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1370 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1371 ( .I(n1478), .Z(n1477) );
  BUFFD0 U1372 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1373 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1374 ( .I(n1481), .Z(n1480) );
  BUFFD0 U1375 ( .I(n1482), .Z(n1481) );
  BUFFD0 U1376 ( .I(n1483), .Z(n1482) );
  BUFFD0 U1377 ( .I(n1484), .Z(n1483) );
  BUFFD0 U1378 ( .I(n1485), .Z(n1484) );
  BUFFD0 U1379 ( .I(n1486), .Z(n1485) );
  BUFFD0 U1380 ( .I(n1487), .Z(n1486) );
  BUFFD0 U1381 ( .I(n1488), .Z(n1487) );
  BUFFD0 U1382 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1383 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1384 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1385 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1386 ( .I(n1438), .Z(n1492) );
  XNR2D0 U1387 ( .A1(n1711), .A2(WriteAddr[3]), .ZN(n1738) );
  BUFFD0 U1388 ( .I(n1499), .Z(n1494) );
  BUFFD0 U1389 ( .I(N69), .Z(n1495) );
  BUFFD0 U1390 ( .I(n1495), .Z(n1496) );
  BUFFD0 U1391 ( .I(n1496), .Z(n1497) );
  BUFFD0 U1392 ( .I(n1497), .Z(n1498) );
  BUFFD0 U1393 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1394 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1395 ( .I(n1502), .Z(n1501) );
  BUFFD0 U1396 ( .I(n1503), .Z(n1502) );
  BUFFD0 U1397 ( .I(n1504), .Z(n1503) );
  BUFFD0 U1398 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1399 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1400 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1401 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1402 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1403 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1404 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1405 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1406 ( .I(n1513), .Z(n1512) );
  BUFFD0 U1407 ( .I(n1514), .Z(n1513) );
  BUFFD0 U1408 ( .I(n1515), .Z(n1514) );
  BUFFD0 U1409 ( .I(n1516), .Z(n1515) );
  BUFFD0 U1410 ( .I(n1517), .Z(n1516) );
  BUFFD0 U1411 ( .I(n1518), .Z(n1517) );
  BUFFD0 U1412 ( .I(n1519), .Z(n1518) );
  BUFFD0 U1413 ( .I(n1520), .Z(n1519) );
  BUFFD0 U1414 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1415 ( .I(n1522), .Z(n1521) );
  BUFFD0 U1416 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1417 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1418 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1419 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1420 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1421 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1422 ( .I(n1529), .Z(n1528) );
  BUFFD0 U1423 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1424 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1425 ( .I(n1532), .Z(n1531) );
  BUFFD0 U1426 ( .I(n1533), .Z(n1532) );
  BUFFD0 U1427 ( .I(n1534), .Z(n1533) );
  BUFFD0 U1428 ( .I(n1535), .Z(n1534) );
  BUFFD0 U1429 ( .I(n1536), .Z(n1535) );
  BUFFD0 U1430 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1431 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1432 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1433 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1434 ( .I(n1541), .Z(n1540) );
  BUFFD0 U1435 ( .I(n1542), .Z(n1541) );
  BUFFD0 U1436 ( .I(n1543), .Z(n1542) );
  BUFFD0 U1437 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1438 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1439 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1440 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1441 ( .I(n1548), .Z(n1547) );
  BUFFD0 U1442 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1443 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1444 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1445 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1446 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1447 ( .I(n1498), .Z(n1553) );
  BUFFD0 U1448 ( .I(n1559), .Z(n1554) );
  BUFFD0 U1449 ( .I(N67), .Z(n1555) );
  BUFFD0 U1450 ( .I(n1555), .Z(n1556) );
  BUFFD0 U1451 ( .I(n1556), .Z(n1557) );
  BUFFD0 U1452 ( .I(n1557), .Z(n1558) );
  BUFFD0 U1453 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1454 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1455 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1456 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1457 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1458 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1459 ( .I(n1566), .Z(n1565) );
  BUFFD0 U1460 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1461 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1462 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1463 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1464 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1465 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1466 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1467 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1468 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1469 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1470 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1471 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1472 ( .I(n1579), .Z(n1578) );
  BUFFD0 U1473 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1474 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1475 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1476 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1477 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1478 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1479 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1480 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1481 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1482 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1483 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1484 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1485 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1486 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1487 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1488 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1489 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1490 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1491 ( .I(n1598), .Z(n1597) );
  BUFFD0 U1492 ( .I(n1599), .Z(n1598) );
  BUFFD0 U1493 ( .I(n1600), .Z(n1599) );
  BUFFD0 U1494 ( .I(n1601), .Z(n1600) );
  BUFFD0 U1495 ( .I(n1602), .Z(n1601) );
  BUFFD0 U1496 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1497 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1498 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1499 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1500 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1501 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1502 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1503 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1504 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1505 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1506 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1507 ( .I(n1558), .Z(n1613) );
  BUFFD0 U1508 ( .I(N71), .Z(n1614) );
  BUFFD0 U1509 ( .I(n1614), .Z(n1615) );
  BUFFD0 U1510 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1511 ( .I(n1618), .Z(n1617) );
  BUFFD0 U1512 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1513 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1514 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1515 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1516 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1517 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1518 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1519 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1520 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1521 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1522 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1523 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1524 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1525 ( .I(n1632), .Z(n1631) );
  BUFFD0 U1526 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1527 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1528 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1529 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1530 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1531 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1532 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1533 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1534 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1535 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1536 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1537 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1538 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1539 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1540 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1541 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1542 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1543 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1544 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1545 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1546 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1547 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1548 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1549 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1550 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1551 ( .I(n1658), .Z(n1657) );
  BUFFD0 U1552 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1553 ( .I(n1660), .Z(n1659) );
  BUFFD0 U1554 ( .I(n1661), .Z(n1660) );
  BUFFD0 U1555 ( .I(n1662), .Z(n1661) );
  BUFFD0 U1556 ( .I(n1663), .Z(n1662) );
  BUFFD0 U1557 ( .I(n1615), .Z(n1663) );
  ND3D0 U1558 ( .A1(n1678), .A2(n1679), .A3(n1677), .ZN(n1798) );
  INVD0 U1559 ( .I(n1780), .ZN(n1791) );
  BUFFD0 U1560 ( .I(n1433), .Z(n1664) );
  INVD1 U1561 ( .I(n1676), .ZN(n1675) );
  BUFFD1 U1562 ( .I(Reset), .Z(n1676) );
  INVD1 U1563 ( .I(n1676), .ZN(n1674) );
  ND2D1 U1564 ( .A1(n1767), .A2(n1791), .ZN(n1718) );
  INVD1 U1565 ( .I(n1785), .ZN(n1784) );
  INVD1 U1566 ( .I(n1793), .ZN(n1795) );
  MAOI22D0 U1567 ( .A1(n5), .A2(n1679), .B1(n1679), .B2(n1763), .ZN(n1767) );
  OAI211D1 U1568 ( .A1(n1798), .A2(n1770), .B(n1767), .C(n1722), .ZN(n1785) );
  INR2D1 U1569 ( .A1(n1763), .B1(n1721), .ZN(n1722) );
  AOI21D1 U1570 ( .A1(n1781), .A2(n1720), .B(n1679), .ZN(n1721) );
  ND2D1 U1571 ( .A1(WriteReq), .A2(n1786), .ZN(n1788) );
  ND2D1 U1572 ( .A1(ReadReq), .A2(n1718), .ZN(n1793) );
  ND2D1 U1573 ( .A1(n1767), .A2(n1798), .ZN(n1786) );
  AOI21D1 U1574 ( .A1(n1758), .A2(n1751), .B(ReadAddr[1]), .ZN(n1732) );
  INVD1 U1575 ( .I(n1731), .ZN(n1758) );
  OA211D0 U1576 ( .A1(n1759), .A2(n1758), .B(n1757), .C(n1756), .Z(n1778) );
  INVD1 U1577 ( .I(n1749), .ZN(n1757) );
  NR3D0 U1578 ( .A1(n1755), .A2(n1754), .A3(n1753), .ZN(n1756) );
  NR3D0 U1579 ( .A1(WriteAddr[2]), .A2(n1787), .A3(ReadAddr[2]), .ZN(n1754) );
  ND2D1 U1580 ( .A1(n1707), .A2(n1278), .ZN(n1708) );
  ND2D1 U1581 ( .A1(n1730), .A2(n1729), .ZN(n1749) );
  XNR2D1 U1582 ( .A1(ReadAddr[1]), .A2(n1787), .ZN(n1730) );
  INVD1 U1583 ( .I(n1746), .ZN(n1750) );
  INVD1 U1584 ( .I(n1740), .ZN(n1729) );
  ND2D1 U1585 ( .A1(n1388), .A2(n1719), .ZN(N50) );
  NR3D0 U1586 ( .A1(n1720), .A2(n1713), .A3(n1712), .ZN(n1714) );
  XNR2D1 U1587 ( .A1(ReadAddr[3]), .A2(n1090), .ZN(n1712) );
  XNR2D1 U1588 ( .A1(ReadAddr[2]), .A2(n1091), .ZN(n1713) );
  XNR2D1 U1589 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n1733) );
  NR2D1 U1590 ( .A1(n1723), .A2(n1719), .ZN(N49) );
  NR2D1 U1591 ( .A1(n1281), .A2(n1719), .ZN(N48) );
  NR2D1 U1592 ( .A1(n1168), .A2(n1719), .ZN(N51) );
  NR2D1 U1593 ( .A1(n1334), .A2(n1719), .ZN(N47) );
  INVD1 U1594 ( .I(ReadReq), .ZN(n1720) );
  INVD1 U1595 ( .I(WriteReq), .ZN(n1770) );
  INVD1 U1596 ( .I(WriteAddr[1]), .ZN(n1787) );
  OAI211D1 U1597 ( .A1(n1787), .A2(ReadAddr[1]), .B(n1751), .C(n1744), .ZN(
        n1760) );
  AOI22D0 U1598 ( .A1(n1686), .A2(WriteAddr[3]), .B1(n1683), .B2(WriteAddr[0]), 
        .ZN(n1744) );
  ND2D1 U1599 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .ZN(n1709) );
  OAI21D1 U1600 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n1709), .ZN(n1724)
         );
  AOI21D1 U1601 ( .A1(n1709), .A2(n1681), .B(n1711), .ZN(n1739) );
  OAI211D1 U1602 ( .A1(n1684), .A2(WriteAddr[1]), .B(n1750), .C(n1747), .ZN(
        n1761) );
  AOI22D0 U1603 ( .A1(n1682), .A2(ReadAddr[3]), .B1(n1680), .B2(ReadAddr[0]), 
        .ZN(n1747) );
  ND2D1 U1604 ( .A1(n1678), .A2(n1781), .ZN(n1763) );
  OAI22D0 U1605 ( .A1(n1795), .A2(n1091), .B1(n1685), .B2(n1793), .ZN(n1700)
         );
  OAI22D0 U1606 ( .A1(n1795), .A2(n1090), .B1(n1686), .B2(n1793), .ZN(n1698)
         );
  NR3D0 U1607 ( .A1(n1678), .A2(n1677), .A3(n1679), .ZN(n1780) );
  ND2D1 U1608 ( .A1(n1685), .A2(WriteAddr[2]), .ZN(n1751) );
  OAI22D0 U1609 ( .A1(n1785), .A2(n915), .B1(n1784), .B2(n1783), .ZN(n1692) );
  AOI21D1 U1610 ( .A1(n1782), .A2(n1781), .B(n1780), .ZN(n1783) );
  OAI22D0 U1611 ( .A1(n1678), .A2(n1779), .B1(n1679), .B2(n1778), .ZN(n1782)
         );
  OAI22D0 U1612 ( .A1(n1785), .A2(n853), .B1(n1784), .B2(n1766), .ZN(n1690) );
  AOI31D0 U1613 ( .A1(n1765), .A2(n5), .A3(n1679), .B(n1764), .ZN(n1766) );
  IOA21D1 U1614 ( .A1(n1781), .A2(n1779), .B(n1748), .ZN(n1765) );
  OAI31D0 U1615 ( .A1(n1763), .A2(n1679), .A3(n1762), .B(n1798), .ZN(n1764) );
  OAI22D0 U1616 ( .A1(n1785), .A2(n791), .B1(n1784), .B2(n1737), .ZN(n1689) );
  AOI22D0 U1617 ( .A1(n1736), .A2(n1781), .B1(n1735), .B2(n1734), .ZN(n1737)
         );
  AOI211D1 U1618 ( .A1(n1685), .A2(n1731), .B(n1796), .C(n1749), .ZN(n1735) );
  AOI221D0 U1619 ( .A1(n1746), .A2(n1758), .B1(n1733), .B2(ReadAddr[1]), .C(
        n1732), .ZN(n1734) );
  AOI21D1 U1620 ( .A1(n1751), .A2(n1750), .B(WriteAddr[1]), .ZN(n1755) );
  NR2D1 U1621 ( .A1(WriteAddr[2]), .A2(n1685), .ZN(n1746) );
  OAI21D1 U1622 ( .A1(n1719), .A2(n1718), .B(n1103), .ZN(n1688) );
  ND4D1 U1623 ( .A1(n1716), .A2(n1718), .A3(n1715), .A4(n1714), .ZN(n1717) );
  XNR2D1 U1624 ( .A1(ReadAddr[0]), .A2(n1089), .ZN(n1716) );
  XNR2D1 U1625 ( .A1(ReadAddr[1]), .A2(n1088), .ZN(n1715) );
  OAI21D1 U1626 ( .A1(n1678), .A2(n1728), .B(n1679), .ZN(n1736) );
  NR4D0 U1627 ( .A1(n1729), .A2(n1727), .A3(n1742), .A4(n1726), .ZN(n1728) );
  XNR2D1 U1628 ( .A1(WriteAddr[2]), .A2(n1723), .ZN(n1727) );
  XNR2D1 U1629 ( .A1(WriteAddr[3]), .A2(n1725), .ZN(n1726) );
  OAI21D1 U1630 ( .A1(n1777), .A2(n1786), .B(n1024), .ZN(n1691) );
  ND4D1 U1631 ( .A1(n1775), .A2(n1786), .A3(n1774), .A4(n1773), .ZN(n1776) );
  XNR2D1 U1632 ( .A1(WriteAddr[0]), .A2(n973), .ZN(n1775) );
  XNR2D1 U1633 ( .A1(WriteAddr[2]), .A2(n972), .ZN(n1774) );
  ND4D1 U1634 ( .A1(n1743), .A2(n1742), .A3(n1741), .A4(n1740), .ZN(n1779) );
  XNR2D1 U1635 ( .A1(n1738), .A2(n1686), .ZN(n1743) );
  XNR2D1 U1636 ( .A1(ReadAddr[2]), .A2(n1739), .ZN(n1741) );
  NR2D1 U1637 ( .A1(n1709), .A2(n1681), .ZN(n1711) );
  NR2D1 U1638 ( .A1(n1787), .A2(n1681), .ZN(n1759) );
  XNR2D1 U1639 ( .A1(ReadAddr[3]), .A2(n1682), .ZN(n1731) );
  XNR2D1 U1640 ( .A1(WriteAddr[0]), .A2(n1683), .ZN(n1740) );
  NR2D1 U1641 ( .A1(n1683), .A2(n1684), .ZN(n1707) );
  XNR2D1 U1642 ( .A1(n1724), .A2(n1684), .ZN(n1742) );
  ND2D1 U1643 ( .A1(WriteCmd), .A2(n1791), .ZN(n1777) );
  OAI32D1 U1644 ( .A1(n1798), .A2(WriteReq), .A3(n1676), .B1(n1797), .B2(n11), 
        .ZN(n1701) );
  AOI21D1 U1645 ( .A1(n1796), .A2(n1798), .B(Reset), .ZN(n1797) );
  OAI22D0 U1646 ( .A1(n1684), .A2(n1791), .B1(n1724), .B2(n1777), .ZN(N68) );
  OAI22D0 U1647 ( .A1(n1493), .A2(n1791), .B1(n1738), .B2(n1777), .ZN(N70) );
  OAI22D0 U1648 ( .A1(n1685), .A2(n1791), .B1(n1710), .B2(n1777), .ZN(N69) );
  INVD1 U1649 ( .I(n1739), .ZN(n1710) );
  OAI22D0 U1650 ( .A1(n1683), .A2(n1791), .B1(WriteAddr[0]), .B2(n1777), .ZN(
        N67) );
  ND3D1 U1651 ( .A1(n1679), .A2(n5), .A3(n1677), .ZN(n1796) );
  NR3D0 U1652 ( .A1(n1772), .A2(n1771), .A3(n1770), .ZN(n1773) );
  XNR2D1 U1653 ( .A1(n1682), .A2(OldWriteAr[3]), .ZN(n1771) );
  XNR2D1 U1654 ( .A1(n1787), .A2(OldWriteAr[1]), .ZN(n1772) );
  OAI21D1 U1655 ( .A1(n1760), .A2(n1761), .B(n1677), .ZN(n1748) );
  OAI31D0 U1656 ( .A1(n1791), .A2(n1676), .A3(ReadReq), .B(n192), .ZN(n1697)
         );
  OAI21D1 U1657 ( .A1(n1789), .A2(n1676), .B(FullFIFO), .ZN(n1790) );
  ND2D1 U1658 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
endmodule


module DPMem1kx32_AWid4_DWid32_1 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [3:0] AddrR;
  input [3:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N9, N44, N45, N46, N47, ClockR, ClockW, Dreadyr, \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N84, N364, N628, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n85, n102,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];

  XNR4D1 U13 ( .A1(n527), .A2(n256), .A3(n511), .A4(n513), .ZN(n3141) );
  XOR4D1 U14 ( .A1(n232), .A2(n499), .A3(n206), .A4(n218), .Z(n3142) );
  XOR4D1 U15 ( .A1(n2932), .A2(n302), .A3(n268), .A4(n2933), .Z(n3145) );
  XOR4D1 U16 ( .A1(n353), .A2(n357), .A3(n336), .A4(n346), .Z(n3148) );
  XNR4D1 U17 ( .A1(n405), .A2(n29), .A3(n135), .A4(n398), .ZN(n3151) );
  XOR4D1 U21 ( .A1(n3136), .A2(n2671), .A3(n3135), .A4(n2670), .Z(n3137) );
  XNR4D1 U22 ( .A1(n2633), .A2(n2639), .A3(n2631), .A4(n2629), .ZN(n3135) );
  XNR4D1 U27 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n3130) );
  XOR4D1 U28 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n3131) );
  XNR4D1 U29 ( .A1(n2593), .A2(n2601), .A3(n2604), .A4(n2600), .ZN(n3133) );
  XNR4D1 U30 ( .A1(n2675), .A2(n2677), .A3(n2676), .A4(n2673), .ZN(n3139) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(n205), .E(n2946), .CP(n2985), .CDN(n3074), .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n207), .E(n2946), .CP(n2985), .CDN(n3092), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n219), .E(n2947), .CP(n2985), .CDN(n3092), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n233), .E(n2946), .CP(n2986), .CDN(n3092), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n246), .E(n2947), .CP(n2986), .CDN(n3092), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n258), .E(n2946), .CP(n2986), .CDN(n3092), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n270), .E(n2946), .CP(n2986), .CDN(n3092), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n281), .E(n2946), .CP(n2986), .CDN(n3092), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n292), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n305), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n311), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n322), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n337), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n349), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n356), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n358), .E(n2946), .CP(n2987), .CDN(n3091), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n33), .E(n2947), .CP(n2987), .CDN(n3091), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n380), .E(n2947), .CP(n2988), .CDN(n3091), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n387), .E(n2947), .CP(n2988), .CDN(n3091), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n105), .E(n2947), .CP(n2988), .CDN(n3090), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n404), .E(n2947), .CP(n2988), .CDN(n3090), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n411), .E(n2947), .CP(n2988), .CDN(n3090), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n140), .E(n2947), .CP(n2988), .CDN(n3090), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n422), .E(n2947), .CP(n2988), .CDN(n3090), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n424), .E(n2947), .CP(n2988), .CDN(n3090), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n430), .E(n2947), .CP(n2988), .CDN(n3090), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n431), .E(n2947), .CP(n2989), .CDN(n3090), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n433), .E(n2947), .CP(n2989), .CDN(n3090), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n434), .E(n2946), .CP(n2989), .CDN(n3090), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n205), .E(n2948), .CP(n2989), .CDN(n3090), .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n207), .E(n2948), .CP(n2989), .CDN(n3070), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n219), .E(n2948), .CP(n2989), .CDN(n3070), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n233), .E(n2948), .CP(n2989), .CDN(n3070), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n246), .E(n2948), .CP(n2990), .CDN(n3089), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n258), .E(n2948), .CP(n2990), .CDN(n3087), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n270), .E(n2948), .CP(n2990), .CDN(n3075), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n281), .E(n2948), .CP(n2990), .CDN(n3106), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n292), .E(n2949), .CP(n2990), .CDN(n3089), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n305), .E(n2948), .CP(n2990), .CDN(n3089), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n311), .E(n2949), .CP(n2990), .CDN(n3089), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n322), .E(n2948), .CP(n2991), .CDN(n3089), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n337), .E(n2949), .CP(n2991), .CDN(n3089), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n349), .E(n2948), .CP(n2991), .CDN(n3089), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n356), .E(n2949), .CP(n2991), .CDN(n3089), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n358), .E(n2948), .CP(n2991), .CDN(n3089), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n33), .E(n2949), .CP(n2991), .CDN(n3089), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n380), .E(n2949), .CP(n2991), .CDN(n3089), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n387), .E(n2949), .CP(n2991), .CDN(n3089), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n105), .E(n2949), .CP(n2991), .CDN(n3097), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n404), .E(n2949), .CP(n2992), .CDN(n3088), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n411), .E(n2949), .CP(n2992), .CDN(n3070), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n140), .E(n2949), .CP(n2992), .CDN(n3097), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n422), .E(n2949), .CP(n2992), .CDN(n3096), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n424), .E(n2949), .CP(n2992), .CDN(n3074), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n430), .E(n2949), .CP(n2992), .CDN(n3097), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n431), .E(n2949), .CP(n2992), .CDN(n3083), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n433), .E(n2949), .CP(n2992), .CDN(n3071), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n434), .E(n2948), .CP(n2992), .CDN(n3097), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(n205), .E(n2954), .CP(n3035), .CDN(n3091), .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n207), .E(n2954), .CP(n3051), .CDN(n3083), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n219), .E(n2954), .CP(n3045), .CDN(n3083), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n233), .E(n2954), .CP(n3025), .CDN(n3083), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n246), .E(n2954), .CP(n3025), .CDN(n3083), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n258), .E(n2954), .CP(n3052), .CDN(n3083), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n270), .E(n2955), .CP(n3027), .CDN(n3083), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n281), .E(n2955), .CP(n3038), .CDN(n3083), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n292), .E(n2955), .CP(n3039), .CDN(n3082), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n305), .E(n2955), .CP(n3037), .CDN(n3082), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n311), .E(n2955), .CP(n2978), .CDN(n3082), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n322), .E(n2955), .CP(n3041), .CDN(n3082), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n337), .E(n2955), .CP(n3032), .CDN(n3082), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n349), .E(n2955), .CP(n3047), .CDN(n3082), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n356), .E(n2955), .CP(n3046), .CDN(n3082), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n358), .E(n2955), .CP(n3048), .CDN(n3082), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n33), .E(n2954), .CP(n3051), .CDN(n3082), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n380), .E(n2954), .CP(n3026), .CDN(n3082), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n387), .E(n2955), .CP(n3050), .CDN(n3082), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n105), .E(n2955), .CP(n3031), .CDN(n3067), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n404), .E(n2955), .CP(n2997), .CDN(n3068), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n411), .E(n2954), .CP(n2997), .CDN(n3071), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n140), .E(n2955), .CP(n2997), .CDN(n3075), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n422), .E(n2954), .CP(n2997), .CDN(n3076), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n424), .E(n2954), .CP(n2997), .CDN(n3105), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n430), .E(n2954), .CP(n2997), .CDN(n3086), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n431), .E(n2955), .CP(n2997), .CDN(n3103), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n433), .E(n2955), .CP(n2997), .CDN(n3069), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n434), .E(n2954), .CP(n2997), .CDN(n3073), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(n205), .E(n2956), .CP(n2998), .CDN(n3072), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n207), .E(n2956), .CP(n2998), .CDN(n3099), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n219), .E(n2956), .CP(n2998), .CDN(n3081), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n233), .E(n2956), .CP(n2998), .CDN(n3099), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n246), .E(n2956), .CP(n2998), .CDN(n3099), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n258), .E(n2956), .CP(n2999), .CDN(n3072), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n270), .E(n2957), .CP(n2999), .CDN(n3062), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n281), .E(n2957), .CP(n2999), .CDN(n3074), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n292), .E(n2957), .CP(n2999), .CDN(n3081), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n305), .E(n2957), .CP(n2999), .CDN(n3081), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n311), .E(n2957), .CP(n2999), .CDN(n3081), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n322), .E(n2957), .CP(n2999), .CDN(n3081), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n337), .E(n2957), .CP(n2999), .CDN(n3081), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n349), .E(n2957), .CP(n2999), .CDN(n3081), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n356), .E(n2957), .CP(n3000), .CDN(n3081), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n358), .E(n2957), .CP(n3000), .CDN(n3081), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n33), .E(n2956), .CP(n3000), .CDN(n3081), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n380), .E(n2957), .CP(n3000), .CDN(n3081), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n387), .E(n2956), .CP(n3000), .CDN(n3081), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n105), .E(n2957), .CP(n3000), .CDN(n3081), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n404), .E(n2956), .CP(n3000), .CDN(n3080), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n411), .E(n2957), .CP(n3000), .CDN(n3064), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n140), .E(n2956), .CP(n3000), .CDN(n3063), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n422), .E(n2957), .CP(n3001), .CDN(n3064), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n424), .E(n2956), .CP(n3001), .CDN(n3070), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n430), .E(n2957), .CP(n3001), .CDN(n3064), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n431), .E(n2957), .CP(n3001), .CDN(n3065), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n433), .E(n2957), .CP(n3001), .CDN(n3098), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n434), .E(n2956), .CP(n3001), .CDN(n3066), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(n205), .E(n2963), .CP(n3003), .CDN(n3075), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n207), .E(n2963), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n219), .E(n2964), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n233), .E(n2963), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n246), .E(n2964), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n258), .E(n2963), .CP(n3004), .CDN(n3076), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n270), .E(n2963), .CP(n3004), .CDN(n3076), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n281), .E(n2963), .CP(n3004), .CDN(n3076), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n292), .E(n2963), .CP(n3004), .CDN(n3075), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n305), .E(n2963), .CP(n3004), .CDN(n3075), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n311), .E(n2963), .CP(n3004), .CDN(n3075), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n322), .E(n2963), .CP(n3004), .CDN(n3075), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n337), .E(n2963), .CP(n3004), .CDN(n3075), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n349), .E(n2963), .CP(n3004), .CDN(n3075), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n356), .E(n2963), .CP(n3005), .CDN(n3075), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n358), .E(n2963), .CP(n3005), .CDN(n3075), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n33), .E(n2964), .CP(n3005), .CDN(n3075), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n380), .E(n2964), .CP(n3005), .CDN(n3075), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n387), .E(n2964), .CP(n3005), .CDN(n3075), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n105), .E(n2964), .CP(n3005), .CDN(n3074), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n404), .E(n2964), .CP(n3005), .CDN(n3074), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n411), .E(n2964), .CP(n3005), .CDN(n3074), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n140), .E(n2964), .CP(n3005), .CDN(n3074), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n422), .E(n2964), .CP(n3006), .CDN(n3074), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n424), .E(n2964), .CP(n3006), .CDN(n3074), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n430), .E(n2964), .CP(n3006), .CDN(n3074), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n431), .E(n2964), .CP(n3006), .CDN(n3074), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n433), .E(n2964), .CP(n3006), .CDN(n3074), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n434), .E(n2963), .CP(n3006), .CDN(n3074), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(n205), .E(n2965), .CP(n3006), .CDN(n3074), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n207), .E(n2965), .CP(n3006), .CDN(n3073), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n219), .E(n2966), .CP(n3006), .CDN(n3067), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n233), .E(n2965), .CP(n3007), .CDN(n3102), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n246), .E(n2966), .CP(n3007), .CDN(n3102), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n258), .E(n2965), .CP(n3007), .CDN(n3101), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n270), .E(n2965), .CP(n3007), .CDN(n3073), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n281), .E(n2965), .CP(n3007), .CDN(n3102), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n292), .E(n2965), .CP(n3008), .CDN(n3067), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n305), .E(n2965), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n311), .E(n2965), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n322), .E(n2965), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n337), .E(n2965), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n349), .E(n2965), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n356), .E(n2965), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n358), .E(n2965), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n33), .E(n2966), .CP(n3008), .CDN(n3102), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n380), .E(n2966), .CP(n3009), .CDN(n3067), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n387), .E(n2966), .CP(n3009), .CDN(n3067), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n105), .E(n2966), .CP(n3009), .CDN(n3073), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n404), .E(n2966), .CP(n3009), .CDN(n3073), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n411), .E(n2966), .CP(n3009), .CDN(n3073), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n140), .E(n2966), .CP(n3009), .CDN(n3073), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n422), .E(n2966), .CP(n3009), .CDN(n3073), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n424), .E(n2966), .CP(n3009), .CDN(n3073), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n430), .E(n2966), .CP(n3009), .CDN(n3073), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n431), .E(n2966), .CP(n3010), .CDN(n3073), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n433), .E(n2966), .CP(n3010), .CDN(n3073), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n434), .E(n2965), .CP(n3010), .CDN(n3073), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(n205), .E(n2971), .CP(n3017), .CDN(n3068), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n207), .E(n2971), .CP(n3017), .CDN(n3078), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n219), .E(n2972), .CP(n3017), .CDN(n3083), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n233), .E(n2971), .CP(n3018), .CDN(n3071), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n246), .E(n2972), .CP(n3018), .CDN(n3103), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n258), .E(n2971), .CP(n3018), .CDN(n3096), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n270), .E(n2971), .CP(n3018), .CDN(n3064), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n281), .E(n2971), .CP(n3018), .CDN(n3096), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n292), .E(n2971), .CP(n3019), .CDN(n3102), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n305), .E(n2971), .CP(n3019), .CDN(n3102), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n311), .E(n2971), .CP(n3019), .CDN(n3102), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n322), .E(n2971), .CP(n3019), .CDN(n3102), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n337), .E(n2971), .CP(n3019), .CDN(n3102), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n349), .E(n2971), .CP(n3019), .CDN(n3102), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n356), .E(n2971), .CP(n3019), .CDN(n3071), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n358), .E(n2971), .CP(n3019), .CDN(n3083), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n33), .E(n2972), .CP(n3019), .CDN(n3102), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n380), .E(n2972), .CP(n3020), .CDN(n3071), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n387), .E(n2972), .CP(n3020), .CDN(n3071), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n105), .E(n2972), .CP(n3020), .CDN(n3067), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n404), .E(n2972), .CP(n3020), .CDN(n3067), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n411), .E(n2972), .CP(n3020), .CDN(n3067), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n140), .E(n2972), .CP(n3020), .CDN(n3067), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n422), .E(n2972), .CP(n3020), .CDN(n3067), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n424), .E(n2972), .CP(n3020), .CDN(n3067), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n430), .E(n2972), .CP(n3020), .CDN(n3067), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n431), .E(n2972), .CP(n3021), .CDN(n3067), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n433), .E(n2972), .CP(n3021), .CDN(n3067), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n434), .E(n2971), .CP(n3021), .CDN(n3067), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(n205), .E(n2974), .CP(n3021), .CDN(n3067), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n207), .E(n2974), .CP(n3021), .CDN(n3066), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n219), .E(n2974), .CP(n3021), .CDN(n3066), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n233), .E(n2974), .CP(n3021), .CDN(n3066), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n246), .E(n2974), .CP(n3022), .CDN(n3066), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n258), .E(n2974), .CP(n3022), .CDN(n3066), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n270), .E(n2973), .CP(n3022), .CDN(n3066), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n281), .E(n2973), .CP(n3022), .CDN(n3066), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n292), .E(n2973), .CP(n3022), .CDN(n3065), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n305), .E(n2974), .CP(n3022), .CDN(n3065), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n311), .E(n2973), .CP(n3022), .CDN(n3065), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n322), .E(n2974), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n337), .E(n2973), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n349), .E(n2974), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n356), .E(n2973), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n358), .E(n2974), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n33), .E(n2973), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n380), .E(n2973), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n387), .E(n2973), .CP(n3023), .CDN(n3065), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n105), .E(n2973), .CP(n3023), .CDN(n3064), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n404), .E(n2973), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n411), .E(n2973), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n140), .E(n2973), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n422), .E(n2973), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n424), .E(n2973), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n430), .E(n2973), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n431), .E(n2974), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n433), .E(n2974), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n434), .E(n2974), .CP(n3024), .CDN(n3064), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(n205), .E(N628), .CP(n2982), .CDN(n3075), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n207), .E(n2943), .CP(n2982), .CDN(n3079), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n219), .E(N628), .CP(n2982), .CDN(n3094), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n233), .E(N628), .CP(n2982), .CDN(n3094), 
        .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n246), .E(N628), .CP(n2982), .CDN(n3092), 
        .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n258), .E(N628), .CP(n2983), .CDN(n3094), 
        .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n270), .E(n2943), .CP(n2983), .CDN(n3077), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n281), .E(n2943), .CP(n2983), .CDN(n3092), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n292), .E(n2943), .CP(n2983), .CDN(n3093), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n305), .E(n2943), .CP(n2983), .CDN(n3093), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n311), .E(n2943), .CP(n2983), .CDN(n3093), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n322), .E(n2943), .CP(n2983), .CDN(n3093), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n337), .E(n2943), .CP(n2983), .CDN(n3093), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n349), .E(n2943), .CP(n2983), .CDN(n3093), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n356), .E(n2943), .CP(n2984), .CDN(n3093), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n358), .E(n2943), .CP(n2984), .CDN(n3093), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n33), .E(n2944), .CP(n2984), .CDN(n3093), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n380), .E(n2944), .CP(n2984), .CDN(n3093), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n387), .E(n2944), .CP(n2984), .CDN(n3093), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n105), .E(n2944), .CP(n2984), .CDN(n3093), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n404), .E(n2944), .CP(n2984), .CDN(n3093), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n411), .E(n2944), .CP(n2984), .CDN(n3092), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n140), .E(n2944), .CP(n2984), .CDN(n3091), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n422), .E(n2944), .CP(n2985), .CDN(n3090), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n424), .E(n2944), .CP(n2985), .CDN(n3093), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n430), .E(n2944), .CP(n2985), .CDN(n3094), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n431), .E(n2944), .CP(n2985), .CDN(n3092), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n433), .E(n2944), .CP(n2985), .CDN(n3091), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n434), .E(n2943), .CP(n2985), .CDN(n3090), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(n205), .E(n2950), .CP(n2993), .CDN(n3109), .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n207), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n219), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n233), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n246), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n258), .E(n2950), .CP(n2994), .CDN(n3088), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n270), .E(n2951), .CP(n2994), .CDN(n3088), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n281), .E(n2951), .CP(n2994), .CDN(n3088), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n292), .E(n2951), .CP(n2994), .CDN(n3087), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n305), .E(n2951), .CP(n2994), .CDN(n3087), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n311), .E(n2951), .CP(n2994), .CDN(n3087), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n322), .E(n2951), .CP(n2994), .CDN(n3087), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n337), .E(n2951), .CP(n2994), .CDN(n3087), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n349), .E(n2951), .CP(n2994), .CDN(n3087), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n356), .E(n2951), .CP(n2995), .CDN(n3087), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n358), .E(n2951), .CP(n2995), .CDN(n3087), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n33), .E(n2950), .CP(n2995), .CDN(n3087), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n380), .E(n2950), .CP(n2995), .CDN(n3087), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n387), .E(n2951), .CP(n2995), .CDN(n3087), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n105), .E(n2950), .CP(n2995), .CDN(n3086), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n404), .E(n2951), .CP(n2995), .CDN(n3086), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n411), .E(n2950), .CP(n2995), .CDN(n3086), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n140), .E(n2951), .CP(n2995), .CDN(n3086), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n422), .E(n2950), .CP(n2996), .CDN(n3086), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n424), .E(n2951), .CP(n2996), .CDN(n3086), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n430), .E(n2950), .CP(n2996), .CDN(n3086), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n431), .E(n2951), .CP(n2996), .CDN(n3086), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n433), .E(n2951), .CP(n2996), .CDN(n3086), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n434), .E(n2950), .CP(n2996), .CDN(n3086), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(n205), .E(n2952), .CP(n2996), .CDN(n3086), .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n207), .E(n2952), .CP(n2996), .CDN(n3085), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n219), .E(n2953), .CP(n2996), .CDN(n3085), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n233), .E(n2952), .CP(n2981), .CDN(n3085), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n246), .E(n2953), .CP(n2977), .CDN(n3085), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n258), .E(n2952), .CP(n3050), .CDN(n3085), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n270), .E(n2952), .CP(n3031), .CDN(n3085), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n281), .E(n2952), .CP(n3041), .CDN(n3085), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n292), .E(n2952), .CP(n3036), .CDN(n3084), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n305), .E(n2952), .CP(n3049), .CDN(n3084), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n311), .E(n2952), .CP(ClockW), .CDN(
        n3084), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n322), .E(n2952), .CP(n2980), .CDN(n3084), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n337), .E(n2952), .CP(n3030), .CDN(n3084), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n349), .E(n2952), .CP(n3029), .CDN(n3084), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n356), .E(n2952), .CP(n3028), .CDN(n3084), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n358), .E(n2952), .CP(n3033), .CDN(n3084), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n33), .E(n2953), .CP(n3032), .CDN(n3084), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n380), .E(n2953), .CP(n3038), .CDN(n3084), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n387), .E(n2953), .CP(n3048), .CDN(n3084), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n105), .E(n2953), .CP(n3044), .CDN(n3083), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n404), .E(n2953), .CP(n3043), .CDN(n3098), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n411), .E(n2953), .CP(n3045), .CDN(n3062), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n140), .E(n2953), .CP(n3034), .CDN(n3098), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n422), .E(n2953), .CP(n3042), .CDN(n3090), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n424), .E(n2953), .CP(n3040), .CDN(n3074), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n430), .E(n2953), .CP(n3039), .CDN(n3098), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n431), .E(n2953), .CP(n3026), .CDN(n3091), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n433), .E(n2952), .CP(n3027), .CDN(n3069), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n434), .E(n2953), .CP(n2981), .CDN(n3098), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(n205), .E(n2959), .CP(n3001), .CDN(n3063), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n207), .E(n2959), .CP(n3001), .CDN(n3080), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n219), .E(n2959), .CP(n3001), .CDN(n3080), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n233), .E(n2959), .CP(n3026), .CDN(n3080), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n246), .E(n2959), .CP(n3027), .CDN(n3080), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n258), .E(n2959), .CP(n3043), .CDN(n3080), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n270), .E(n2958), .CP(n3038), .CDN(n3080), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n281), .E(n2958), .CP(n3039), .CDN(n3080), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n292), .E(n2958), .CP(n3036), .CDN(n3079), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n305), .E(n2959), .CP(n3052), .CDN(n3079), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n311), .E(n2958), .CP(n2981), .CDN(n3079), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n322), .E(n2959), .CP(n3040), .CDN(n3079), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n337), .E(n2958), .CP(n3044), .CDN(n3079), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n349), .E(n2959), .CP(n3043), .CDN(n3079), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n356), .E(n2958), .CP(n3045), .CDN(n3079), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n358), .E(n2959), .CP(n3034), .CDN(n3079), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n33), .E(n2958), .CP(n3035), .CDN(n3079), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n380), .E(n2958), .CP(n3041), .CDN(n3079), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n387), .E(n2958), .CP(n2979), .CDN(n3079), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n105), .E(n2958), .CP(n2978), .CDN(n3078), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n404), .E(n2958), .CP(n3046), .CDN(n3078), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n411), .E(n2958), .CP(n3048), .CDN(n3078), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n140), .E(n2958), .CP(n3047), .CDN(n3078), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n422), .E(n2958), .CP(n3050), .CDN(n3078), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n424), .E(n2958), .CP(n3051), .CDN(n3078), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n430), .E(n2958), .CP(n3034), .CDN(n3078), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n431), .E(n2959), .CP(n2977), .CDN(n3078), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n433), .E(n2959), .CP(n3049), .CDN(n3078), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n434), .E(n2959), .CP(n3049), .CDN(n3078), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(n205), .E(n2962), .CP(n3051), .CDN(n3078), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n207), .E(n2962), .CP(n3050), .CDN(n3084), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n219), .E(n2962), .CP(n3040), .CDN(n3063), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n233), .E(n2962), .CP(n3052), .CDN(n3063), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n246), .E(n2962), .CP(n3033), .CDN(n3083), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n258), .E(n2962), .CP(n3031), .CDN(n3077), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n270), .E(N364), .CP(n2980), .CDN(n3074), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n281), .E(n2960), .CP(n2978), .CDN(n3085), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n292), .E(n2960), .CP(n2981), .CDN(n3077), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n305), .E(n2962), .CP(ClockW), .CDN(n3077), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n311), .E(N364), .CP(n3030), .CDN(n3077), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n322), .E(N364), .CP(n3028), .CDN(n3077), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n337), .E(N364), .CP(n3035), .CDN(n3077), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n349), .E(N364), .CP(n3049), .CDN(n3077), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n356), .E(N364), .CP(ClockW), .CDN(n3077), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n358), .E(N364), .CP(n3033), .CDN(n3077), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n33), .E(n2960), .CP(n3032), .CDN(n3077), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n380), .E(n2960), .CP(n3036), .CDN(n3077), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n387), .E(n2960), .CP(n3030), .CDN(n3077), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n105), .E(n2960), .CP(n3029), .CDN(n3076), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n404), .E(n2960), .CP(n3002), .CDN(n3078), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n411), .E(n2960), .CP(n3002), .CDN(n3114), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n140), .E(n2962), .CP(n3002), .CDN(n3079), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n422), .E(n2960), .CP(n3002), .CDN(n3077), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n424), .E(n2962), .CP(n3002), .CDN(n3068), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n430), .E(n2962), .CP(n3002), .CDN(n3100), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n431), .E(n2962), .CP(n3002), .CDN(n3069), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n433), .E(n2962), .CP(n3002), .CDN(n3068), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n434), .E(n2962), .CP(n3002), .CDN(n3100), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(n205), .E(n2967), .CP(n3010), .CDN(n3073), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n207), .E(n2967), .CP(n3010), .CDN(n3072), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n219), .E(n2968), .CP(n3010), .CDN(n3072), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n233), .E(n2967), .CP(n3010), .CDN(n3072), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n246), .E(n2968), .CP(n3011), .CDN(n3072), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n258), .E(n2967), .CP(n3011), .CDN(n3072), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n270), .E(n2967), .CP(n3011), .CDN(n3072), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n281), .E(n2967), .CP(n3011), .CDN(n3072), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n292), .E(n2967), .CP(n3011), .CDN(n3071), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n305), .E(n2967), .CP(n3011), .CDN(n3071), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n311), .E(n2967), .CP(n3011), .CDN(n3071), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n322), .E(n2967), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n337), .E(n2967), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n349), .E(n2967), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n356), .E(n2967), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n358), .E(n2967), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n33), .E(n2968), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n380), .E(n2968), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n387), .E(n2968), .CP(n3012), .CDN(n3071), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n105), .E(n2968), .CP(n3012), .CDN(n3070), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n404), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n411), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n140), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n422), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n424), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n430), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n431), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n433), .E(n2968), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n434), .E(n2967), .CP(n3013), .CDN(n3070), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(n205), .E(n2969), .CP(n3014), .CDN(n3070), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n207), .E(n2969), .CP(n3014), .CDN(n3104), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n219), .E(n2970), .CP(n3014), .CDN(n3069), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n233), .E(n2969), .CP(n3014), .CDN(n3091), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n246), .E(n2970), .CP(n3014), .CDN(n3068), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n258), .E(n2969), .CP(n3015), .CDN(n3104), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n270), .E(n2969), .CP(n3015), .CDN(n3072), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n281), .E(n2969), .CP(n3015), .CDN(n3072), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n292), .E(n2969), .CP(n3015), .CDN(n3069), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n305), .E(n2969), .CP(n3015), .CDN(n3069), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n311), .E(n2969), .CP(n3015), .CDN(n3069), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n322), .E(n2969), .CP(n3015), .CDN(n3069), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n337), .E(n2969), .CP(n3015), .CDN(n3069), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n349), .E(n2969), .CP(n3015), .CDN(n3069), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n356), .E(n2969), .CP(n3016), .CDN(n3069), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n358), .E(n2969), .CP(n3016), .CDN(n3069), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n33), .E(n2970), .CP(n3016), .CDN(n3069), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n380), .E(n2970), .CP(n3016), .CDN(n3069), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n387), .E(n2970), .CP(n3016), .CDN(n3069), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n105), .E(n2970), .CP(n3016), .CDN(n3068), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n404), .E(n2970), .CP(n3016), .CDN(n3068), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n411), .E(n2970), .CP(n3016), .CDN(n3068), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n140), .E(n2970), .CP(n3016), .CDN(n3068), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n422), .E(n2970), .CP(n3017), .CDN(n3068), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n424), .E(n2970), .CP(n3017), .CDN(n3068), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n430), .E(n2970), .CP(n3017), .CDN(n3068), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n431), .E(n2969), .CP(n3017), .CDN(n3068), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n433), .E(n2970), .CP(n3017), .CDN(n3068), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n434), .E(n2970), .CP(n3017), .CDN(n3068), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(n205), .E(n2975), .CP(n3041), .CDN(n3064), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n207), .E(n2976), .CP(n3025), .CDN(n3063), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n219), .E(n2976), .CP(ClockW), .CDN(n3063), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n233), .E(n2975), .CP(n2981), .CDN(n3063), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n246), .E(n2976), .CP(n2977), .CDN(n3063), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n258), .E(n2975), .CP(n3040), .CDN(n3063), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n270), .E(n2975), .CP(n2980), .CDN(n3063), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n281), .E(n2975), .CP(n2978), .CDN(n3063), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n292), .E(n2975), .CP(n3039), .CDN(n3101), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n305), .E(n2975), .CP(n3038), .CDN(n3075), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n311), .E(n2975), .CP(n3044), .CDN(n3090), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n322), .E(n2975), .CP(n3046), .CDN(n3072), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n337), .E(n2975), .CP(ClockW), .CDN(n3064), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n349), .E(n2975), .CP(n3037), .CDN(n3090), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n356), .E(n2975), .CP(n3034), .CDN(n3064), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n358), .E(n2975), .CP(n3027), .CDN(n3092), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n33), .E(n2976), .CP(n3030), .CDN(n3091), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n380), .E(n2976), .CP(n3029), .CDN(n3073), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n387), .E(n2976), .CP(n3028), .CDN(n3092), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n105), .E(n2976), .CP(n3033), .CDN(n3062), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n404), .E(n2976), .CP(n3032), .CDN(n3062), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n411), .E(n2976), .CP(n3031), .CDN(n3062), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n140), .E(n2976), .CP(n3035), .CDN(n3062), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n422), .E(n2976), .CP(n3032), .CDN(n3062), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n424), .E(n2976), .CP(n3026), .CDN(n3062), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n430), .E(n2976), .CP(n2979), .CDN(n3062), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n431), .E(n2975), .CP(n3036), .CDN(n3062), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n433), .E(n2975), .CP(n3042), .CDN(n3062), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n434), .E(n2976), .CP(n2980), .CDN(n3062), 
        .Q(\Storage[0][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n436), .CP(ClockR), .CDN(n3062), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n500), .E(n2947), .CP(n2986), .CDN(n3092), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n511), .E(n2946), .CP(n2986), .CDN(n3092), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n514), .E(n2947), .CP(n2986), .CDN(n3092), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n527), .E(n2946), .CP(n2986), .CDN(n3092), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n500), .E(n2948), .CP(n2989), .CDN(n3089), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n511), .E(n2948), .CP(n2989), .CDN(n3088), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n514), .E(n2948), .CP(n2990), .CDN(n3087), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n527), .E(n2948), .CP(n2990), .CDN(n3074), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n500), .E(n2954), .CP(n3037), .CDN(n3083), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n511), .E(n2954), .CP(n2979), .CDN(n3083), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n514), .E(n2954), .CP(n2979), .CDN(n3083), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n527), .E(n2954), .CP(n3035), .CDN(n3083), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n500), .E(n2956), .CP(n2998), .CDN(n3099), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n511), .E(n2956), .CP(n2998), .CDN(n3090), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n514), .E(n2956), .CP(n2998), .CDN(n3092), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n527), .E(n2956), .CP(n2998), .CDN(n3091), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n500), .E(n2964), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n511), .E(n2963), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n514), .E(n2964), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n527), .E(n2963), .CP(n3003), .CDN(n3076), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n500), .E(n2966), .CP(n3007), .CDN(n3101), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n511), .E(n2965), .CP(n3007), .CDN(n3073), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n514), .E(n2966), .CP(n3007), .CDN(n3102), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n527), .E(n2965), .CP(n3007), .CDN(n3101), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n500), .E(n2972), .CP(n3018), .CDN(n3068), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n511), .E(n2971), .CP(n3018), .CDN(n3105), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n514), .E(n2972), .CP(n3018), .CDN(n3102), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n527), .E(n2971), .CP(n3018), .CDN(n3096), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n500), .E(n2974), .CP(n3021), .CDN(n3066), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n511), .E(n2974), .CP(n3021), .CDN(n3066), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n514), .E(n2974), .CP(n3022), .CDN(n3066), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n527), .E(n2974), .CP(n3022), .CDN(n3066), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n500), .E(N628), .CP(n2982), .CDN(n3094), 
        .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n511), .E(N628), .CP(n2982), .CDN(n3101), 
        .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n514), .E(N628), .CP(n2982), .CDN(n3092), 
        .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n527), .E(N628), .CP(n2982), .CDN(n3094), 
        .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n500), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n511), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n514), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n527), .E(n2950), .CP(n2993), .CDN(n3088), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n500), .E(n2953), .CP(n3048), .CDN(n3085), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n511), .E(n2952), .CP(n3042), .CDN(n3085), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n514), .E(n2953), .CP(n3052), .CDN(n3085), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n527), .E(n2952), .CP(n2978), .CDN(n3085), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n500), .E(n2959), .CP(n3047), .CDN(n3080), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n511), .E(n2959), .CP(n3033), .CDN(n3080), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n514), .E(n2959), .CP(n3037), .CDN(n3080), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n527), .E(n2959), .CP(n3025), .CDN(n3080), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n500), .E(n2962), .CP(n2977), .CDN(n3083), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n511), .E(n2962), .CP(n2979), .CDN(n3077), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n514), .E(n2962), .CP(n3029), .CDN(n3063), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n527), .E(n2962), .CP(n3028), .CDN(n3075), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n500), .E(n2968), .CP(n3010), .CDN(n3072), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n511), .E(n2967), .CP(n3010), .CDN(n3072), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n514), .E(n2968), .CP(n3011), .CDN(n3072), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n527), .E(n2967), .CP(n3011), .CDN(n3072), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n500), .E(n2970), .CP(n3014), .CDN(n3104), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n511), .E(n2969), .CP(n3014), .CDN(n3072), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n514), .E(n2970), .CP(n3014), .CDN(n3105), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n527), .E(n2969), .CP(n3014), .CDN(n3105), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n500), .E(n2976), .CP(n3043), .CDN(n3063), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n511), .E(n2975), .CP(n3044), .CDN(n3063), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n514), .E(n2976), .CP(n3045), .CDN(n3063), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n527), .E(n2975), .CP(n3042), .CDN(n3063), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n529), .E(n3056), .CP(n3053), .CDN(n3094), 
        .Q(DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n595), .E(n3055), .CP(n3053), .CDN(n3089), 
        .Q(DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n175), .E(n3056), .CP(n3053), .CDN(n3095), 
        .Q(DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n176), .E(n3055), .CP(ClockR), .CDN(n3064), 
        .Q(DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n177), .E(n3056), .CP(ClockR), .CDN(n3066), 
        .Q(DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n859), .E(n3055), .CP(n3053), .CDN(n3062), 
        .Q(DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n178), .E(n3055), .CP(n3053), .CDN(n3063), 
        .Q(DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n179), .E(n3055), .CP(ClockR), .CDN(n3085), 
        .Q(DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n1057), .E(n3055), .CP(ClockR), .CDN(n3109), 
        .Q(DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n1123), .E(n3056), .CP(n3053), .CDN(n3077), 
        .Q(DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n1188), .E(n3055), .CP(ClockR), .CDN(n3084), 
        .Q(DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n1254), .E(n3055), .CP(ClockR), .CDN(n3095), 
        .Q(DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n1320), .E(n3055), .CP(n3053), .CDN(n3090), 
        .Q(DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n1386), .E(n3055), .CP(n3053), .CDN(n3087), 
        .Q(DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n180), .E(n3055), .CP(ClockR), .CDN(n3086), 
        .Q(DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n1515), .E(n3055), .CP(n3053), .CDN(n3090), 
        .Q(DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n1578), .E(n3055), .CP(n3053), .CDN(n3082), 
        .Q(DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n1641), .E(n3055), .CP(ClockR), .CDN(n3088), 
        .Q(DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n1703), .E(n3055), .CP(n3053), .CDN(n3070), 
        .Q(DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n1765), .E(n3055), .CP(n3053), .CDN(n3064), 
        .Q(DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n1828), .E(n3056), .CP(n3053), .CDN(n3065), 
        .Q(DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n1891), .E(n3056), .CP(n3053), .CDN(n3073), 
        .Q(DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n1952), .E(n3056), .CP(n3053), .CDN(n3091), 
        .Q(DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n2010), .E(n3056), .CP(n3053), .CDN(n3082), 
        .Q(DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n2067), .E(n3056), .CP(n3053), .CDN(n3082), 
        .Q(DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n2127), .E(n3056), .CP(n3053), .CDN(n3090), 
        .Q(DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n2186), .E(n3056), .CP(n3053), .CDN(n3082), 
        .Q(DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n181), .E(n3056), .CP(ClockR), .CDN(n3092), 
        .Q(DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n2304), .E(n3056), .CP(ClockR), .CDN(n3086), 
        .Q(DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n2360), .E(n3056), .CP(ClockR), .CDN(n3112), 
        .Q(DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n2419), .E(n183), .CP(ClockR), .CDN(n3091), 
        .Q(DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n182), .E(n183), .CP(ClockR), .CDN(n3082), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(n2542), .E(n183), .CP(ClockR), .CDN(n3067), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  BUFFD0 U3 ( .I(N84), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(n5), .Z(n4) );
  BUFFD0 U7 ( .I(n6), .Z(n5) );
  BUFFD0 U8 ( .I(n7), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(n10), .Z(n9) );
  BUFFD0 U12 ( .I(n11), .Z(n10) );
  BUFFD0 U18 ( .I(n12), .Z(n11) );
  BUFFD0 U19 ( .I(n13), .Z(n12) );
  BUFFD0 U20 ( .I(n14), .Z(n13) );
  BUFFD0 U23 ( .I(n15), .Z(n14) );
  BUFFD0 U24 ( .I(n17), .Z(n15) );
  BUFFD0 U25 ( .I(n18), .Z(n16) );
  BUFFD0 U26 ( .I(n19), .Z(n17) );
  BUFFD0 U31 ( .I(n20), .Z(n18) );
  BUFFD0 U32 ( .I(n21), .Z(n19) );
  BUFFD0 U33 ( .I(n22), .Z(n20) );
  BUFFD0 U34 ( .I(n23), .Z(n21) );
  BUFFD0 U35 ( .I(n24), .Z(n22) );
  BUFFD0 U36 ( .I(n25), .Z(n23) );
  BUFFD0 U37 ( .I(n26), .Z(n24) );
  BUFFD0 U38 ( .I(n27), .Z(n25) );
  BUFFD0 U39 ( .I(n28), .Z(n26) );
  BUFFD0 U40 ( .I(n3152), .Z(n27) );
  BUFFD0 U41 ( .I(n32), .Z(n28) );
  BUFFD0 U42 ( .I(n30), .Z(n29) );
  BUFFD0 U43 ( .I(n31), .Z(n30) );
  BUFFD0 U44 ( .I(n412), .Z(n31) );
  BUFFD0 U45 ( .I(n3151), .Z(n32) );
  BUFFD0 U46 ( .I(n34), .Z(n33) );
  BUFFD0 U47 ( .I(n35), .Z(n34) );
  BUFFD0 U48 ( .I(n36), .Z(n35) );
  BUFFD0 U49 ( .I(n37), .Z(n36) );
  BUFFD0 U50 ( .I(n38), .Z(n37) );
  BUFFD0 U51 ( .I(n39), .Z(n38) );
  BUFFD0 U52 ( .I(n40), .Z(n39) );
  BUFFD0 U53 ( .I(n41), .Z(n40) );
  BUFFD0 U54 ( .I(n42), .Z(n41) );
  BUFFD0 U55 ( .I(n43), .Z(n42) );
  BUFFD0 U56 ( .I(n44), .Z(n43) );
  BUFFD0 U57 ( .I(n45), .Z(n44) );
  BUFFD0 U58 ( .I(n46), .Z(n45) );
  BUFFD0 U59 ( .I(n47), .Z(n46) );
  BUFFD0 U60 ( .I(n48), .Z(n47) );
  BUFFD0 U61 ( .I(n49), .Z(n48) );
  BUFFD0 U62 ( .I(n51), .Z(n49) );
  BUFFD0 U63 ( .I(n57), .Z(n50) );
  BUFFD0 U64 ( .I(n52), .Z(n51) );
  BUFFD0 U65 ( .I(n53), .Z(n52) );
  BUFFD0 U66 ( .I(n54), .Z(n53) );
  BUFFD0 U67 ( .I(n55), .Z(n54) );
  BUFFD0 U68 ( .I(n56), .Z(n55) );
  BUFFD0 U69 ( .I(n365), .Z(n56) );
  BUFFD0 U70 ( .I(n58), .Z(n57) );
  BUFFD0 U71 ( .I(n59), .Z(n58) );
  BUFFD0 U72 ( .I(n60), .Z(n59) );
  BUFFD0 U73 ( .I(n61), .Z(n60) );
  BUFFD0 U74 ( .I(n62), .Z(n61) );
  BUFFD0 U75 ( .I(n63), .Z(n62) );
  BUFFD0 U76 ( .I(n64), .Z(n63) );
  BUFFD0 U77 ( .I(n85), .Z(n64) );
  BUFFD0 U78 ( .I(n102), .Z(n85) );
  BUFFD0 U79 ( .I(n104), .Z(n102) );
  BUFFD0 U80 ( .I(n364), .Z(n104) );
  BUFFD0 U81 ( .I(n106), .Z(n105) );
  BUFFD0 U82 ( .I(n107), .Z(n106) );
  BUFFD0 U83 ( .I(n108), .Z(n107) );
  BUFFD0 U84 ( .I(n109), .Z(n108) );
  BUFFD0 U85 ( .I(n110), .Z(n109) );
  BUFFD0 U86 ( .I(n111), .Z(n110) );
  BUFFD0 U87 ( .I(n112), .Z(n111) );
  BUFFD0 U88 ( .I(n113), .Z(n112) );
  BUFFD0 U89 ( .I(n114), .Z(n113) );
  BUFFD0 U90 ( .I(n115), .Z(n114) );
  BUFFD0 U91 ( .I(n116), .Z(n115) );
  BUFFD0 U92 ( .I(n117), .Z(n116) );
  BUFFD0 U93 ( .I(n118), .Z(n117) );
  BUFFD0 U94 ( .I(n119), .Z(n118) );
  BUFFD0 U95 ( .I(n120), .Z(n119) );
  BUFFD0 U96 ( .I(n121), .Z(n120) );
  BUFFD0 U97 ( .I(n122), .Z(n121) );
  BUFFD0 U98 ( .I(n123), .Z(n122) );
  BUFFD0 U99 ( .I(n124), .Z(n123) );
  BUFFD0 U100 ( .I(n125), .Z(n124) );
  BUFFD0 U101 ( .I(n126), .Z(n125) );
  BUFFD0 U102 ( .I(n127), .Z(n126) );
  BUFFD0 U103 ( .I(n128), .Z(n127) );
  BUFFD0 U104 ( .I(n129), .Z(n128) );
  BUFFD0 U105 ( .I(n130), .Z(n129) );
  BUFFD0 U106 ( .I(n131), .Z(n130) );
  BUFFD0 U107 ( .I(n132), .Z(n131) );
  BUFFD0 U108 ( .I(n133), .Z(n132) );
  BUFFD0 U109 ( .I(n134), .Z(n133) );
  BUFFD0 U110 ( .I(n136), .Z(n134) );
  BUFFD0 U111 ( .I(n137), .Z(n135) );
  BUFFD0 U112 ( .I(n389), .Z(n136) );
  BUFFD0 U113 ( .I(n138), .Z(n137) );
  BUFFD0 U114 ( .I(n139), .Z(n138) );
  BUFFD0 U115 ( .I(n388), .Z(n139) );
  BUFFD0 U116 ( .I(n141), .Z(n140) );
  BUFFD0 U117 ( .I(n142), .Z(n141) );
  BUFFD0 U118 ( .I(n143), .Z(n142) );
  BUFFD0 U119 ( .I(n144), .Z(n143) );
  BUFFD0 U120 ( .I(n145), .Z(n144) );
  BUFFD0 U121 ( .I(n146), .Z(n145) );
  BUFFD0 U122 ( .I(n147), .Z(n146) );
  BUFFD0 U123 ( .I(n148), .Z(n147) );
  BUFFD0 U124 ( .I(n149), .Z(n148) );
  BUFFD0 U125 ( .I(n150), .Z(n149) );
  BUFFD0 U126 ( .I(n151), .Z(n150) );
  BUFFD0 U127 ( .I(n152), .Z(n151) );
  BUFFD0 U128 ( .I(n153), .Z(n152) );
  BUFFD0 U129 ( .I(n154), .Z(n153) );
  BUFFD0 U130 ( .I(n155), .Z(n154) );
  BUFFD0 U131 ( .I(n156), .Z(n155) );
  BUFFD0 U132 ( .I(n157), .Z(n156) );
  BUFFD0 U133 ( .I(n158), .Z(n157) );
  BUFFD0 U134 ( .I(n159), .Z(n158) );
  BUFFD0 U135 ( .I(n160), .Z(n159) );
  BUFFD0 U136 ( .I(n161), .Z(n160) );
  BUFFD0 U137 ( .I(n162), .Z(n161) );
  BUFFD0 U138 ( .I(n163), .Z(n162) );
  BUFFD0 U139 ( .I(n164), .Z(n163) );
  BUFFD0 U140 ( .I(n165), .Z(n164) );
  BUFFD0 U141 ( .I(n166), .Z(n165) );
  BUFFD0 U142 ( .I(n167), .Z(n166) );
  BUFFD0 U143 ( .I(n168), .Z(n167) );
  BUFFD0 U144 ( .I(n169), .Z(n168) );
  BUFFD0 U145 ( .I(n170), .Z(n169) );
  BUFFD0 U146 ( .I(n171), .Z(n170) );
  BUFFD0 U147 ( .I(n172), .Z(n171) );
  BUFFD0 U148 ( .I(n173), .Z(n172) );
  BUFFD0 U149 ( .I(n174), .Z(n173) );
  BUFFD0 U150 ( .I(n413), .Z(n174) );
  CKBD0 U151 ( .CLK(N50), .C(n530) );
  CKBD0 U152 ( .CLK(N51), .C(n596) );
  BUFFD0 U153 ( .I(n661), .Z(n175) );
  BUFFD0 U154 ( .I(n727), .Z(n176) );
  BUFFD0 U155 ( .I(n793), .Z(n177) );
  CKBD0 U156 ( .CLK(N55), .C(n860) );
  BUFFD0 U157 ( .I(n925), .Z(n178) );
  BUFFD0 U158 ( .I(n991), .Z(n179) );
  BUFFD0 U159 ( .I(n1452), .Z(n180) );
  BUFFD0 U160 ( .I(n2245), .Z(n181) );
  CKBD0 U161 ( .CLK(n2696), .C(n2686) );
  CKBD0 U162 ( .CLK(n2695), .C(n2685) );
  BUFFD0 U163 ( .I(n2478), .Z(n182) );
  XOR3D4 U164 ( .A1(n2707), .A2(n2706), .A3(n3140), .Z(N82) );
  XOR3D0 U165 ( .A1(n2700), .A2(n3139), .A3(n3138), .Z(n3140) );
  BUFFD0 U166 ( .I(n2713), .Z(n183) );
  XNR3D1 U167 ( .A1(n2602), .A2(n3133), .A3(n184), .ZN(n3134) );
  XNR3D1 U168 ( .A1(n2594), .A2(n2612), .A3(n3132), .ZN(n184) );
  CKBD0 U169 ( .CLK(n203), .C(n433) );
  CKBD0 U170 ( .CLK(n204), .C(n434) );
  CKBD0 U171 ( .CLK(n202), .C(n431) );
  CKBD0 U172 ( .CLK(n199), .C(n422) );
  CKBD0 U173 ( .CLK(n338), .C(n337) );
  CKBD0 U174 ( .CLK(n306), .C(n305) );
  CKBD0 U175 ( .CLK(n359), .C(n358) );
  CKBD0 U176 ( .CLK(n312), .C(n311) );
  CKBD0 U177 ( .CLK(n293), .C(n292) );
  CKBD0 U178 ( .CLK(n271), .C(n270) );
  CKBD0 U179 ( .CLK(n259), .C(n258) );
  CKBD0 U180 ( .CLK(n501), .C(n500) );
  CKBD0 U181 ( .CLK(n208), .C(n207) );
  CKBD0 U182 ( .CLK(n282), .C(n281) );
  CKBD0 U183 ( .CLK(n247), .C(n246) );
  CKBXD0 U184 ( .I(N44), .Z(n3059) );
  BUFFD1 U185 ( .I(DataI[12]), .Z(n2923) );
  BUFFD1 U186 ( .I(DataI[9]), .Z(n2920) );
  BUFFD1 U187 ( .I(DataI[6]), .Z(n2917) );
  INVD0 U188 ( .I(N47), .ZN(n2900) );
  OR2D1 U189 ( .A1(n3124), .A2(n3120), .Z(n185) );
  OR2D1 U190 ( .A1(n3129), .A2(n3125), .Z(n186) );
  OR2D1 U191 ( .A1(n3127), .A2(n3126), .Z(n187) );
  OR2D1 U192 ( .A1(n3127), .A2(n3125), .Z(n188) );
  OR2D1 U193 ( .A1(n3129), .A2(n3126), .Z(n189) );
  INVD0 U194 ( .I(n2945), .ZN(n2943) );
  NR2XD0 U195 ( .A1(n3129), .A2(n3128), .ZN(N628) );
  INVD0 U196 ( .I(n2961), .ZN(n2960) );
  NR2XD0 U197 ( .A1(n3128), .A2(n3121), .ZN(N364) );
  OR2D1 U198 ( .A1(n3129), .A2(n3124), .Z(n190) );
  OR2D1 U199 ( .A1(n3125), .A2(n3121), .Z(n191) );
  OR2D1 U200 ( .A1(n3126), .A2(n3120), .Z(n192) );
  OR2D1 U201 ( .A1(n3127), .A2(n3124), .Z(n193) );
  OR2D1 U202 ( .A1(n3125), .A2(n3120), .Z(n194) );
  OR2D1 U203 ( .A1(n3126), .A2(n3121), .Z(n195) );
  OR2D1 U204 ( .A1(n3124), .A2(n3121), .Z(n196) );
  OR2D1 U205 ( .A1(n3128), .A2(n3127), .Z(n197) );
  OR2D1 U206 ( .A1(n3128), .A2(n3120), .Z(n198) );
  BUFFD0 U207 ( .I(n423), .Z(n199) );
  BUFFD0 U208 ( .I(n2916), .Z(n200) );
  BUFFD0 U209 ( .I(n425), .Z(n201) );
  BUFFD0 U210 ( .I(n432), .Z(n202) );
  BUFFD0 U211 ( .I(DataI[1]), .Z(n2914) );
  BUFFD0 U212 ( .I(n2914), .Z(n203) );
  BUFFD0 U213 ( .I(n435), .Z(n204) );
  XOR3D0 U214 ( .A1(n3142), .A2(n2928), .A3(n3141), .Z(n3143) );
  CKBD0 U215 ( .CLK(n1), .C(n205) );
  XOR3D0 U216 ( .A1(n432), .A2(DataI[1]), .A3(n2), .Z(N84) );
  XOR3D0 U217 ( .A1(n423), .A2(n2916), .A3(n3149), .Z(n3150) );
  XOR3D0 U218 ( .A1(n3145), .A2(n384), .A3(n3144), .Z(n3146) );
  XOR3D0 U219 ( .A1(n435), .A2(n16), .A3(n3150), .Z(n3152) );
  XOR3D0 U220 ( .A1(n50), .A2(n376), .A3(n3146), .Z(n3147) );
  XOR3D0 U221 ( .A1(n308), .A2(n2929), .A3(n3143), .Z(n3144) );
  BUFFD0 U222 ( .I(DataI[31]), .Z(n2942) );
  BUFFD0 U223 ( .I(n216), .Z(n206) );
  BUFFD0 U224 ( .I(n209), .Z(n208) );
  BUFFD0 U225 ( .I(n210), .Z(n209) );
  BUFFD0 U226 ( .I(n211), .Z(n210) );
  BUFFD0 U227 ( .I(n212), .Z(n211) );
  BUFFD0 U228 ( .I(n213), .Z(n212) );
  BUFFD0 U229 ( .I(n214), .Z(n213) );
  BUFFD0 U230 ( .I(n215), .Z(n214) );
  BUFFD0 U231 ( .I(n217), .Z(n215) );
  BUFFD0 U232 ( .I(n2942), .Z(n216) );
  BUFFD0 U233 ( .I(n206), .Z(n217) );
  BUFFD0 U234 ( .I(n2941), .Z(n218) );
  BUFFD0 U235 ( .I(n220), .Z(n219) );
  BUFFD0 U236 ( .I(n221), .Z(n220) );
  BUFFD0 U237 ( .I(n222), .Z(n221) );
  BUFFD0 U238 ( .I(n223), .Z(n222) );
  BUFFD0 U239 ( .I(n224), .Z(n223) );
  BUFFD0 U240 ( .I(n225), .Z(n224) );
  BUFFD0 U241 ( .I(n226), .Z(n225) );
  BUFFD0 U242 ( .I(n227), .Z(n226) );
  BUFFD0 U243 ( .I(n228), .Z(n227) );
  BUFFD0 U244 ( .I(n229), .Z(n228) );
  BUFFD0 U245 ( .I(n230), .Z(n229) );
  BUFFD0 U246 ( .I(n231), .Z(n230) );
  CKBD0 U247 ( .CLK(DataI[30]), .C(n2941) );
  BUFFD0 U248 ( .I(n218), .Z(n231) );
  BUFFD0 U249 ( .I(n2940), .Z(n232) );
  BUFFD0 U250 ( .I(n234), .Z(n233) );
  BUFFD0 U251 ( .I(n235), .Z(n234) );
  BUFFD0 U252 ( .I(n236), .Z(n235) );
  BUFFD0 U253 ( .I(n237), .Z(n236) );
  BUFFD0 U254 ( .I(n238), .Z(n237) );
  BUFFD0 U255 ( .I(n239), .Z(n238) );
  BUFFD0 U256 ( .I(n240), .Z(n239) );
  BUFFD0 U257 ( .I(n241), .Z(n240) );
  BUFFD0 U258 ( .I(n242), .Z(n241) );
  BUFFD0 U259 ( .I(n243), .Z(n242) );
  BUFFD0 U260 ( .I(n244), .Z(n243) );
  BUFFD0 U261 ( .I(n245), .Z(n244) );
  CKBD0 U262 ( .CLK(DataI[29]), .C(n2940) );
  BUFFD0 U263 ( .I(n232), .Z(n245) );
  BUFFD0 U264 ( .I(n248), .Z(n247) );
  BUFFD0 U265 ( .I(n249), .Z(n248) );
  BUFFD0 U266 ( .I(n250), .Z(n249) );
  BUFFD0 U267 ( .I(n251), .Z(n250) );
  BUFFD0 U268 ( .I(n252), .Z(n251) );
  BUFFD0 U269 ( .I(n253), .Z(n252) );
  BUFFD0 U270 ( .I(n254), .Z(n253) );
  BUFFD0 U271 ( .I(n255), .Z(n254) );
  BUFFD0 U272 ( .I(n257), .Z(n255) );
  BUFFD0 U273 ( .I(n2935), .Z(n256) );
  BUFFD0 U274 ( .I(n256), .Z(n257) );
  CKBD1 U275 ( .CLK(DataI[24]), .C(n2935) );
  BUFFD0 U276 ( .I(n260), .Z(n259) );
  BUFFD0 U277 ( .I(n261), .Z(n260) );
  BUFFD0 U278 ( .I(n262), .Z(n261) );
  BUFFD0 U279 ( .I(n263), .Z(n262) );
  BUFFD0 U280 ( .I(n264), .Z(n263) );
  BUFFD0 U281 ( .I(n265), .Z(n264) );
  BUFFD0 U282 ( .I(n266), .Z(n265) );
  BUFFD0 U283 ( .I(n267), .Z(n266) );
  BUFFD0 U284 ( .I(n269), .Z(n267) );
  BUFFD0 U285 ( .I(n2934), .Z(n268) );
  BUFFD0 U286 ( .I(n268), .Z(n269) );
  CKBD1 U287 ( .CLK(DataI[23]), .C(n2934) );
  BUFFD0 U288 ( .I(n272), .Z(n271) );
  BUFFD0 U289 ( .I(n273), .Z(n272) );
  BUFFD0 U290 ( .I(n274), .Z(n273) );
  BUFFD0 U291 ( .I(n275), .Z(n274) );
  BUFFD0 U292 ( .I(n276), .Z(n275) );
  BUFFD0 U293 ( .I(n277), .Z(n276) );
  BUFFD0 U294 ( .I(n278), .Z(n277) );
  BUFFD0 U295 ( .I(n279), .Z(n278) );
  BUFFD0 U296 ( .I(n280), .Z(n279) );
  CKBD0 U297 ( .CLK(DataI[22]), .C(n2933) );
  BUFFD0 U298 ( .I(n2933), .Z(n280) );
  BUFFD0 U299 ( .I(n283), .Z(n282) );
  BUFFD0 U300 ( .I(n284), .Z(n283) );
  BUFFD0 U301 ( .I(n285), .Z(n284) );
  BUFFD0 U302 ( .I(n286), .Z(n285) );
  BUFFD0 U303 ( .I(n287), .Z(n286) );
  BUFFD0 U304 ( .I(n288), .Z(n287) );
  BUFFD0 U305 ( .I(n289), .Z(n288) );
  BUFFD0 U306 ( .I(n290), .Z(n289) );
  BUFFD0 U307 ( .I(n291), .Z(n290) );
  CKBD0 U308 ( .CLK(DataI[21]), .C(n2932) );
  BUFFD0 U309 ( .I(n2932), .Z(n291) );
  BUFFD0 U310 ( .I(n294), .Z(n293) );
  BUFFD0 U311 ( .I(n295), .Z(n294) );
  BUFFD0 U312 ( .I(n296), .Z(n295) );
  BUFFD0 U313 ( .I(n297), .Z(n296) );
  BUFFD0 U314 ( .I(n298), .Z(n297) );
  BUFFD0 U315 ( .I(n299), .Z(n298) );
  BUFFD0 U316 ( .I(n300), .Z(n299) );
  BUFFD0 U317 ( .I(n301), .Z(n300) );
  BUFFD0 U318 ( .I(n303), .Z(n301) );
  BUFFD0 U319 ( .I(n2931), .Z(n302) );
  BUFFD0 U320 ( .I(n302), .Z(n303) );
  CKBD1 U321 ( .CLK(DataI[20]), .C(n2931) );
  BUFFD0 U322 ( .I(DataI[19]), .Z(n2930) );
  BUFFD0 U323 ( .I(n308), .Z(n304) );
  BUFFD0 U324 ( .I(n307), .Z(n306) );
  BUFFD0 U325 ( .I(n309), .Z(n307) );
  BUFFD0 U326 ( .I(n310), .Z(n308) );
  BUFFD0 U327 ( .I(n304), .Z(n309) );
  BUFFD0 U328 ( .I(n2930), .Z(n310) );
  BUFFD0 U329 ( .I(n313), .Z(n312) );
  BUFFD0 U330 ( .I(n314), .Z(n313) );
  BUFFD0 U331 ( .I(n315), .Z(n314) );
  BUFFD0 U332 ( .I(n316), .Z(n315) );
  BUFFD0 U333 ( .I(n317), .Z(n316) );
  BUFFD0 U334 ( .I(n318), .Z(n317) );
  BUFFD0 U335 ( .I(n319), .Z(n318) );
  BUFFD0 U336 ( .I(n320), .Z(n319) );
  BUFFD0 U337 ( .I(n321), .Z(n320) );
  CKBD0 U338 ( .CLK(DataI[18]), .C(n2929) );
  BUFFD0 U339 ( .I(n2929), .Z(n321) );
  BUFFD0 U340 ( .I(n323), .Z(n322) );
  BUFFD0 U341 ( .I(n324), .Z(n323) );
  BUFFD0 U342 ( .I(n325), .Z(n324) );
  BUFFD0 U343 ( .I(n326), .Z(n325) );
  BUFFD0 U344 ( .I(n327), .Z(n326) );
  BUFFD0 U345 ( .I(n328), .Z(n327) );
  BUFFD0 U346 ( .I(n329), .Z(n328) );
  BUFFD0 U347 ( .I(n330), .Z(n329) );
  BUFFD0 U348 ( .I(n331), .Z(n330) );
  BUFFD0 U349 ( .I(n332), .Z(n331) );
  BUFFD0 U350 ( .I(n333), .Z(n332) );
  BUFFD0 U351 ( .I(n334), .Z(n333) );
  BUFFD0 U352 ( .I(n335), .Z(n334) );
  CKBD0 U353 ( .CLK(DataI[17]), .C(n2928) );
  BUFFD0 U354 ( .I(n2928), .Z(n335) );
  BUFFD0 U355 ( .I(DataI[16]), .Z(n2927) );
  BUFFD0 U356 ( .I(n340), .Z(n336) );
  BUFFD0 U357 ( .I(n339), .Z(n338) );
  BUFFD0 U358 ( .I(n342), .Z(n339) );
  BUFFD0 U359 ( .I(n341), .Z(n340) );
  BUFFD0 U360 ( .I(n2927), .Z(n341) );
  BUFFD0 U361 ( .I(n336), .Z(n342) );
  BUFFD0 U362 ( .I(n346), .Z(n343) );
  BUFFD0 U363 ( .I(n343), .Z(n344) );
  BUFFD0 U364 ( .I(n344), .Z(n345) );
  BUFFD0 U365 ( .I(n347), .Z(n346) );
  BUFFD0 U366 ( .I(n348), .Z(n347) );
  BUFFD0 U367 ( .I(n2926), .Z(n348) );
  CKBD0 U368 ( .CLK(n345), .C(n349) );
  CKBD0 U369 ( .CLK(DataI[15]), .C(n2926) );
  BUFFD0 U370 ( .I(n353), .Z(n350) );
  BUFFD0 U371 ( .I(n350), .Z(n351) );
  BUFFD0 U372 ( .I(n351), .Z(n352) );
  BUFFD0 U373 ( .I(n354), .Z(n353) );
  BUFFD0 U374 ( .I(n355), .Z(n354) );
  BUFFD0 U375 ( .I(n2925), .Z(n355) );
  CKBD0 U376 ( .CLK(n352), .C(n356) );
  CKBD0 U377 ( .CLK(DataI[14]), .C(n2925) );
  BUFFD0 U378 ( .I(DataI[13]), .Z(n2924) );
  BUFFD0 U379 ( .I(n361), .Z(n357) );
  BUFFD0 U380 ( .I(n360), .Z(n359) );
  BUFFD0 U381 ( .I(n363), .Z(n360) );
  BUFFD0 U382 ( .I(n362), .Z(n361) );
  BUFFD0 U383 ( .I(n2924), .Z(n362) );
  BUFFD0 U384 ( .I(n357), .Z(n363) );
  BUFFD0 U385 ( .I(n370), .Z(n364) );
  BUFFD0 U386 ( .I(n366), .Z(n365) );
  BUFFD0 U387 ( .I(n367), .Z(n366) );
  BUFFD0 U388 ( .I(n368), .Z(n367) );
  BUFFD0 U389 ( .I(n369), .Z(n368) );
  BUFFD0 U390 ( .I(n371), .Z(n369) );
  BUFFD0 U391 ( .I(n372), .Z(n370) );
  BUFFD0 U392 ( .I(n373), .Z(n371) );
  BUFFD0 U393 ( .I(n2923), .Z(n372) );
  BUFFD0 U394 ( .I(n50), .Z(n373) );
  BUFFD0 U395 ( .I(n376), .Z(n374) );
  BUFFD0 U396 ( .I(n374), .Z(n375) );
  BUFFD0 U397 ( .I(n377), .Z(n376) );
  BUFFD0 U398 ( .I(n378), .Z(n377) );
  BUFFD0 U399 ( .I(n379), .Z(n378) );
  BUFFD0 U400 ( .I(n2922), .Z(n379) );
  CKBD0 U401 ( .CLK(n375), .C(n380) );
  CKBD0 U402 ( .CLK(DataI[11]), .C(n2922) );
  BUFFD0 U403 ( .I(n384), .Z(n381) );
  BUFFD0 U404 ( .I(n381), .Z(n382) );
  BUFFD0 U405 ( .I(n382), .Z(n383) );
  BUFFD0 U406 ( .I(n385), .Z(n384) );
  BUFFD0 U407 ( .I(n386), .Z(n385) );
  BUFFD0 U408 ( .I(n2921), .Z(n386) );
  CKBD0 U409 ( .CLK(n383), .C(n387) );
  CKBD0 U410 ( .CLK(DataI[10]), .C(n2921) );
  BUFFD0 U411 ( .I(n394), .Z(n388) );
  BUFFD0 U412 ( .I(n390), .Z(n389) );
  BUFFD0 U413 ( .I(n391), .Z(n390) );
  BUFFD0 U414 ( .I(n392), .Z(n391) );
  BUFFD0 U415 ( .I(n393), .Z(n392) );
  BUFFD0 U416 ( .I(n395), .Z(n393) );
  BUFFD0 U417 ( .I(n396), .Z(n394) );
  BUFFD0 U418 ( .I(n397), .Z(n395) );
  BUFFD0 U419 ( .I(n2920), .Z(n396) );
  BUFFD0 U420 ( .I(n135), .Z(n397) );
  BUFFD0 U421 ( .I(n399), .Z(n398) );
  BUFFD0 U422 ( .I(n400), .Z(n399) );
  BUFFD0 U423 ( .I(n401), .Z(n400) );
  BUFFD0 U424 ( .I(n402), .Z(n401) );
  BUFFD0 U425 ( .I(n403), .Z(n402) );
  BUFFD0 U426 ( .I(n2919), .Z(n403) );
  CKBD0 U427 ( .CLK(n398), .C(n404) );
  CKBD0 U428 ( .CLK(DataI[8]), .C(n2919) );
  BUFFD0 U429 ( .I(n406), .Z(n405) );
  BUFFD0 U430 ( .I(n407), .Z(n406) );
  BUFFD0 U431 ( .I(n408), .Z(n407) );
  BUFFD0 U432 ( .I(n409), .Z(n408) );
  BUFFD0 U433 ( .I(n410), .Z(n409) );
  BUFFD0 U434 ( .I(n2918), .Z(n410) );
  CKBD0 U435 ( .CLK(n405), .C(n411) );
  CKBD0 U436 ( .CLK(DataI[7]), .C(n2918) );
  BUFFD0 U437 ( .I(n418), .Z(n412) );
  BUFFD0 U438 ( .I(n414), .Z(n413) );
  BUFFD0 U439 ( .I(n415), .Z(n414) );
  BUFFD0 U440 ( .I(n416), .Z(n415) );
  BUFFD0 U441 ( .I(n417), .Z(n416) );
  BUFFD0 U442 ( .I(n419), .Z(n417) );
  BUFFD0 U443 ( .I(n420), .Z(n418) );
  BUFFD0 U444 ( .I(n421), .Z(n419) );
  BUFFD0 U445 ( .I(n2917), .Z(n420) );
  BUFFD0 U446 ( .I(n412), .Z(n421) );
  BUFFD0 U447 ( .I(DataI[5]), .Z(n423) );
  CKBD0 U448 ( .CLK(n200), .C(n424) );
  CKBD0 U449 ( .CLK(DataI[4]), .C(n2916) );
  BUFFD0 U450 ( .I(n426), .Z(n425) );
  BUFFD0 U451 ( .I(n427), .Z(n426) );
  BUFFD0 U452 ( .I(n428), .Z(n427) );
  BUFFD0 U453 ( .I(n429), .Z(n428) );
  BUFFD0 U454 ( .I(n2915), .Z(n429) );
  CKBD0 U455 ( .CLK(n201), .C(n430) );
  CKBD0 U456 ( .CLK(DataI[3]), .C(n2915) );
  BUFFD0 U457 ( .I(DataI[2]), .Z(n432) );
  BUFFD0 U458 ( .I(DataI[0]), .Z(n435) );
  BUFFD0 U459 ( .I(n440), .Z(n436) );
  BUFFD0 U460 ( .I(n3116), .Z(n437) );
  BUFFD0 U461 ( .I(n437), .Z(n438) );
  BUFFD0 U462 ( .I(n438), .Z(n439) );
  BUFFD0 U463 ( .I(n441), .Z(n440) );
  BUFFD0 U464 ( .I(n442), .Z(n441) );
  BUFFD0 U465 ( .I(n443), .Z(n442) );
  BUFFD0 U466 ( .I(n444), .Z(n443) );
  BUFFD0 U467 ( .I(n445), .Z(n444) );
  BUFFD0 U468 ( .I(n446), .Z(n445) );
  BUFFD0 U469 ( .I(n447), .Z(n446) );
  BUFFD0 U470 ( .I(n448), .Z(n447) );
  BUFFD0 U471 ( .I(n449), .Z(n448) );
  BUFFD0 U472 ( .I(n450), .Z(n449) );
  BUFFD0 U473 ( .I(n451), .Z(n450) );
  BUFFD0 U474 ( .I(n452), .Z(n451) );
  BUFFD0 U475 ( .I(n453), .Z(n452) );
  BUFFD0 U476 ( .I(n454), .Z(n453) );
  BUFFD0 U477 ( .I(n455), .Z(n454) );
  BUFFD0 U478 ( .I(n456), .Z(n455) );
  BUFFD0 U479 ( .I(n457), .Z(n456) );
  BUFFD0 U480 ( .I(n458), .Z(n457) );
  BUFFD0 U481 ( .I(n459), .Z(n458) );
  BUFFD0 U482 ( .I(n460), .Z(n459) );
  BUFFD0 U483 ( .I(n461), .Z(n460) );
  BUFFD0 U484 ( .I(n462), .Z(n461) );
  BUFFD0 U485 ( .I(n463), .Z(n462) );
  BUFFD0 U486 ( .I(n464), .Z(n463) );
  BUFFD0 U487 ( .I(n465), .Z(n464) );
  BUFFD0 U488 ( .I(n466), .Z(n465) );
  BUFFD0 U489 ( .I(n467), .Z(n466) );
  BUFFD0 U490 ( .I(n468), .Z(n467) );
  BUFFD0 U491 ( .I(n469), .Z(n468) );
  BUFFD0 U492 ( .I(n470), .Z(n469) );
  BUFFD0 U493 ( .I(n471), .Z(n470) );
  BUFFD0 U494 ( .I(n472), .Z(n471) );
  BUFFD0 U495 ( .I(n473), .Z(n472) );
  BUFFD0 U496 ( .I(n474), .Z(n473) );
  BUFFD0 U497 ( .I(n475), .Z(n474) );
  BUFFD0 U498 ( .I(n476), .Z(n475) );
  BUFFD0 U499 ( .I(n477), .Z(n476) );
  BUFFD0 U500 ( .I(n478), .Z(n477) );
  BUFFD0 U501 ( .I(n479), .Z(n478) );
  BUFFD0 U502 ( .I(n480), .Z(n479) );
  BUFFD0 U503 ( .I(n481), .Z(n480) );
  BUFFD0 U504 ( .I(n482), .Z(n481) );
  BUFFD0 U505 ( .I(n483), .Z(n482) );
  BUFFD0 U506 ( .I(n484), .Z(n483) );
  BUFFD0 U507 ( .I(n485), .Z(n484) );
  BUFFD0 U508 ( .I(n486), .Z(n485) );
  BUFFD0 U509 ( .I(n487), .Z(n486) );
  BUFFD0 U510 ( .I(n488), .Z(n487) );
  BUFFD0 U511 ( .I(n489), .Z(n488) );
  BUFFD0 U512 ( .I(n490), .Z(n489) );
  BUFFD0 U513 ( .I(n491), .Z(n490) );
  BUFFD0 U514 ( .I(n492), .Z(n491) );
  BUFFD0 U515 ( .I(n493), .Z(n492) );
  BUFFD0 U516 ( .I(n494), .Z(n493) );
  BUFFD0 U517 ( .I(n496), .Z(n494) );
  BUFFD0 U518 ( .I(n498), .Z(n495) );
  BUFFD0 U519 ( .I(n497), .Z(n496) );
  BUFFD0 U520 ( .I(n439), .Z(n497) );
  BUFFD0 U521 ( .I(Dreadyr), .Z(n498) );
  OR2D0 U522 ( .A1(n2713), .A2(n495), .Z(n3116) );
  BUFFD0 U523 ( .I(DataI[28]), .Z(n2939) );
  BUFFD0 U524 ( .I(n509), .Z(n499) );
  BUFFD0 U525 ( .I(n502), .Z(n501) );
  BUFFD0 U526 ( .I(n503), .Z(n502) );
  BUFFD0 U527 ( .I(n504), .Z(n503) );
  BUFFD0 U528 ( .I(n505), .Z(n504) );
  BUFFD0 U529 ( .I(n506), .Z(n505) );
  BUFFD0 U530 ( .I(n507), .Z(n506) );
  BUFFD0 U531 ( .I(n508), .Z(n507) );
  BUFFD0 U532 ( .I(n510), .Z(n508) );
  BUFFD0 U533 ( .I(n2939), .Z(n509) );
  BUFFD0 U534 ( .I(n499), .Z(n510) );
  CKBXD0 U535 ( .I(n512), .Z(n511) );
  CKBXD0 U536 ( .I(n2938), .Z(n512) );
  CKBXD0 U537 ( .I(DataI[27]), .Z(n2938) );
  BUFFD0 U538 ( .I(n2937), .Z(n513) );
  BUFFD0 U539 ( .I(n515), .Z(n514) );
  BUFFD0 U540 ( .I(n516), .Z(n515) );
  BUFFD0 U541 ( .I(n517), .Z(n516) );
  BUFFD0 U542 ( .I(n518), .Z(n517) );
  BUFFD0 U543 ( .I(n519), .Z(n518) );
  BUFFD0 U544 ( .I(n520), .Z(n519) );
  BUFFD0 U545 ( .I(n521), .Z(n520) );
  BUFFD0 U546 ( .I(n522), .Z(n521) );
  BUFFD0 U547 ( .I(n523), .Z(n522) );
  BUFFD0 U548 ( .I(n524), .Z(n523) );
  BUFFD0 U549 ( .I(n525), .Z(n524) );
  BUFFD0 U550 ( .I(n526), .Z(n525) );
  CKBD0 U551 ( .CLK(DataI[26]), .C(n2937) );
  BUFFD0 U552 ( .I(n513), .Z(n526) );
  CKBXD0 U553 ( .I(n528), .Z(n527) );
  CKBXD0 U554 ( .I(n2936), .Z(n528) );
  CKBXD0 U555 ( .I(DataI[25]), .Z(n2936) );
  BUFFD0 U556 ( .I(n532), .Z(n529) );
  BUFFD0 U557 ( .I(n530), .Z(n531) );
  BUFFD0 U558 ( .I(n533), .Z(n532) );
  BUFFD0 U559 ( .I(n534), .Z(n533) );
  BUFFD0 U560 ( .I(n535), .Z(n534) );
  BUFFD0 U561 ( .I(n536), .Z(n535) );
  BUFFD0 U562 ( .I(n537), .Z(n536) );
  BUFFD0 U563 ( .I(n538), .Z(n537) );
  BUFFD0 U564 ( .I(n539), .Z(n538) );
  BUFFD0 U565 ( .I(n540), .Z(n539) );
  BUFFD0 U566 ( .I(n541), .Z(n540) );
  BUFFD0 U567 ( .I(n542), .Z(n541) );
  BUFFD0 U568 ( .I(n543), .Z(n542) );
  BUFFD0 U569 ( .I(n544), .Z(n543) );
  BUFFD0 U570 ( .I(n545), .Z(n544) );
  BUFFD0 U571 ( .I(n546), .Z(n545) );
  BUFFD0 U572 ( .I(n547), .Z(n546) );
  BUFFD0 U573 ( .I(n548), .Z(n547) );
  BUFFD0 U574 ( .I(n549), .Z(n548) );
  BUFFD0 U575 ( .I(n550), .Z(n549) );
  BUFFD0 U576 ( .I(n551), .Z(n550) );
  BUFFD0 U577 ( .I(n552), .Z(n551) );
  BUFFD0 U578 ( .I(n553), .Z(n552) );
  BUFFD0 U579 ( .I(n554), .Z(n553) );
  BUFFD0 U580 ( .I(n555), .Z(n554) );
  BUFFD0 U581 ( .I(n556), .Z(n555) );
  BUFFD0 U582 ( .I(n557), .Z(n556) );
  BUFFD0 U583 ( .I(n558), .Z(n557) );
  BUFFD0 U584 ( .I(n559), .Z(n558) );
  BUFFD0 U585 ( .I(n560), .Z(n559) );
  BUFFD0 U586 ( .I(n561), .Z(n560) );
  BUFFD0 U587 ( .I(n562), .Z(n561) );
  BUFFD0 U588 ( .I(n563), .Z(n562) );
  BUFFD0 U589 ( .I(n564), .Z(n563) );
  BUFFD0 U590 ( .I(n565), .Z(n564) );
  BUFFD0 U591 ( .I(n566), .Z(n565) );
  BUFFD0 U592 ( .I(n567), .Z(n566) );
  BUFFD0 U593 ( .I(n568), .Z(n567) );
  BUFFD0 U594 ( .I(n569), .Z(n568) );
  BUFFD0 U595 ( .I(n570), .Z(n569) );
  BUFFD0 U596 ( .I(n571), .Z(n570) );
  BUFFD0 U597 ( .I(n572), .Z(n571) );
  BUFFD0 U598 ( .I(n573), .Z(n572) );
  BUFFD0 U599 ( .I(n574), .Z(n573) );
  BUFFD0 U600 ( .I(n575), .Z(n574) );
  BUFFD0 U601 ( .I(n576), .Z(n575) );
  BUFFD0 U602 ( .I(n577), .Z(n576) );
  BUFFD0 U603 ( .I(n578), .Z(n577) );
  BUFFD0 U604 ( .I(n579), .Z(n578) );
  BUFFD0 U605 ( .I(n580), .Z(n579) );
  BUFFD0 U606 ( .I(n581), .Z(n580) );
  BUFFD0 U607 ( .I(n582), .Z(n581) );
  BUFFD0 U608 ( .I(n583), .Z(n582) );
  BUFFD0 U609 ( .I(n584), .Z(n583) );
  BUFFD0 U610 ( .I(n585), .Z(n584) );
  BUFFD0 U611 ( .I(n586), .Z(n585) );
  BUFFD0 U612 ( .I(n587), .Z(n586) );
  BUFFD0 U613 ( .I(n588), .Z(n587) );
  BUFFD0 U614 ( .I(n589), .Z(n588) );
  BUFFD0 U615 ( .I(n590), .Z(n589) );
  BUFFD0 U616 ( .I(n591), .Z(n590) );
  BUFFD0 U617 ( .I(n592), .Z(n591) );
  BUFFD0 U618 ( .I(n593), .Z(n592) );
  BUFFD0 U619 ( .I(n594), .Z(n593) );
  BUFFD0 U620 ( .I(n531), .Z(n594) );
  BUFFD0 U621 ( .I(n598), .Z(n595) );
  BUFFD0 U622 ( .I(n596), .Z(n597) );
  BUFFD0 U623 ( .I(n599), .Z(n598) );
  BUFFD0 U624 ( .I(n600), .Z(n599) );
  BUFFD0 U625 ( .I(n601), .Z(n600) );
  BUFFD0 U626 ( .I(n602), .Z(n601) );
  BUFFD0 U627 ( .I(n603), .Z(n602) );
  BUFFD0 U628 ( .I(n604), .Z(n603) );
  BUFFD0 U629 ( .I(n605), .Z(n604) );
  BUFFD0 U630 ( .I(n606), .Z(n605) );
  BUFFD0 U631 ( .I(n607), .Z(n606) );
  BUFFD0 U632 ( .I(n608), .Z(n607) );
  BUFFD0 U633 ( .I(n609), .Z(n608) );
  BUFFD0 U634 ( .I(n610), .Z(n609) );
  BUFFD0 U635 ( .I(n611), .Z(n610) );
  BUFFD0 U636 ( .I(n612), .Z(n611) );
  BUFFD0 U637 ( .I(n613), .Z(n612) );
  BUFFD0 U638 ( .I(n614), .Z(n613) );
  BUFFD0 U639 ( .I(n615), .Z(n614) );
  BUFFD0 U640 ( .I(n616), .Z(n615) );
  BUFFD0 U641 ( .I(n617), .Z(n616) );
  BUFFD0 U642 ( .I(n618), .Z(n617) );
  BUFFD0 U643 ( .I(n619), .Z(n618) );
  BUFFD0 U644 ( .I(n620), .Z(n619) );
  BUFFD0 U645 ( .I(n621), .Z(n620) );
  BUFFD0 U646 ( .I(n622), .Z(n621) );
  BUFFD0 U647 ( .I(n623), .Z(n622) );
  BUFFD0 U648 ( .I(n624), .Z(n623) );
  BUFFD0 U649 ( .I(n625), .Z(n624) );
  BUFFD0 U650 ( .I(n626), .Z(n625) );
  BUFFD0 U651 ( .I(n627), .Z(n626) );
  BUFFD0 U652 ( .I(n628), .Z(n627) );
  BUFFD0 U653 ( .I(n629), .Z(n628) );
  BUFFD0 U654 ( .I(n630), .Z(n629) );
  BUFFD0 U655 ( .I(n631), .Z(n630) );
  BUFFD0 U656 ( .I(n632), .Z(n631) );
  BUFFD0 U657 ( .I(n633), .Z(n632) );
  BUFFD0 U658 ( .I(n634), .Z(n633) );
  BUFFD0 U659 ( .I(n635), .Z(n634) );
  BUFFD0 U660 ( .I(n636), .Z(n635) );
  BUFFD0 U661 ( .I(n637), .Z(n636) );
  BUFFD0 U662 ( .I(n638), .Z(n637) );
  BUFFD0 U663 ( .I(n639), .Z(n638) );
  BUFFD0 U664 ( .I(n640), .Z(n639) );
  BUFFD0 U665 ( .I(n641), .Z(n640) );
  BUFFD0 U666 ( .I(n642), .Z(n641) );
  BUFFD0 U667 ( .I(n643), .Z(n642) );
  BUFFD0 U668 ( .I(n644), .Z(n643) );
  BUFFD0 U669 ( .I(n645), .Z(n644) );
  BUFFD0 U670 ( .I(n646), .Z(n645) );
  BUFFD0 U671 ( .I(n647), .Z(n646) );
  BUFFD0 U672 ( .I(n648), .Z(n647) );
  BUFFD0 U673 ( .I(n649), .Z(n648) );
  BUFFD0 U674 ( .I(n650), .Z(n649) );
  BUFFD0 U675 ( .I(n651), .Z(n650) );
  BUFFD0 U676 ( .I(n652), .Z(n651) );
  BUFFD0 U677 ( .I(n653), .Z(n652) );
  BUFFD0 U678 ( .I(n654), .Z(n653) );
  BUFFD0 U679 ( .I(n655), .Z(n654) );
  BUFFD0 U680 ( .I(n656), .Z(n655) );
  BUFFD0 U681 ( .I(n657), .Z(n656) );
  BUFFD0 U682 ( .I(n658), .Z(n657) );
  BUFFD0 U683 ( .I(n659), .Z(n658) );
  BUFFD0 U684 ( .I(n660), .Z(n659) );
  BUFFD0 U685 ( .I(n597), .Z(n660) );
  CKBD0 U686 ( .CLK(N52), .C(n662) );
  BUFFD0 U687 ( .I(n664), .Z(n661) );
  BUFFD0 U688 ( .I(n662), .Z(n663) );
  BUFFD0 U689 ( .I(n665), .Z(n664) );
  BUFFD0 U690 ( .I(n666), .Z(n665) );
  BUFFD0 U691 ( .I(n667), .Z(n666) );
  BUFFD0 U692 ( .I(n668), .Z(n667) );
  BUFFD0 U693 ( .I(n669), .Z(n668) );
  BUFFD0 U694 ( .I(n670), .Z(n669) );
  BUFFD0 U695 ( .I(n671), .Z(n670) );
  BUFFD0 U696 ( .I(n672), .Z(n671) );
  BUFFD0 U697 ( .I(n673), .Z(n672) );
  BUFFD0 U698 ( .I(n674), .Z(n673) );
  BUFFD0 U699 ( .I(n675), .Z(n674) );
  BUFFD0 U700 ( .I(n676), .Z(n675) );
  BUFFD0 U701 ( .I(n677), .Z(n676) );
  BUFFD0 U702 ( .I(n678), .Z(n677) );
  BUFFD0 U703 ( .I(n679), .Z(n678) );
  BUFFD0 U704 ( .I(n680), .Z(n679) );
  BUFFD0 U705 ( .I(n681), .Z(n680) );
  BUFFD0 U706 ( .I(n682), .Z(n681) );
  BUFFD0 U707 ( .I(n683), .Z(n682) );
  BUFFD0 U708 ( .I(n684), .Z(n683) );
  BUFFD0 U709 ( .I(n685), .Z(n684) );
  BUFFD0 U710 ( .I(n686), .Z(n685) );
  BUFFD0 U711 ( .I(n687), .Z(n686) );
  BUFFD0 U712 ( .I(n688), .Z(n687) );
  BUFFD0 U713 ( .I(n689), .Z(n688) );
  BUFFD0 U714 ( .I(n690), .Z(n689) );
  BUFFD0 U715 ( .I(n691), .Z(n690) );
  BUFFD0 U716 ( .I(n692), .Z(n691) );
  BUFFD0 U717 ( .I(n693), .Z(n692) );
  BUFFD0 U718 ( .I(n694), .Z(n693) );
  BUFFD0 U719 ( .I(n695), .Z(n694) );
  BUFFD0 U720 ( .I(n696), .Z(n695) );
  BUFFD0 U721 ( .I(n697), .Z(n696) );
  BUFFD0 U722 ( .I(n698), .Z(n697) );
  BUFFD0 U723 ( .I(n699), .Z(n698) );
  BUFFD0 U724 ( .I(n700), .Z(n699) );
  BUFFD0 U725 ( .I(n701), .Z(n700) );
  BUFFD0 U726 ( .I(n702), .Z(n701) );
  BUFFD0 U727 ( .I(n703), .Z(n702) );
  BUFFD0 U728 ( .I(n704), .Z(n703) );
  BUFFD0 U729 ( .I(n705), .Z(n704) );
  BUFFD0 U730 ( .I(n706), .Z(n705) );
  BUFFD0 U731 ( .I(n707), .Z(n706) );
  BUFFD0 U732 ( .I(n708), .Z(n707) );
  BUFFD0 U733 ( .I(n709), .Z(n708) );
  BUFFD0 U734 ( .I(n710), .Z(n709) );
  BUFFD0 U735 ( .I(n711), .Z(n710) );
  BUFFD0 U736 ( .I(n712), .Z(n711) );
  BUFFD0 U737 ( .I(n713), .Z(n712) );
  BUFFD0 U738 ( .I(n714), .Z(n713) );
  BUFFD0 U739 ( .I(n715), .Z(n714) );
  BUFFD0 U740 ( .I(n716), .Z(n715) );
  BUFFD0 U741 ( .I(n717), .Z(n716) );
  BUFFD0 U742 ( .I(n718), .Z(n717) );
  BUFFD0 U743 ( .I(n719), .Z(n718) );
  BUFFD0 U744 ( .I(n720), .Z(n719) );
  BUFFD0 U745 ( .I(n721), .Z(n720) );
  BUFFD0 U746 ( .I(n722), .Z(n721) );
  BUFFD0 U747 ( .I(n723), .Z(n722) );
  BUFFD0 U748 ( .I(n724), .Z(n723) );
  BUFFD0 U749 ( .I(n725), .Z(n724) );
  BUFFD0 U750 ( .I(n726), .Z(n725) );
  BUFFD0 U751 ( .I(n663), .Z(n726) );
  CKBD0 U752 ( .CLK(N53), .C(n728) );
  BUFFD0 U753 ( .I(n730), .Z(n727) );
  BUFFD0 U754 ( .I(n728), .Z(n729) );
  BUFFD0 U755 ( .I(n731), .Z(n730) );
  BUFFD0 U756 ( .I(n732), .Z(n731) );
  BUFFD0 U757 ( .I(n733), .Z(n732) );
  BUFFD0 U758 ( .I(n734), .Z(n733) );
  BUFFD0 U759 ( .I(n735), .Z(n734) );
  BUFFD0 U760 ( .I(n736), .Z(n735) );
  BUFFD0 U761 ( .I(n737), .Z(n736) );
  BUFFD0 U762 ( .I(n738), .Z(n737) );
  BUFFD0 U763 ( .I(n739), .Z(n738) );
  BUFFD0 U764 ( .I(n740), .Z(n739) );
  BUFFD0 U765 ( .I(n741), .Z(n740) );
  BUFFD0 U766 ( .I(n742), .Z(n741) );
  BUFFD0 U767 ( .I(n743), .Z(n742) );
  BUFFD0 U768 ( .I(n744), .Z(n743) );
  BUFFD0 U769 ( .I(n745), .Z(n744) );
  BUFFD0 U770 ( .I(n746), .Z(n745) );
  BUFFD0 U771 ( .I(n747), .Z(n746) );
  BUFFD0 U772 ( .I(n748), .Z(n747) );
  BUFFD0 U773 ( .I(n749), .Z(n748) );
  BUFFD0 U774 ( .I(n750), .Z(n749) );
  BUFFD0 U775 ( .I(n751), .Z(n750) );
  BUFFD0 U776 ( .I(n752), .Z(n751) );
  BUFFD0 U777 ( .I(n753), .Z(n752) );
  BUFFD0 U778 ( .I(n754), .Z(n753) );
  BUFFD0 U779 ( .I(n755), .Z(n754) );
  BUFFD0 U780 ( .I(n756), .Z(n755) );
  BUFFD0 U781 ( .I(n757), .Z(n756) );
  BUFFD0 U782 ( .I(n758), .Z(n757) );
  BUFFD0 U783 ( .I(n759), .Z(n758) );
  BUFFD0 U784 ( .I(n760), .Z(n759) );
  BUFFD0 U785 ( .I(n761), .Z(n760) );
  BUFFD0 U786 ( .I(n762), .Z(n761) );
  BUFFD0 U787 ( .I(n763), .Z(n762) );
  BUFFD0 U788 ( .I(n764), .Z(n763) );
  BUFFD0 U789 ( .I(n765), .Z(n764) );
  BUFFD0 U790 ( .I(n766), .Z(n765) );
  BUFFD0 U791 ( .I(n767), .Z(n766) );
  BUFFD0 U792 ( .I(n768), .Z(n767) );
  BUFFD0 U793 ( .I(n769), .Z(n768) );
  BUFFD0 U794 ( .I(n770), .Z(n769) );
  BUFFD0 U795 ( .I(n771), .Z(n770) );
  BUFFD0 U796 ( .I(n772), .Z(n771) );
  BUFFD0 U797 ( .I(n773), .Z(n772) );
  BUFFD0 U798 ( .I(n774), .Z(n773) );
  BUFFD0 U799 ( .I(n775), .Z(n774) );
  BUFFD0 U800 ( .I(n776), .Z(n775) );
  BUFFD0 U801 ( .I(n777), .Z(n776) );
  BUFFD0 U802 ( .I(n778), .Z(n777) );
  BUFFD0 U803 ( .I(n779), .Z(n778) );
  BUFFD0 U804 ( .I(n780), .Z(n779) );
  BUFFD0 U805 ( .I(n781), .Z(n780) );
  BUFFD0 U806 ( .I(n782), .Z(n781) );
  BUFFD0 U807 ( .I(n783), .Z(n782) );
  BUFFD0 U808 ( .I(n784), .Z(n783) );
  BUFFD0 U809 ( .I(n785), .Z(n784) );
  BUFFD0 U810 ( .I(n786), .Z(n785) );
  BUFFD0 U811 ( .I(n787), .Z(n786) );
  BUFFD0 U812 ( .I(n788), .Z(n787) );
  BUFFD0 U813 ( .I(n789), .Z(n788) );
  BUFFD0 U814 ( .I(n790), .Z(n789) );
  BUFFD0 U815 ( .I(n791), .Z(n790) );
  BUFFD0 U816 ( .I(n792), .Z(n791) );
  BUFFD0 U817 ( .I(n729), .Z(n792) );
  BUFFD0 U818 ( .I(n796), .Z(n793) );
  BUFFD0 U819 ( .I(N54), .Z(n794) );
  BUFFD0 U820 ( .I(n794), .Z(n795) );
  BUFFD0 U821 ( .I(n797), .Z(n796) );
  BUFFD0 U822 ( .I(n798), .Z(n797) );
  BUFFD0 U823 ( .I(n799), .Z(n798) );
  BUFFD0 U824 ( .I(n800), .Z(n799) );
  BUFFD0 U825 ( .I(n801), .Z(n800) );
  BUFFD0 U826 ( .I(n802), .Z(n801) );
  BUFFD0 U827 ( .I(n803), .Z(n802) );
  BUFFD0 U828 ( .I(n804), .Z(n803) );
  BUFFD0 U829 ( .I(n805), .Z(n804) );
  BUFFD0 U830 ( .I(n806), .Z(n805) );
  BUFFD0 U831 ( .I(n807), .Z(n806) );
  BUFFD0 U832 ( .I(n808), .Z(n807) );
  BUFFD0 U833 ( .I(n809), .Z(n808) );
  BUFFD0 U834 ( .I(n810), .Z(n809) );
  BUFFD0 U835 ( .I(n811), .Z(n810) );
  BUFFD0 U836 ( .I(n812), .Z(n811) );
  BUFFD0 U837 ( .I(n813), .Z(n812) );
  BUFFD0 U838 ( .I(n814), .Z(n813) );
  BUFFD0 U839 ( .I(n815), .Z(n814) );
  BUFFD0 U840 ( .I(n816), .Z(n815) );
  BUFFD0 U841 ( .I(n817), .Z(n816) );
  BUFFD0 U842 ( .I(n818), .Z(n817) );
  BUFFD0 U843 ( .I(n819), .Z(n818) );
  BUFFD0 U844 ( .I(n820), .Z(n819) );
  BUFFD0 U845 ( .I(n821), .Z(n820) );
  BUFFD0 U846 ( .I(n822), .Z(n821) );
  BUFFD0 U847 ( .I(n823), .Z(n822) );
  BUFFD0 U848 ( .I(n824), .Z(n823) );
  BUFFD0 U849 ( .I(n825), .Z(n824) );
  BUFFD0 U850 ( .I(n826), .Z(n825) );
  BUFFD0 U851 ( .I(n827), .Z(n826) );
  BUFFD0 U852 ( .I(n828), .Z(n827) );
  BUFFD0 U853 ( .I(n829), .Z(n828) );
  BUFFD0 U854 ( .I(n830), .Z(n829) );
  BUFFD0 U855 ( .I(n831), .Z(n830) );
  BUFFD0 U856 ( .I(n832), .Z(n831) );
  BUFFD0 U857 ( .I(n833), .Z(n832) );
  BUFFD0 U858 ( .I(n834), .Z(n833) );
  BUFFD0 U859 ( .I(n835), .Z(n834) );
  BUFFD0 U860 ( .I(n836), .Z(n835) );
  BUFFD0 U861 ( .I(n837), .Z(n836) );
  BUFFD0 U862 ( .I(n838), .Z(n837) );
  BUFFD0 U863 ( .I(n839), .Z(n838) );
  BUFFD0 U864 ( .I(n840), .Z(n839) );
  BUFFD0 U865 ( .I(n841), .Z(n840) );
  BUFFD0 U866 ( .I(n842), .Z(n841) );
  BUFFD0 U867 ( .I(n843), .Z(n842) );
  BUFFD0 U868 ( .I(n844), .Z(n843) );
  BUFFD0 U869 ( .I(n845), .Z(n844) );
  BUFFD0 U870 ( .I(n846), .Z(n845) );
  BUFFD0 U871 ( .I(n847), .Z(n846) );
  BUFFD0 U872 ( .I(n848), .Z(n847) );
  BUFFD0 U873 ( .I(n849), .Z(n848) );
  BUFFD0 U874 ( .I(n850), .Z(n849) );
  BUFFD0 U875 ( .I(n851), .Z(n850) );
  BUFFD0 U876 ( .I(n852), .Z(n851) );
  BUFFD0 U877 ( .I(n853), .Z(n852) );
  BUFFD0 U878 ( .I(n854), .Z(n853) );
  BUFFD0 U879 ( .I(n855), .Z(n854) );
  BUFFD0 U880 ( .I(n856), .Z(n855) );
  BUFFD0 U881 ( .I(n857), .Z(n856) );
  BUFFD0 U882 ( .I(n858), .Z(n857) );
  BUFFD0 U883 ( .I(n795), .Z(n858) );
  BUFFD0 U884 ( .I(n862), .Z(n859) );
  BUFFD0 U885 ( .I(n860), .Z(n861) );
  BUFFD0 U886 ( .I(n863), .Z(n862) );
  BUFFD0 U887 ( .I(n864), .Z(n863) );
  BUFFD0 U888 ( .I(n865), .Z(n864) );
  BUFFD0 U889 ( .I(n866), .Z(n865) );
  BUFFD0 U890 ( .I(n867), .Z(n866) );
  BUFFD0 U891 ( .I(n868), .Z(n867) );
  BUFFD0 U892 ( .I(n869), .Z(n868) );
  BUFFD0 U893 ( .I(n870), .Z(n869) );
  BUFFD0 U894 ( .I(n871), .Z(n870) );
  BUFFD0 U895 ( .I(n872), .Z(n871) );
  BUFFD0 U896 ( .I(n873), .Z(n872) );
  BUFFD0 U897 ( .I(n874), .Z(n873) );
  BUFFD0 U898 ( .I(n875), .Z(n874) );
  BUFFD0 U899 ( .I(n876), .Z(n875) );
  BUFFD0 U900 ( .I(n877), .Z(n876) );
  BUFFD0 U901 ( .I(n878), .Z(n877) );
  BUFFD0 U902 ( .I(n879), .Z(n878) );
  BUFFD0 U903 ( .I(n880), .Z(n879) );
  BUFFD0 U904 ( .I(n881), .Z(n880) );
  BUFFD0 U905 ( .I(n882), .Z(n881) );
  BUFFD0 U906 ( .I(n883), .Z(n882) );
  BUFFD0 U907 ( .I(n884), .Z(n883) );
  BUFFD0 U908 ( .I(n885), .Z(n884) );
  BUFFD0 U909 ( .I(n886), .Z(n885) );
  BUFFD0 U910 ( .I(n887), .Z(n886) );
  BUFFD0 U911 ( .I(n888), .Z(n887) );
  BUFFD0 U912 ( .I(n889), .Z(n888) );
  BUFFD0 U913 ( .I(n890), .Z(n889) );
  BUFFD0 U914 ( .I(n891), .Z(n890) );
  BUFFD0 U915 ( .I(n892), .Z(n891) );
  BUFFD0 U916 ( .I(n893), .Z(n892) );
  BUFFD0 U917 ( .I(n894), .Z(n893) );
  BUFFD0 U918 ( .I(n895), .Z(n894) );
  BUFFD0 U919 ( .I(n896), .Z(n895) );
  BUFFD0 U920 ( .I(n897), .Z(n896) );
  BUFFD0 U921 ( .I(n898), .Z(n897) );
  BUFFD0 U922 ( .I(n899), .Z(n898) );
  BUFFD0 U923 ( .I(n900), .Z(n899) );
  BUFFD0 U924 ( .I(n901), .Z(n900) );
  BUFFD0 U925 ( .I(n902), .Z(n901) );
  BUFFD0 U926 ( .I(n903), .Z(n902) );
  BUFFD0 U927 ( .I(n904), .Z(n903) );
  BUFFD0 U928 ( .I(n905), .Z(n904) );
  BUFFD0 U929 ( .I(n906), .Z(n905) );
  BUFFD0 U930 ( .I(n907), .Z(n906) );
  BUFFD0 U931 ( .I(n908), .Z(n907) );
  BUFFD0 U932 ( .I(n909), .Z(n908) );
  BUFFD0 U933 ( .I(n910), .Z(n909) );
  BUFFD0 U934 ( .I(n911), .Z(n910) );
  BUFFD0 U935 ( .I(n912), .Z(n911) );
  BUFFD0 U936 ( .I(n913), .Z(n912) );
  BUFFD0 U937 ( .I(n914), .Z(n913) );
  BUFFD0 U938 ( .I(n915), .Z(n914) );
  BUFFD0 U939 ( .I(n916), .Z(n915) );
  BUFFD0 U940 ( .I(n917), .Z(n916) );
  BUFFD0 U941 ( .I(n918), .Z(n917) );
  BUFFD0 U942 ( .I(n919), .Z(n918) );
  BUFFD0 U943 ( .I(n920), .Z(n919) );
  BUFFD0 U944 ( .I(n921), .Z(n920) );
  BUFFD0 U945 ( .I(n922), .Z(n921) );
  BUFFD0 U946 ( .I(n923), .Z(n922) );
  BUFFD0 U947 ( .I(n924), .Z(n923) );
  BUFFD0 U948 ( .I(n861), .Z(n924) );
  CKBD0 U949 ( .CLK(N56), .C(n926) );
  BUFFD0 U950 ( .I(n928), .Z(n925) );
  BUFFD0 U951 ( .I(n926), .Z(n927) );
  BUFFD0 U952 ( .I(n929), .Z(n928) );
  BUFFD0 U953 ( .I(n930), .Z(n929) );
  BUFFD0 U954 ( .I(n931), .Z(n930) );
  BUFFD0 U955 ( .I(n932), .Z(n931) );
  BUFFD0 U956 ( .I(n933), .Z(n932) );
  BUFFD0 U957 ( .I(n934), .Z(n933) );
  BUFFD0 U958 ( .I(n935), .Z(n934) );
  BUFFD0 U959 ( .I(n936), .Z(n935) );
  BUFFD0 U960 ( .I(n937), .Z(n936) );
  BUFFD0 U961 ( .I(n938), .Z(n937) );
  BUFFD0 U962 ( .I(n939), .Z(n938) );
  BUFFD0 U963 ( .I(n940), .Z(n939) );
  BUFFD0 U964 ( .I(n941), .Z(n940) );
  BUFFD0 U965 ( .I(n942), .Z(n941) );
  BUFFD0 U966 ( .I(n943), .Z(n942) );
  BUFFD0 U967 ( .I(n944), .Z(n943) );
  BUFFD0 U968 ( .I(n945), .Z(n944) );
  BUFFD0 U969 ( .I(n946), .Z(n945) );
  BUFFD0 U970 ( .I(n947), .Z(n946) );
  BUFFD0 U971 ( .I(n948), .Z(n947) );
  BUFFD0 U972 ( .I(n949), .Z(n948) );
  BUFFD0 U973 ( .I(n950), .Z(n949) );
  BUFFD0 U974 ( .I(n951), .Z(n950) );
  BUFFD0 U975 ( .I(n952), .Z(n951) );
  BUFFD0 U976 ( .I(n953), .Z(n952) );
  BUFFD0 U977 ( .I(n954), .Z(n953) );
  BUFFD0 U978 ( .I(n955), .Z(n954) );
  BUFFD0 U979 ( .I(n956), .Z(n955) );
  BUFFD0 U980 ( .I(n957), .Z(n956) );
  BUFFD0 U981 ( .I(n958), .Z(n957) );
  BUFFD0 U982 ( .I(n959), .Z(n958) );
  BUFFD0 U983 ( .I(n960), .Z(n959) );
  BUFFD0 U984 ( .I(n961), .Z(n960) );
  BUFFD0 U985 ( .I(n962), .Z(n961) );
  BUFFD0 U986 ( .I(n963), .Z(n962) );
  BUFFD0 U987 ( .I(n964), .Z(n963) );
  BUFFD0 U988 ( .I(n965), .Z(n964) );
  BUFFD0 U989 ( .I(n966), .Z(n965) );
  BUFFD0 U990 ( .I(n967), .Z(n966) );
  BUFFD0 U991 ( .I(n968), .Z(n967) );
  BUFFD0 U992 ( .I(n969), .Z(n968) );
  BUFFD0 U993 ( .I(n970), .Z(n969) );
  BUFFD0 U994 ( .I(n971), .Z(n970) );
  BUFFD0 U995 ( .I(n972), .Z(n971) );
  BUFFD0 U996 ( .I(n973), .Z(n972) );
  BUFFD0 U997 ( .I(n974), .Z(n973) );
  BUFFD0 U998 ( .I(n975), .Z(n974) );
  BUFFD0 U999 ( .I(n976), .Z(n975) );
  BUFFD0 U1000 ( .I(n977), .Z(n976) );
  BUFFD0 U1001 ( .I(n978), .Z(n977) );
  BUFFD0 U1002 ( .I(n979), .Z(n978) );
  BUFFD0 U1003 ( .I(n980), .Z(n979) );
  BUFFD0 U1004 ( .I(n981), .Z(n980) );
  BUFFD0 U1005 ( .I(n982), .Z(n981) );
  BUFFD0 U1006 ( .I(n983), .Z(n982) );
  BUFFD0 U1007 ( .I(n984), .Z(n983) );
  BUFFD0 U1008 ( .I(n985), .Z(n984) );
  BUFFD0 U1009 ( .I(n986), .Z(n985) );
  BUFFD0 U1010 ( .I(n987), .Z(n986) );
  BUFFD0 U1011 ( .I(n988), .Z(n987) );
  BUFFD0 U1012 ( .I(n989), .Z(n988) );
  BUFFD0 U1013 ( .I(n990), .Z(n989) );
  BUFFD0 U1014 ( .I(n927), .Z(n990) );
  BUFFD0 U1015 ( .I(n994), .Z(n991) );
  BUFFD0 U1016 ( .I(N57), .Z(n992) );
  BUFFD0 U1017 ( .I(n992), .Z(n993) );
  BUFFD0 U1018 ( .I(n995), .Z(n994) );
  BUFFD0 U1019 ( .I(n996), .Z(n995) );
  BUFFD0 U1020 ( .I(n997), .Z(n996) );
  BUFFD0 U1021 ( .I(n998), .Z(n997) );
  BUFFD0 U1022 ( .I(n999), .Z(n998) );
  BUFFD0 U1023 ( .I(n1000), .Z(n999) );
  BUFFD0 U1024 ( .I(n1001), .Z(n1000) );
  BUFFD0 U1025 ( .I(n1002), .Z(n1001) );
  BUFFD0 U1026 ( .I(n1003), .Z(n1002) );
  BUFFD0 U1027 ( .I(n1004), .Z(n1003) );
  BUFFD0 U1028 ( .I(n1005), .Z(n1004) );
  BUFFD0 U1029 ( .I(n1006), .Z(n1005) );
  BUFFD0 U1030 ( .I(n1007), .Z(n1006) );
  BUFFD0 U1031 ( .I(n1008), .Z(n1007) );
  BUFFD0 U1032 ( .I(n1009), .Z(n1008) );
  BUFFD0 U1033 ( .I(n1010), .Z(n1009) );
  BUFFD0 U1034 ( .I(n1011), .Z(n1010) );
  BUFFD0 U1035 ( .I(n1012), .Z(n1011) );
  BUFFD0 U1036 ( .I(n1013), .Z(n1012) );
  BUFFD0 U1037 ( .I(n1014), .Z(n1013) );
  BUFFD0 U1038 ( .I(n1015), .Z(n1014) );
  BUFFD0 U1039 ( .I(n1016), .Z(n1015) );
  BUFFD0 U1040 ( .I(n1017), .Z(n1016) );
  BUFFD0 U1041 ( .I(n1018), .Z(n1017) );
  BUFFD0 U1042 ( .I(n1019), .Z(n1018) );
  BUFFD0 U1043 ( .I(n1020), .Z(n1019) );
  BUFFD0 U1044 ( .I(n1021), .Z(n1020) );
  BUFFD0 U1045 ( .I(n1022), .Z(n1021) );
  BUFFD0 U1046 ( .I(n1023), .Z(n1022) );
  BUFFD0 U1047 ( .I(n1024), .Z(n1023) );
  BUFFD0 U1048 ( .I(n1025), .Z(n1024) );
  BUFFD0 U1049 ( .I(n1026), .Z(n1025) );
  BUFFD0 U1050 ( .I(n1027), .Z(n1026) );
  BUFFD0 U1051 ( .I(n1028), .Z(n1027) );
  BUFFD0 U1052 ( .I(n1029), .Z(n1028) );
  BUFFD0 U1053 ( .I(n1030), .Z(n1029) );
  BUFFD0 U1054 ( .I(n1031), .Z(n1030) );
  BUFFD0 U1055 ( .I(n1032), .Z(n1031) );
  BUFFD0 U1056 ( .I(n1033), .Z(n1032) );
  BUFFD0 U1057 ( .I(n1034), .Z(n1033) );
  BUFFD0 U1058 ( .I(n1035), .Z(n1034) );
  BUFFD0 U1059 ( .I(n1036), .Z(n1035) );
  BUFFD0 U1060 ( .I(n1037), .Z(n1036) );
  BUFFD0 U1061 ( .I(n1038), .Z(n1037) );
  BUFFD0 U1062 ( .I(n1039), .Z(n1038) );
  BUFFD0 U1063 ( .I(n1040), .Z(n1039) );
  BUFFD0 U1064 ( .I(n1041), .Z(n1040) );
  BUFFD0 U1065 ( .I(n1042), .Z(n1041) );
  BUFFD0 U1066 ( .I(n1043), .Z(n1042) );
  BUFFD0 U1067 ( .I(n1044), .Z(n1043) );
  BUFFD0 U1068 ( .I(n1045), .Z(n1044) );
  BUFFD0 U1069 ( .I(n1046), .Z(n1045) );
  BUFFD0 U1070 ( .I(n1047), .Z(n1046) );
  BUFFD0 U1071 ( .I(n1048), .Z(n1047) );
  BUFFD0 U1072 ( .I(n1049), .Z(n1048) );
  BUFFD0 U1073 ( .I(n1050), .Z(n1049) );
  BUFFD0 U1074 ( .I(n1051), .Z(n1050) );
  BUFFD0 U1075 ( .I(n1052), .Z(n1051) );
  BUFFD0 U1076 ( .I(n1053), .Z(n1052) );
  BUFFD0 U1077 ( .I(n1054), .Z(n1053) );
  BUFFD0 U1078 ( .I(n1055), .Z(n1054) );
  BUFFD0 U1079 ( .I(n1056), .Z(n1055) );
  BUFFD0 U1080 ( .I(n993), .Z(n1056) );
  BUFFD0 U1081 ( .I(n1061), .Z(n1057) );
  BUFFD0 U1082 ( .I(n2612), .Z(n1058) );
  BUFFD0 U1083 ( .I(n1058), .Z(n1059) );
  BUFFD0 U1084 ( .I(n1059), .Z(n1060) );
  BUFFD0 U1085 ( .I(n1062), .Z(n1061) );
  BUFFD0 U1086 ( .I(n1063), .Z(n1062) );
  BUFFD0 U1087 ( .I(n1064), .Z(n1063) );
  BUFFD0 U1088 ( .I(n1065), .Z(n1064) );
  BUFFD0 U1089 ( .I(n1066), .Z(n1065) );
  BUFFD0 U1090 ( .I(n1067), .Z(n1066) );
  BUFFD0 U1091 ( .I(n1068), .Z(n1067) );
  BUFFD0 U1092 ( .I(n1069), .Z(n1068) );
  BUFFD0 U1093 ( .I(n1070), .Z(n1069) );
  BUFFD0 U1094 ( .I(n1071), .Z(n1070) );
  BUFFD0 U1095 ( .I(n1072), .Z(n1071) );
  BUFFD0 U1096 ( .I(n1073), .Z(n1072) );
  BUFFD0 U1097 ( .I(n1074), .Z(n1073) );
  BUFFD0 U1098 ( .I(n1075), .Z(n1074) );
  BUFFD0 U1099 ( .I(n1076), .Z(n1075) );
  BUFFD0 U1100 ( .I(n1077), .Z(n1076) );
  BUFFD0 U1101 ( .I(n1078), .Z(n1077) );
  BUFFD0 U1102 ( .I(n1079), .Z(n1078) );
  BUFFD0 U1103 ( .I(n1080), .Z(n1079) );
  BUFFD0 U1104 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1105 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1106 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1107 ( .I(n1084), .Z(n1083) );
  BUFFD0 U1108 ( .I(n1085), .Z(n1084) );
  BUFFD0 U1109 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1110 ( .I(n1087), .Z(n1086) );
  BUFFD0 U1111 ( .I(n1088), .Z(n1087) );
  BUFFD0 U1112 ( .I(n1089), .Z(n1088) );
  BUFFD0 U1113 ( .I(n1090), .Z(n1089) );
  BUFFD0 U1114 ( .I(n1091), .Z(n1090) );
  BUFFD0 U1115 ( .I(n1092), .Z(n1091) );
  BUFFD0 U1116 ( .I(n1093), .Z(n1092) );
  BUFFD0 U1117 ( .I(n1094), .Z(n1093) );
  BUFFD0 U1118 ( .I(n1095), .Z(n1094) );
  BUFFD0 U1119 ( .I(n1096), .Z(n1095) );
  BUFFD0 U1120 ( .I(n1097), .Z(n1096) );
  BUFFD0 U1121 ( .I(n1098), .Z(n1097) );
  BUFFD0 U1122 ( .I(n1099), .Z(n1098) );
  BUFFD0 U1123 ( .I(n1100), .Z(n1099) );
  BUFFD0 U1124 ( .I(n1101), .Z(n1100) );
  BUFFD0 U1125 ( .I(n1102), .Z(n1101) );
  BUFFD0 U1126 ( .I(n1103), .Z(n1102) );
  BUFFD0 U1127 ( .I(n1104), .Z(n1103) );
  BUFFD0 U1128 ( .I(n1105), .Z(n1104) );
  BUFFD0 U1129 ( .I(n1106), .Z(n1105) );
  BUFFD0 U1130 ( .I(n1107), .Z(n1106) );
  BUFFD0 U1131 ( .I(n1108), .Z(n1107) );
  BUFFD0 U1132 ( .I(n1109), .Z(n1108) );
  BUFFD0 U1133 ( .I(n1110), .Z(n1109) );
  BUFFD0 U1134 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1135 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1136 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1137 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1138 ( .I(n1115), .Z(n1114) );
  BUFFD0 U1139 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1140 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1141 ( .I(n1118), .Z(n1117) );
  BUFFD0 U1142 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1143 ( .I(n1060), .Z(n1119) );
  BUFFD0 U1144 ( .I(N58), .Z(n1120) );
  BUFFD0 U1145 ( .I(n1120), .Z(n1121) );
  BUFFD0 U1146 ( .I(n1121), .Z(n1122) );
  BUFFD0 U1147 ( .I(n1127), .Z(n1123) );
  BUFFD0 U1148 ( .I(N59), .Z(n1124) );
  BUFFD0 U1149 ( .I(n1124), .Z(n1125) );
  BUFFD0 U1150 ( .I(n1125), .Z(n1126) );
  BUFFD0 U1151 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1152 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1153 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1154 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1155 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1156 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1157 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1158 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1159 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1160 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1161 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1162 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1163 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1164 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1165 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1166 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1167 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1168 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1169 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1170 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1171 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1172 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1173 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1174 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1175 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1176 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1177 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1178 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1179 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1180 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1181 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1182 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1183 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1184 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1185 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1186 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1187 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1188 ( .I(n1165), .Z(n1164) );
  BUFFD0 U1189 ( .I(n1166), .Z(n1165) );
  BUFFD0 U1190 ( .I(n1167), .Z(n1166) );
  BUFFD0 U1191 ( .I(n1168), .Z(n1167) );
  BUFFD0 U1192 ( .I(n1169), .Z(n1168) );
  BUFFD0 U1193 ( .I(n1170), .Z(n1169) );
  BUFFD0 U1194 ( .I(n1171), .Z(n1170) );
  BUFFD0 U1195 ( .I(n1172), .Z(n1171) );
  BUFFD0 U1196 ( .I(n1173), .Z(n1172) );
  BUFFD0 U1197 ( .I(n1174), .Z(n1173) );
  BUFFD0 U1198 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1199 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1200 ( .I(n1177), .Z(n1176) );
  BUFFD0 U1201 ( .I(n1178), .Z(n1177) );
  BUFFD0 U1202 ( .I(n1179), .Z(n1178) );
  BUFFD0 U1203 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1204 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1205 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1206 ( .I(n1183), .Z(n1182) );
  BUFFD0 U1207 ( .I(n1184), .Z(n1183) );
  BUFFD0 U1208 ( .I(n2594), .Z(n1184) );
  BUFFD0 U1209 ( .I(n1126), .Z(n1185) );
  BUFFD0 U1210 ( .I(n1185), .Z(n1186) );
  BUFFD0 U1211 ( .I(n1186), .Z(n1187) );
  BUFFD0 U1212 ( .I(n1192), .Z(n1188) );
  BUFFD0 U1213 ( .I(N60), .Z(n1189) );
  BUFFD0 U1214 ( .I(n1189), .Z(n1190) );
  BUFFD0 U1215 ( .I(n1190), .Z(n1191) );
  BUFFD0 U1216 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1217 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1218 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1219 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1220 ( .I(n1197), .Z(n1196) );
  BUFFD0 U1221 ( .I(n1198), .Z(n1197) );
  BUFFD0 U1222 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1223 ( .I(n1200), .Z(n1199) );
  BUFFD0 U1224 ( .I(n1201), .Z(n1200) );
  BUFFD0 U1225 ( .I(n1202), .Z(n1201) );
  BUFFD0 U1226 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1227 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1228 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1229 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1230 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1231 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1232 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1233 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1234 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1235 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1236 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1237 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1238 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1239 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1240 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1241 ( .I(n1218), .Z(n1217) );
  BUFFD0 U1242 ( .I(n1219), .Z(n1218) );
  BUFFD0 U1243 ( .I(n1220), .Z(n1219) );
  BUFFD0 U1244 ( .I(n1221), .Z(n1220) );
  BUFFD0 U1245 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1246 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1247 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1248 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1249 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1250 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1251 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1252 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1253 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1254 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1255 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1256 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1257 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1258 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1259 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1260 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1261 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1262 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1263 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1264 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1265 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1266 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1267 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1268 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1269 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1270 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1271 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1272 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1273 ( .I(n2601), .Z(n1249) );
  BUFFD0 U1274 ( .I(n1191), .Z(n1250) );
  BUFFD0 U1275 ( .I(n1250), .Z(n1251) );
  BUFFD0 U1276 ( .I(n1251), .Z(n1252) );
  BUFFD0 U1277 ( .I(n1252), .Z(n1253) );
  BUFFD0 U1278 ( .I(n1258), .Z(n1254) );
  BUFFD0 U1279 ( .I(n2593), .Z(n1255) );
  BUFFD0 U1280 ( .I(n1255), .Z(n1256) );
  BUFFD0 U1281 ( .I(n1256), .Z(n1257) );
  BUFFD0 U1282 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1283 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1284 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1285 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1286 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1287 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1288 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1289 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1290 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1291 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1292 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1293 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1294 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1295 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1296 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1297 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1298 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1299 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1300 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1301 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1302 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1303 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1304 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1305 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1306 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1307 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1308 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1309 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1310 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1311 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1312 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1313 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1314 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1315 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1316 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1317 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1318 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1319 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1320 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1321 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1322 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1323 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1324 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1325 ( .I(n1302), .Z(n1301) );
  BUFFD0 U1326 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1327 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1328 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1329 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1330 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1331 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1332 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1333 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1334 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1335 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1336 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1337 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1338 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1339 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1340 ( .I(n1257), .Z(n1316) );
  BUFFD0 U1341 ( .I(N61), .Z(n1317) );
  BUFFD0 U1342 ( .I(n1317), .Z(n1318) );
  BUFFD0 U1343 ( .I(n1318), .Z(n1319) );
  BUFFD0 U1344 ( .I(n1324), .Z(n1320) );
  BUFFD0 U1345 ( .I(n2600), .Z(n1321) );
  BUFFD0 U1346 ( .I(n1321), .Z(n1322) );
  BUFFD0 U1347 ( .I(n1322), .Z(n1323) );
  BUFFD0 U1348 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1349 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1350 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1351 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1352 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1353 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1354 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1355 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1356 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1357 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1358 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1359 ( .I(n1336), .Z(n1335) );
  BUFFD0 U1360 ( .I(n1337), .Z(n1336) );
  BUFFD0 U1361 ( .I(n1338), .Z(n1337) );
  BUFFD0 U1362 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1363 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1364 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1365 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1366 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1367 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1368 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1369 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1370 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1371 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1372 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1373 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1374 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1375 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1376 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1377 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1378 ( .I(n1355), .Z(n1354) );
  BUFFD0 U1379 ( .I(n1356), .Z(n1355) );
  BUFFD0 U1380 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1381 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1382 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1383 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1384 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1385 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1386 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1387 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1388 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1389 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1390 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1391 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1392 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1393 ( .I(n1370), .Z(n1369) );
  BUFFD0 U1394 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1395 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1396 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1397 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1398 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1399 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1400 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1401 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1402 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1403 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1404 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1405 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1406 ( .I(n1323), .Z(n1382) );
  BUFFD0 U1407 ( .I(N62), .Z(n1383) );
  BUFFD0 U1408 ( .I(n1383), .Z(n1384) );
  BUFFD0 U1409 ( .I(n1384), .Z(n1385) );
  BUFFD0 U1410 ( .I(n1390), .Z(n1386) );
  BUFFD0 U1411 ( .I(N63), .Z(n1387) );
  BUFFD0 U1412 ( .I(n1387), .Z(n1388) );
  BUFFD0 U1413 ( .I(n1388), .Z(n1389) );
  BUFFD0 U1414 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1415 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1416 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1417 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1418 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1419 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1420 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1421 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1422 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1423 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1424 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1425 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1426 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1427 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1428 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1429 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1430 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1431 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1432 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1433 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1434 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1435 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1436 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1437 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1438 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1439 ( .I(n1416), .Z(n1415) );
  BUFFD0 U1440 ( .I(n1417), .Z(n1416) );
  BUFFD0 U1441 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1442 ( .I(n1419), .Z(n1418) );
  BUFFD0 U1443 ( .I(n1420), .Z(n1419) );
  BUFFD0 U1444 ( .I(n1421), .Z(n1420) );
  BUFFD0 U1445 ( .I(n1422), .Z(n1421) );
  BUFFD0 U1446 ( .I(n1423), .Z(n1422) );
  BUFFD0 U1447 ( .I(n1424), .Z(n1423) );
  BUFFD0 U1448 ( .I(n1425), .Z(n1424) );
  BUFFD0 U1449 ( .I(n1426), .Z(n1425) );
  BUFFD0 U1450 ( .I(n1427), .Z(n1426) );
  BUFFD0 U1451 ( .I(n1428), .Z(n1427) );
  BUFFD0 U1452 ( .I(n1429), .Z(n1428) );
  BUFFD0 U1453 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1454 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1455 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1456 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1457 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1458 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1459 ( .I(n1436), .Z(n1435) );
  BUFFD0 U1460 ( .I(n1437), .Z(n1436) );
  BUFFD0 U1461 ( .I(n1438), .Z(n1437) );
  BUFFD0 U1462 ( .I(n1439), .Z(n1438) );
  BUFFD0 U1463 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1464 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1465 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1466 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1467 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1468 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1469 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1470 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1471 ( .I(n2604), .Z(n1447) );
  BUFFD0 U1472 ( .I(n1389), .Z(n1448) );
  BUFFD0 U1473 ( .I(n1448), .Z(n1449) );
  BUFFD0 U1474 ( .I(n1449), .Z(n1450) );
  BUFFD0 U1475 ( .I(n1450), .Z(n1451) );
  BUFFD0 U1476 ( .I(n1456), .Z(n1452) );
  BUFFD0 U1477 ( .I(n2602), .Z(n1453) );
  BUFFD0 U1478 ( .I(n1453), .Z(n1454) );
  BUFFD0 U1479 ( .I(n1454), .Z(n1455) );
  BUFFD0 U1480 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1481 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1482 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1483 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1484 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1485 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1486 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1487 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1488 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1489 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1490 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1491 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1492 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1493 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1494 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1495 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1496 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1497 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1498 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1499 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1500 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1501 ( .I(n1478), .Z(n1477) );
  BUFFD0 U1502 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1503 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1504 ( .I(n1481), .Z(n1480) );
  BUFFD0 U1505 ( .I(n1482), .Z(n1481) );
  BUFFD0 U1506 ( .I(n1483), .Z(n1482) );
  BUFFD0 U1507 ( .I(n1484), .Z(n1483) );
  BUFFD0 U1508 ( .I(n1485), .Z(n1484) );
  BUFFD0 U1509 ( .I(n1486), .Z(n1485) );
  BUFFD0 U1510 ( .I(n1487), .Z(n1486) );
  BUFFD0 U1511 ( .I(n1488), .Z(n1487) );
  BUFFD0 U1512 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1513 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1514 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1515 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1516 ( .I(n1493), .Z(n1492) );
  BUFFD0 U1517 ( .I(n1494), .Z(n1493) );
  BUFFD0 U1518 ( .I(n1495), .Z(n1494) );
  BUFFD0 U1519 ( .I(n1496), .Z(n1495) );
  BUFFD0 U1520 ( .I(n1497), .Z(n1496) );
  BUFFD0 U1521 ( .I(n1498), .Z(n1497) );
  BUFFD0 U1522 ( .I(n1499), .Z(n1498) );
  BUFFD0 U1523 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1524 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1525 ( .I(n1502), .Z(n1501) );
  BUFFD0 U1526 ( .I(n1503), .Z(n1502) );
  BUFFD0 U1527 ( .I(n1504), .Z(n1503) );
  BUFFD0 U1528 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1529 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1530 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1531 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1532 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1533 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1534 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1535 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1536 ( .I(n1513), .Z(n1512) );
  BUFFD0 U1537 ( .I(n1514), .Z(n1513) );
  BUFFD0 U1538 ( .I(n1455), .Z(n1514) );
  BUFFD0 U1539 ( .I(n1519), .Z(n1515) );
  BUFFD0 U1540 ( .I(n2624), .Z(n1516) );
  BUFFD0 U1541 ( .I(n1516), .Z(n1517) );
  BUFFD0 U1542 ( .I(n1517), .Z(n1518) );
  BUFFD0 U1543 ( .I(n1520), .Z(n1519) );
  BUFFD0 U1544 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1545 ( .I(n1522), .Z(n1521) );
  BUFFD0 U1546 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1547 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1548 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1549 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1550 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1551 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1552 ( .I(n1529), .Z(n1528) );
  BUFFD0 U1553 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1554 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1555 ( .I(n1532), .Z(n1531) );
  BUFFD0 U1556 ( .I(n1533), .Z(n1532) );
  BUFFD0 U1557 ( .I(n1534), .Z(n1533) );
  BUFFD0 U1558 ( .I(n1535), .Z(n1534) );
  BUFFD0 U1559 ( .I(n1536), .Z(n1535) );
  BUFFD0 U1560 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1561 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1562 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1563 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1564 ( .I(n1541), .Z(n1540) );
  BUFFD0 U1565 ( .I(n1542), .Z(n1541) );
  BUFFD0 U1566 ( .I(n1543), .Z(n1542) );
  BUFFD0 U1567 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1568 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1569 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1570 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1571 ( .I(n1548), .Z(n1547) );
  BUFFD0 U1572 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1573 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1574 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1575 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1576 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1577 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1578 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1579 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1580 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1581 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1582 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1583 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1584 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1585 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1586 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1587 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1588 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1589 ( .I(n1566), .Z(n1565) );
  BUFFD0 U1590 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1591 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1592 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1593 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1594 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1595 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1596 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1597 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1598 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1599 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1600 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1601 ( .I(n1518), .Z(n1577) );
  BUFFD0 U1602 ( .I(n1582), .Z(n1578) );
  BUFFD0 U1603 ( .I(N66), .Z(n1579) );
  BUFFD0 U1604 ( .I(n1579), .Z(n1580) );
  BUFFD0 U1605 ( .I(n1580), .Z(n1581) );
  BUFFD0 U1606 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1607 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1608 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1609 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1610 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1611 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1612 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1613 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1614 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1615 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1616 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1617 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1618 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1619 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1620 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1621 ( .I(n1598), .Z(n1597) );
  BUFFD0 U1622 ( .I(n1599), .Z(n1598) );
  BUFFD0 U1623 ( .I(n1600), .Z(n1599) );
  BUFFD0 U1624 ( .I(n1601), .Z(n1600) );
  BUFFD0 U1625 ( .I(n1602), .Z(n1601) );
  BUFFD0 U1626 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1627 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1628 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1629 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1630 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1631 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1632 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1633 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1634 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1635 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1636 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1637 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1638 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1639 ( .I(n1616), .Z(n1615) );
  BUFFD0 U1640 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1641 ( .I(n1618), .Z(n1617) );
  BUFFD0 U1642 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1643 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1644 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1645 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1646 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1647 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1648 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1649 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1650 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1651 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1652 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1653 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1654 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1655 ( .I(n1632), .Z(n1631) );
  BUFFD0 U1656 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1657 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1658 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1659 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1660 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1661 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1662 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1663 ( .I(n2628), .Z(n1639) );
  BUFFD0 U1664 ( .I(n1581), .Z(n1640) );
  BUFFD0 U1665 ( .I(n1645), .Z(n1641) );
  BUFFD0 U1666 ( .I(N67), .Z(n1642) );
  BUFFD0 U1667 ( .I(n1642), .Z(n1643) );
  BUFFD0 U1668 ( .I(n1643), .Z(n1644) );
  BUFFD0 U1669 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1670 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1671 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1672 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1673 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1674 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1675 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1676 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1677 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1678 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1679 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1680 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1681 ( .I(n1658), .Z(n1657) );
  BUFFD0 U1682 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1683 ( .I(n1660), .Z(n1659) );
  BUFFD0 U1684 ( .I(n1661), .Z(n1660) );
  BUFFD0 U1685 ( .I(n1662), .Z(n1661) );
  BUFFD0 U1686 ( .I(n1663), .Z(n1662) );
  BUFFD0 U1687 ( .I(n1664), .Z(n1663) );
  BUFFD0 U1688 ( .I(n1665), .Z(n1664) );
  BUFFD0 U1689 ( .I(n1666), .Z(n1665) );
  BUFFD0 U1690 ( .I(n1667), .Z(n1666) );
  BUFFD0 U1691 ( .I(n1668), .Z(n1667) );
  BUFFD0 U1692 ( .I(n1669), .Z(n1668) );
  BUFFD0 U1693 ( .I(n1670), .Z(n1669) );
  BUFFD0 U1694 ( .I(n1671), .Z(n1670) );
  BUFFD0 U1695 ( .I(n1672), .Z(n1671) );
  BUFFD0 U1696 ( .I(n1673), .Z(n1672) );
  BUFFD0 U1697 ( .I(n1674), .Z(n1673) );
  BUFFD0 U1698 ( .I(n1675), .Z(n1674) );
  BUFFD0 U1699 ( .I(n1676), .Z(n1675) );
  BUFFD0 U1700 ( .I(n1677), .Z(n1676) );
  BUFFD0 U1701 ( .I(n1678), .Z(n1677) );
  BUFFD0 U1702 ( .I(n1679), .Z(n1678) );
  BUFFD0 U1703 ( .I(n1680), .Z(n1679) );
  BUFFD0 U1704 ( .I(n1681), .Z(n1680) );
  BUFFD0 U1705 ( .I(n1682), .Z(n1681) );
  BUFFD0 U1706 ( .I(n1683), .Z(n1682) );
  BUFFD0 U1707 ( .I(n1684), .Z(n1683) );
  BUFFD0 U1708 ( .I(n1685), .Z(n1684) );
  BUFFD0 U1709 ( .I(n1686), .Z(n1685) );
  BUFFD0 U1710 ( .I(n1687), .Z(n1686) );
  BUFFD0 U1711 ( .I(n1688), .Z(n1687) );
  BUFFD0 U1712 ( .I(n1689), .Z(n1688) );
  BUFFD0 U1713 ( .I(n1690), .Z(n1689) );
  BUFFD0 U1714 ( .I(n1691), .Z(n1690) );
  BUFFD0 U1715 ( .I(n1692), .Z(n1691) );
  BUFFD0 U1716 ( .I(n1693), .Z(n1692) );
  BUFFD0 U1717 ( .I(n1694), .Z(n1693) );
  BUFFD0 U1718 ( .I(n1695), .Z(n1694) );
  BUFFD0 U1719 ( .I(n1696), .Z(n1695) );
  BUFFD0 U1720 ( .I(n1697), .Z(n1696) );
  BUFFD0 U1721 ( .I(n1698), .Z(n1697) );
  BUFFD0 U1722 ( .I(n1699), .Z(n1698) );
  BUFFD0 U1723 ( .I(n1700), .Z(n1699) );
  BUFFD0 U1724 ( .I(n1701), .Z(n1700) );
  BUFFD0 U1725 ( .I(n1702), .Z(n1701) );
  BUFFD0 U1726 ( .I(n2639), .Z(n1702) );
  BUFFD0 U1727 ( .I(n1707), .Z(n1703) );
  BUFFD0 U1728 ( .I(n2633), .Z(n1704) );
  BUFFD0 U1729 ( .I(n1704), .Z(n1705) );
  BUFFD0 U1730 ( .I(n1705), .Z(n1706) );
  BUFFD0 U1731 ( .I(n1708), .Z(n1707) );
  BUFFD0 U1732 ( .I(n1709), .Z(n1708) );
  BUFFD0 U1733 ( .I(n1710), .Z(n1709) );
  BUFFD0 U1734 ( .I(n1711), .Z(n1710) );
  BUFFD0 U1735 ( .I(n1712), .Z(n1711) );
  BUFFD0 U1736 ( .I(n1713), .Z(n1712) );
  BUFFD0 U1737 ( .I(n1714), .Z(n1713) );
  BUFFD0 U1738 ( .I(n1715), .Z(n1714) );
  BUFFD0 U1739 ( .I(n1716), .Z(n1715) );
  BUFFD0 U1740 ( .I(n1717), .Z(n1716) );
  BUFFD0 U1741 ( .I(n1718), .Z(n1717) );
  BUFFD0 U1742 ( .I(n1719), .Z(n1718) );
  BUFFD0 U1743 ( .I(n1720), .Z(n1719) );
  BUFFD0 U1744 ( .I(n1721), .Z(n1720) );
  BUFFD0 U1745 ( .I(n1722), .Z(n1721) );
  BUFFD0 U1746 ( .I(n1723), .Z(n1722) );
  BUFFD0 U1747 ( .I(n1724), .Z(n1723) );
  BUFFD0 U1748 ( .I(n1725), .Z(n1724) );
  BUFFD0 U1749 ( .I(n1726), .Z(n1725) );
  BUFFD0 U1750 ( .I(n1727), .Z(n1726) );
  BUFFD0 U1751 ( .I(n1728), .Z(n1727) );
  BUFFD0 U1752 ( .I(n1729), .Z(n1728) );
  BUFFD0 U1753 ( .I(n1730), .Z(n1729) );
  BUFFD0 U1754 ( .I(n1731), .Z(n1730) );
  BUFFD0 U1755 ( .I(n1732), .Z(n1731) );
  BUFFD0 U1756 ( .I(n1733), .Z(n1732) );
  BUFFD0 U1757 ( .I(n1734), .Z(n1733) );
  BUFFD0 U1758 ( .I(n1735), .Z(n1734) );
  BUFFD0 U1759 ( .I(n1736), .Z(n1735) );
  BUFFD0 U1760 ( .I(n1737), .Z(n1736) );
  BUFFD0 U1761 ( .I(n1738), .Z(n1737) );
  BUFFD0 U1762 ( .I(n1739), .Z(n1738) );
  BUFFD0 U1763 ( .I(n1740), .Z(n1739) );
  BUFFD0 U1764 ( .I(n1741), .Z(n1740) );
  BUFFD0 U1765 ( .I(n1742), .Z(n1741) );
  BUFFD0 U1766 ( .I(n1743), .Z(n1742) );
  BUFFD0 U1767 ( .I(n1744), .Z(n1743) );
  BUFFD0 U1768 ( .I(n1745), .Z(n1744) );
  BUFFD0 U1769 ( .I(n1746), .Z(n1745) );
  BUFFD0 U1770 ( .I(n1747), .Z(n1746) );
  BUFFD0 U1771 ( .I(n1748), .Z(n1747) );
  BUFFD0 U1772 ( .I(n1749), .Z(n1748) );
  BUFFD0 U1773 ( .I(n1750), .Z(n1749) );
  BUFFD0 U1774 ( .I(n1751), .Z(n1750) );
  BUFFD0 U1775 ( .I(n1752), .Z(n1751) );
  BUFFD0 U1776 ( .I(n1753), .Z(n1752) );
  BUFFD0 U1777 ( .I(n1754), .Z(n1753) );
  BUFFD0 U1778 ( .I(n1755), .Z(n1754) );
  BUFFD0 U1779 ( .I(n1756), .Z(n1755) );
  BUFFD0 U1780 ( .I(n1757), .Z(n1756) );
  BUFFD0 U1781 ( .I(n1758), .Z(n1757) );
  BUFFD0 U1782 ( .I(n1759), .Z(n1758) );
  BUFFD0 U1783 ( .I(n1760), .Z(n1759) );
  BUFFD0 U1784 ( .I(n1761), .Z(n1760) );
  BUFFD0 U1785 ( .I(n1762), .Z(n1761) );
  BUFFD0 U1786 ( .I(n1763), .Z(n1762) );
  BUFFD0 U1787 ( .I(n1764), .Z(n1763) );
  BUFFD0 U1788 ( .I(n1706), .Z(n1764) );
  BUFFD0 U1789 ( .I(n1769), .Z(n1765) );
  BUFFD0 U1790 ( .I(n2629), .Z(n1766) );
  BUFFD0 U1791 ( .I(n1766), .Z(n1767) );
  BUFFD0 U1792 ( .I(n1767), .Z(n1768) );
  BUFFD0 U1793 ( .I(n1770), .Z(n1769) );
  BUFFD0 U1794 ( .I(n1771), .Z(n1770) );
  BUFFD0 U1795 ( .I(n1772), .Z(n1771) );
  BUFFD0 U1796 ( .I(n1773), .Z(n1772) );
  BUFFD0 U1797 ( .I(n1774), .Z(n1773) );
  BUFFD0 U1798 ( .I(n1775), .Z(n1774) );
  BUFFD0 U1799 ( .I(n1776), .Z(n1775) );
  BUFFD0 U1800 ( .I(n1777), .Z(n1776) );
  BUFFD0 U1801 ( .I(n1778), .Z(n1777) );
  BUFFD0 U1802 ( .I(n1779), .Z(n1778) );
  BUFFD0 U1803 ( .I(n1780), .Z(n1779) );
  BUFFD0 U1804 ( .I(n1781), .Z(n1780) );
  BUFFD0 U1805 ( .I(n1782), .Z(n1781) );
  BUFFD0 U1806 ( .I(n1783), .Z(n1782) );
  BUFFD0 U1807 ( .I(n1784), .Z(n1783) );
  BUFFD0 U1808 ( .I(n1785), .Z(n1784) );
  BUFFD0 U1809 ( .I(n1786), .Z(n1785) );
  BUFFD0 U1810 ( .I(n1787), .Z(n1786) );
  BUFFD0 U1811 ( .I(n1788), .Z(n1787) );
  BUFFD0 U1812 ( .I(n1789), .Z(n1788) );
  BUFFD0 U1813 ( .I(n1790), .Z(n1789) );
  BUFFD0 U1814 ( .I(n1791), .Z(n1790) );
  BUFFD0 U1815 ( .I(n1792), .Z(n1791) );
  BUFFD0 U1816 ( .I(n1793), .Z(n1792) );
  BUFFD0 U1817 ( .I(n1794), .Z(n1793) );
  BUFFD0 U1818 ( .I(n1795), .Z(n1794) );
  BUFFD0 U1819 ( .I(n1796), .Z(n1795) );
  BUFFD0 U1820 ( .I(n1797), .Z(n1796) );
  BUFFD0 U1821 ( .I(n1798), .Z(n1797) );
  BUFFD0 U1822 ( .I(n1799), .Z(n1798) );
  BUFFD0 U1823 ( .I(n1800), .Z(n1799) );
  BUFFD0 U1824 ( .I(n1801), .Z(n1800) );
  BUFFD0 U1825 ( .I(n1802), .Z(n1801) );
  BUFFD0 U1826 ( .I(n1803), .Z(n1802) );
  BUFFD0 U1827 ( .I(n1804), .Z(n1803) );
  BUFFD0 U1828 ( .I(n1805), .Z(n1804) );
  BUFFD0 U1829 ( .I(n1806), .Z(n1805) );
  BUFFD0 U1830 ( .I(n1807), .Z(n1806) );
  BUFFD0 U1831 ( .I(n1808), .Z(n1807) );
  BUFFD0 U1832 ( .I(n1809), .Z(n1808) );
  BUFFD0 U1833 ( .I(n1810), .Z(n1809) );
  BUFFD0 U1834 ( .I(n1811), .Z(n1810) );
  BUFFD0 U1835 ( .I(n1812), .Z(n1811) );
  BUFFD0 U1836 ( .I(n1813), .Z(n1812) );
  BUFFD0 U1837 ( .I(n1814), .Z(n1813) );
  BUFFD0 U1838 ( .I(n1815), .Z(n1814) );
  BUFFD0 U1839 ( .I(n1816), .Z(n1815) );
  BUFFD0 U1840 ( .I(n1817), .Z(n1816) );
  BUFFD0 U1841 ( .I(n1818), .Z(n1817) );
  BUFFD0 U1842 ( .I(n1819), .Z(n1818) );
  BUFFD0 U1843 ( .I(n1820), .Z(n1819) );
  BUFFD0 U1844 ( .I(n1821), .Z(n1820) );
  BUFFD0 U1845 ( .I(n1822), .Z(n1821) );
  BUFFD0 U1846 ( .I(n1823), .Z(n1822) );
  BUFFD0 U1847 ( .I(n1824), .Z(n1823) );
  BUFFD0 U1848 ( .I(n1825), .Z(n1824) );
  BUFFD0 U1849 ( .I(n1826), .Z(n1825) );
  BUFFD0 U1850 ( .I(n1827), .Z(n1826) );
  BUFFD0 U1851 ( .I(n1768), .Z(n1827) );
  BUFFD0 U1852 ( .I(n1832), .Z(n1828) );
  BUFFD0 U1853 ( .I(N70), .Z(n1829) );
  BUFFD0 U1854 ( .I(n1829), .Z(n1830) );
  BUFFD0 U1855 ( .I(n1830), .Z(n1831) );
  BUFFD0 U1856 ( .I(n1833), .Z(n1832) );
  BUFFD0 U1857 ( .I(n1834), .Z(n1833) );
  BUFFD0 U1858 ( .I(n1835), .Z(n1834) );
  BUFFD0 U1859 ( .I(n1836), .Z(n1835) );
  BUFFD0 U1860 ( .I(n1837), .Z(n1836) );
  BUFFD0 U1861 ( .I(n1838), .Z(n1837) );
  BUFFD0 U1862 ( .I(n1839), .Z(n1838) );
  BUFFD0 U1863 ( .I(n1840), .Z(n1839) );
  BUFFD0 U1864 ( .I(n1841), .Z(n1840) );
  BUFFD0 U1865 ( .I(n1842), .Z(n1841) );
  BUFFD0 U1866 ( .I(n1843), .Z(n1842) );
  BUFFD0 U1867 ( .I(n1844), .Z(n1843) );
  BUFFD0 U1868 ( .I(n1845), .Z(n1844) );
  BUFFD0 U1869 ( .I(n1846), .Z(n1845) );
  BUFFD0 U1870 ( .I(n1847), .Z(n1846) );
  BUFFD0 U1871 ( .I(n1848), .Z(n1847) );
  BUFFD0 U1872 ( .I(n1849), .Z(n1848) );
  BUFFD0 U1873 ( .I(n1850), .Z(n1849) );
  BUFFD0 U1874 ( .I(n1851), .Z(n1850) );
  BUFFD0 U1875 ( .I(n1852), .Z(n1851) );
  BUFFD0 U1876 ( .I(n1853), .Z(n1852) );
  BUFFD0 U1877 ( .I(n1854), .Z(n1853) );
  BUFFD0 U1878 ( .I(n1855), .Z(n1854) );
  BUFFD0 U1879 ( .I(n1856), .Z(n1855) );
  BUFFD0 U1880 ( .I(n1857), .Z(n1856) );
  BUFFD0 U1881 ( .I(n1858), .Z(n1857) );
  BUFFD0 U1882 ( .I(n1859), .Z(n1858) );
  BUFFD0 U1883 ( .I(n1860), .Z(n1859) );
  BUFFD0 U1884 ( .I(n1861), .Z(n1860) );
  BUFFD0 U1885 ( .I(n1862), .Z(n1861) );
  BUFFD0 U1886 ( .I(n1863), .Z(n1862) );
  BUFFD0 U1887 ( .I(n1864), .Z(n1863) );
  BUFFD0 U1888 ( .I(n1865), .Z(n1864) );
  BUFFD0 U1889 ( .I(n1866), .Z(n1865) );
  BUFFD0 U1890 ( .I(n1867), .Z(n1866) );
  BUFFD0 U1891 ( .I(n1868), .Z(n1867) );
  BUFFD0 U1892 ( .I(n1869), .Z(n1868) );
  BUFFD0 U1893 ( .I(n1870), .Z(n1869) );
  BUFFD0 U1894 ( .I(n1871), .Z(n1870) );
  BUFFD0 U1895 ( .I(n1872), .Z(n1871) );
  BUFFD0 U1896 ( .I(n1873), .Z(n1872) );
  BUFFD0 U1897 ( .I(n1874), .Z(n1873) );
  BUFFD0 U1898 ( .I(n1875), .Z(n1874) );
  BUFFD0 U1899 ( .I(n1876), .Z(n1875) );
  BUFFD0 U1900 ( .I(n1877), .Z(n1876) );
  BUFFD0 U1901 ( .I(n1878), .Z(n1877) );
  BUFFD0 U1902 ( .I(n1879), .Z(n1878) );
  BUFFD0 U1903 ( .I(n1880), .Z(n1879) );
  BUFFD0 U1904 ( .I(n1881), .Z(n1880) );
  BUFFD0 U1905 ( .I(n1882), .Z(n1881) );
  BUFFD0 U1906 ( .I(n1883), .Z(n1882) );
  BUFFD0 U1907 ( .I(n1884), .Z(n1883) );
  BUFFD0 U1908 ( .I(n1885), .Z(n1884) );
  BUFFD0 U1909 ( .I(n1886), .Z(n1885) );
  BUFFD0 U1910 ( .I(n1887), .Z(n1886) );
  BUFFD0 U1911 ( .I(n1888), .Z(n1887) );
  BUFFD0 U1912 ( .I(n1889), .Z(n1888) );
  BUFFD0 U1913 ( .I(n2631), .Z(n1889) );
  BUFFD0 U1914 ( .I(n1831), .Z(n1890) );
  BUFFD0 U1915 ( .I(n1895), .Z(n1891) );
  BUFFD0 U1916 ( .I(N71), .Z(n1892) );
  BUFFD0 U1917 ( .I(n1892), .Z(n1893) );
  BUFFD0 U1918 ( .I(n1893), .Z(n1894) );
  BUFFD0 U1919 ( .I(n1896), .Z(n1895) );
  BUFFD0 U1920 ( .I(n1897), .Z(n1896) );
  BUFFD0 U1921 ( .I(n1898), .Z(n1897) );
  BUFFD0 U1922 ( .I(n1899), .Z(n1898) );
  BUFFD0 U1923 ( .I(n1900), .Z(n1899) );
  BUFFD0 U1924 ( .I(n1901), .Z(n1900) );
  BUFFD0 U1925 ( .I(n1902), .Z(n1901) );
  BUFFD0 U1926 ( .I(n1903), .Z(n1902) );
  BUFFD0 U1927 ( .I(n1904), .Z(n1903) );
  BUFFD0 U1928 ( .I(n1905), .Z(n1904) );
  BUFFD0 U1929 ( .I(n1906), .Z(n1905) );
  BUFFD0 U1930 ( .I(n1907), .Z(n1906) );
  BUFFD0 U1931 ( .I(n1908), .Z(n1907) );
  BUFFD0 U1932 ( .I(n1909), .Z(n1908) );
  BUFFD0 U1933 ( .I(n1910), .Z(n1909) );
  BUFFD0 U1934 ( .I(n1911), .Z(n1910) );
  BUFFD0 U1935 ( .I(n1912), .Z(n1911) );
  BUFFD0 U1936 ( .I(n1913), .Z(n1912) );
  BUFFD0 U1937 ( .I(n1914), .Z(n1913) );
  BUFFD0 U1938 ( .I(n1915), .Z(n1914) );
  BUFFD0 U1939 ( .I(n1916), .Z(n1915) );
  BUFFD0 U1940 ( .I(n1917), .Z(n1916) );
  BUFFD0 U1941 ( .I(n1918), .Z(n1917) );
  BUFFD0 U1942 ( .I(n1919), .Z(n1918) );
  BUFFD0 U1943 ( .I(n1920), .Z(n1919) );
  BUFFD0 U1944 ( .I(n1921), .Z(n1920) );
  BUFFD0 U1945 ( .I(n1922), .Z(n1921) );
  BUFFD0 U1946 ( .I(n1923), .Z(n1922) );
  BUFFD0 U1947 ( .I(n1924), .Z(n1923) );
  BUFFD0 U1948 ( .I(n1925), .Z(n1924) );
  BUFFD0 U1949 ( .I(n1926), .Z(n1925) );
  BUFFD0 U1950 ( .I(n1927), .Z(n1926) );
  BUFFD0 U1951 ( .I(n1928), .Z(n1927) );
  BUFFD0 U1952 ( .I(n1929), .Z(n1928) );
  BUFFD0 U1953 ( .I(n1930), .Z(n1929) );
  BUFFD0 U1954 ( .I(n1931), .Z(n1930) );
  BUFFD0 U1955 ( .I(n1932), .Z(n1931) );
  BUFFD0 U1956 ( .I(n1933), .Z(n1932) );
  BUFFD0 U1957 ( .I(n1934), .Z(n1933) );
  BUFFD0 U1958 ( .I(n1935), .Z(n1934) );
  BUFFD0 U1959 ( .I(n1936), .Z(n1935) );
  BUFFD0 U1960 ( .I(n1937), .Z(n1936) );
  BUFFD0 U1961 ( .I(n1938), .Z(n1937) );
  BUFFD0 U1962 ( .I(n1939), .Z(n1938) );
  BUFFD0 U1963 ( .I(n1940), .Z(n1939) );
  BUFFD0 U1964 ( .I(n1941), .Z(n1940) );
  BUFFD0 U1965 ( .I(n1942), .Z(n1941) );
  BUFFD0 U1966 ( .I(n1943), .Z(n1942) );
  BUFFD0 U1967 ( .I(n1944), .Z(n1943) );
  BUFFD0 U1968 ( .I(n1945), .Z(n1944) );
  BUFFD0 U1969 ( .I(n1946), .Z(n1945) );
  BUFFD0 U1970 ( .I(n1947), .Z(n1946) );
  BUFFD0 U1971 ( .I(n1948), .Z(n1947) );
  BUFFD0 U1972 ( .I(n1949), .Z(n1948) );
  BUFFD0 U1973 ( .I(n1950), .Z(n1949) );
  BUFFD0 U1974 ( .I(n1951), .Z(n1950) );
  BUFFD0 U1975 ( .I(n2671), .Z(n1951) );
  BUFFD0 U1976 ( .I(n1956), .Z(n1952) );
  BUFFD0 U1977 ( .I(N72), .Z(n1953) );
  BUFFD0 U1978 ( .I(n1953), .Z(n1954) );
  BUFFD0 U1979 ( .I(n1954), .Z(n1955) );
  BUFFD0 U1980 ( .I(n1957), .Z(n1956) );
  BUFFD0 U1981 ( .I(n1958), .Z(n1957) );
  BUFFD0 U1982 ( .I(n1959), .Z(n1958) );
  BUFFD0 U1983 ( .I(n1960), .Z(n1959) );
  BUFFD0 U1984 ( .I(n1961), .Z(n1960) );
  BUFFD0 U1985 ( .I(n1962), .Z(n1961) );
  BUFFD0 U1986 ( .I(n1963), .Z(n1962) );
  BUFFD0 U1987 ( .I(n1964), .Z(n1963) );
  BUFFD0 U1988 ( .I(n1965), .Z(n1964) );
  BUFFD0 U1989 ( .I(n1966), .Z(n1965) );
  BUFFD0 U1990 ( .I(n1967), .Z(n1966) );
  BUFFD0 U1991 ( .I(n1968), .Z(n1967) );
  BUFFD0 U1992 ( .I(n1969), .Z(n1968) );
  BUFFD0 U1993 ( .I(n1970), .Z(n1969) );
  BUFFD0 U1994 ( .I(n1971), .Z(n1970) );
  BUFFD0 U1995 ( .I(n1972), .Z(n1971) );
  BUFFD0 U1996 ( .I(n1973), .Z(n1972) );
  BUFFD0 U1997 ( .I(n1974), .Z(n1973) );
  BUFFD0 U1998 ( .I(n1975), .Z(n1974) );
  BUFFD0 U1999 ( .I(n1976), .Z(n1975) );
  BUFFD0 U2000 ( .I(n1977), .Z(n1976) );
  BUFFD0 U2001 ( .I(n1978), .Z(n1977) );
  BUFFD0 U2002 ( .I(n1979), .Z(n1978) );
  BUFFD0 U2003 ( .I(n1980), .Z(n1979) );
  BUFFD0 U2004 ( .I(n1981), .Z(n1980) );
  BUFFD0 U2005 ( .I(n1982), .Z(n1981) );
  BUFFD0 U2006 ( .I(n1983), .Z(n1982) );
  BUFFD0 U2007 ( .I(n1984), .Z(n1983) );
  BUFFD0 U2008 ( .I(n1985), .Z(n1984) );
  BUFFD0 U2009 ( .I(n1986), .Z(n1985) );
  BUFFD0 U2010 ( .I(n1987), .Z(n1986) );
  BUFFD0 U2011 ( .I(n1988), .Z(n1987) );
  BUFFD0 U2012 ( .I(n1989), .Z(n1988) );
  BUFFD0 U2013 ( .I(n1990), .Z(n1989) );
  BUFFD0 U2014 ( .I(n1991), .Z(n1990) );
  BUFFD0 U2015 ( .I(n1992), .Z(n1991) );
  BUFFD0 U2016 ( .I(n1993), .Z(n1992) );
  BUFFD0 U2017 ( .I(n1994), .Z(n1993) );
  BUFFD0 U2018 ( .I(n1995), .Z(n1994) );
  BUFFD0 U2019 ( .I(n1996), .Z(n1995) );
  BUFFD0 U2020 ( .I(n1997), .Z(n1996) );
  BUFFD0 U2021 ( .I(n1998), .Z(n1997) );
  BUFFD0 U2022 ( .I(n1999), .Z(n1998) );
  BUFFD0 U2023 ( .I(n2000), .Z(n1999) );
  BUFFD0 U2024 ( .I(n2001), .Z(n2000) );
  BUFFD0 U2025 ( .I(n2002), .Z(n2001) );
  BUFFD0 U2026 ( .I(n2003), .Z(n2002) );
  BUFFD0 U2027 ( .I(n2004), .Z(n2003) );
  BUFFD0 U2028 ( .I(n2005), .Z(n2004) );
  BUFFD0 U2029 ( .I(n2006), .Z(n2005) );
  BUFFD0 U2030 ( .I(n2007), .Z(n2006) );
  BUFFD0 U2031 ( .I(n2008), .Z(n2007) );
  BUFFD0 U2032 ( .I(n2009), .Z(n2008) );
  BUFFD0 U2033 ( .I(n2700), .Z(n2009) );
  BUFFD0 U2034 ( .I(n2014), .Z(n2010) );
  BUFFD0 U2035 ( .I(n2706), .Z(n2011) );
  BUFFD0 U2036 ( .I(n2011), .Z(n2012) );
  BUFFD0 U2037 ( .I(n2012), .Z(n2013) );
  BUFFD0 U2038 ( .I(n2015), .Z(n2014) );
  BUFFD0 U2039 ( .I(n2016), .Z(n2015) );
  BUFFD0 U2040 ( .I(n2017), .Z(n2016) );
  BUFFD0 U2041 ( .I(n2018), .Z(n2017) );
  BUFFD0 U2042 ( .I(n2019), .Z(n2018) );
  BUFFD0 U2043 ( .I(n2020), .Z(n2019) );
  BUFFD0 U2044 ( .I(n2021), .Z(n2020) );
  BUFFD0 U2045 ( .I(n2022), .Z(n2021) );
  BUFFD0 U2046 ( .I(n2023), .Z(n2022) );
  BUFFD0 U2047 ( .I(n2024), .Z(n2023) );
  BUFFD0 U2048 ( .I(n2025), .Z(n2024) );
  BUFFD0 U2049 ( .I(n2026), .Z(n2025) );
  BUFFD0 U2050 ( .I(n2027), .Z(n2026) );
  BUFFD0 U2051 ( .I(n2028), .Z(n2027) );
  BUFFD0 U2052 ( .I(n2029), .Z(n2028) );
  BUFFD0 U2053 ( .I(n2030), .Z(n2029) );
  BUFFD0 U2054 ( .I(n2031), .Z(n2030) );
  BUFFD0 U2055 ( .I(n2032), .Z(n2031) );
  BUFFD0 U2056 ( .I(n2033), .Z(n2032) );
  BUFFD0 U2057 ( .I(n2034), .Z(n2033) );
  BUFFD0 U2058 ( .I(n2035), .Z(n2034) );
  BUFFD0 U2059 ( .I(n2036), .Z(n2035) );
  BUFFD0 U2060 ( .I(n2037), .Z(n2036) );
  BUFFD0 U2061 ( .I(n2038), .Z(n2037) );
  BUFFD0 U2062 ( .I(n2039), .Z(n2038) );
  BUFFD0 U2063 ( .I(n2040), .Z(n2039) );
  BUFFD0 U2064 ( .I(n2041), .Z(n2040) );
  BUFFD0 U2065 ( .I(n2042), .Z(n2041) );
  BUFFD0 U2066 ( .I(n2043), .Z(n2042) );
  BUFFD0 U2067 ( .I(n2044), .Z(n2043) );
  BUFFD0 U2068 ( .I(n2045), .Z(n2044) );
  BUFFD0 U2069 ( .I(n2046), .Z(n2045) );
  BUFFD0 U2070 ( .I(n2047), .Z(n2046) );
  BUFFD0 U2071 ( .I(n2048), .Z(n2047) );
  BUFFD0 U2072 ( .I(n2049), .Z(n2048) );
  BUFFD0 U2073 ( .I(n2050), .Z(n2049) );
  BUFFD0 U2074 ( .I(n2051), .Z(n2050) );
  BUFFD0 U2075 ( .I(n2052), .Z(n2051) );
  BUFFD0 U2076 ( .I(n2053), .Z(n2052) );
  BUFFD0 U2077 ( .I(n2054), .Z(n2053) );
  BUFFD0 U2078 ( .I(n2055), .Z(n2054) );
  BUFFD0 U2079 ( .I(n2056), .Z(n2055) );
  BUFFD0 U2080 ( .I(n2057), .Z(n2056) );
  BUFFD0 U2081 ( .I(n2058), .Z(n2057) );
  BUFFD0 U2082 ( .I(n2059), .Z(n2058) );
  BUFFD0 U2083 ( .I(n2060), .Z(n2059) );
  BUFFD0 U2084 ( .I(n2061), .Z(n2060) );
  BUFFD0 U2085 ( .I(n2062), .Z(n2061) );
  BUFFD0 U2086 ( .I(n2063), .Z(n2062) );
  BUFFD0 U2087 ( .I(n2064), .Z(n2063) );
  BUFFD0 U2088 ( .I(n2065), .Z(n2064) );
  BUFFD0 U2089 ( .I(n2066), .Z(n2065) );
  BUFFD0 U2090 ( .I(n2013), .Z(n2066) );
  BUFFD0 U2091 ( .I(n2071), .Z(n2067) );
  BUFFD0 U2092 ( .I(n2670), .Z(n2068) );
  BUFFD0 U2093 ( .I(n2068), .Z(n2069) );
  BUFFD0 U2094 ( .I(n2069), .Z(n2070) );
  BUFFD0 U2095 ( .I(n2072), .Z(n2071) );
  BUFFD0 U2096 ( .I(n2073), .Z(n2072) );
  BUFFD0 U2097 ( .I(n2074), .Z(n2073) );
  BUFFD0 U2098 ( .I(n2075), .Z(n2074) );
  BUFFD0 U2099 ( .I(n2076), .Z(n2075) );
  BUFFD0 U2100 ( .I(n2077), .Z(n2076) );
  BUFFD0 U2101 ( .I(n2078), .Z(n2077) );
  BUFFD0 U2102 ( .I(n2079), .Z(n2078) );
  BUFFD0 U2103 ( .I(n2080), .Z(n2079) );
  BUFFD0 U2104 ( .I(n2081), .Z(n2080) );
  BUFFD0 U2105 ( .I(n2082), .Z(n2081) );
  BUFFD0 U2106 ( .I(n2083), .Z(n2082) );
  BUFFD0 U2107 ( .I(n2084), .Z(n2083) );
  BUFFD0 U2108 ( .I(n2085), .Z(n2084) );
  BUFFD0 U2109 ( .I(n2086), .Z(n2085) );
  BUFFD0 U2110 ( .I(n2087), .Z(n2086) );
  BUFFD0 U2111 ( .I(n2088), .Z(n2087) );
  BUFFD0 U2112 ( .I(n2089), .Z(n2088) );
  BUFFD0 U2113 ( .I(n2090), .Z(n2089) );
  BUFFD0 U2114 ( .I(n2091), .Z(n2090) );
  BUFFD0 U2115 ( .I(n2092), .Z(n2091) );
  BUFFD0 U2116 ( .I(n2093), .Z(n2092) );
  BUFFD0 U2117 ( .I(n2094), .Z(n2093) );
  BUFFD0 U2118 ( .I(n2095), .Z(n2094) );
  BUFFD0 U2119 ( .I(n2096), .Z(n2095) );
  BUFFD0 U2120 ( .I(n2097), .Z(n2096) );
  BUFFD0 U2121 ( .I(n2098), .Z(n2097) );
  BUFFD0 U2122 ( .I(n2099), .Z(n2098) );
  BUFFD0 U2123 ( .I(n2100), .Z(n2099) );
  BUFFD0 U2124 ( .I(n2101), .Z(n2100) );
  BUFFD0 U2125 ( .I(n2102), .Z(n2101) );
  BUFFD0 U2126 ( .I(n2103), .Z(n2102) );
  BUFFD0 U2127 ( .I(n2104), .Z(n2103) );
  BUFFD0 U2128 ( .I(n2105), .Z(n2104) );
  BUFFD0 U2129 ( .I(n2106), .Z(n2105) );
  BUFFD0 U2130 ( .I(n2107), .Z(n2106) );
  BUFFD0 U2131 ( .I(n2108), .Z(n2107) );
  BUFFD0 U2132 ( .I(n2109), .Z(n2108) );
  BUFFD0 U2133 ( .I(n2110), .Z(n2109) );
  BUFFD0 U2134 ( .I(n2111), .Z(n2110) );
  BUFFD0 U2135 ( .I(n2112), .Z(n2111) );
  BUFFD0 U2136 ( .I(n2113), .Z(n2112) );
  BUFFD0 U2137 ( .I(n2114), .Z(n2113) );
  BUFFD0 U2138 ( .I(n2115), .Z(n2114) );
  BUFFD0 U2139 ( .I(n2116), .Z(n2115) );
  BUFFD0 U2140 ( .I(n2117), .Z(n2116) );
  BUFFD0 U2141 ( .I(n2118), .Z(n2117) );
  BUFFD0 U2142 ( .I(n2119), .Z(n2118) );
  BUFFD0 U2143 ( .I(n2120), .Z(n2119) );
  BUFFD0 U2144 ( .I(n2121), .Z(n2120) );
  BUFFD0 U2145 ( .I(n2122), .Z(n2121) );
  BUFFD0 U2146 ( .I(n2123), .Z(n2122) );
  BUFFD0 U2147 ( .I(n2124), .Z(n2123) );
  BUFFD0 U2148 ( .I(n2125), .Z(n2124) );
  BUFFD0 U2149 ( .I(n2126), .Z(n2125) );
  BUFFD0 U2150 ( .I(n2070), .Z(n2126) );
  BUFFD0 U2151 ( .I(n2131), .Z(n2127) );
  BUFFD0 U2152 ( .I(n2681), .Z(n2128) );
  BUFFD0 U2153 ( .I(n2128), .Z(n2129) );
  BUFFD0 U2154 ( .I(n2129), .Z(n2130) );
  BUFFD0 U2155 ( .I(n2132), .Z(n2131) );
  BUFFD0 U2156 ( .I(n2133), .Z(n2132) );
  BUFFD0 U2157 ( .I(n2134), .Z(n2133) );
  BUFFD0 U2158 ( .I(n2135), .Z(n2134) );
  BUFFD0 U2159 ( .I(n2136), .Z(n2135) );
  BUFFD0 U2160 ( .I(n2137), .Z(n2136) );
  BUFFD0 U2161 ( .I(n2138), .Z(n2137) );
  BUFFD0 U2162 ( .I(n2139), .Z(n2138) );
  BUFFD0 U2163 ( .I(n2140), .Z(n2139) );
  BUFFD0 U2164 ( .I(n2141), .Z(n2140) );
  BUFFD0 U2165 ( .I(n2142), .Z(n2141) );
  BUFFD0 U2166 ( .I(n2143), .Z(n2142) );
  BUFFD0 U2167 ( .I(n2144), .Z(n2143) );
  BUFFD0 U2168 ( .I(n2145), .Z(n2144) );
  BUFFD0 U2169 ( .I(n2146), .Z(n2145) );
  BUFFD0 U2170 ( .I(n2147), .Z(n2146) );
  BUFFD0 U2171 ( .I(n2148), .Z(n2147) );
  BUFFD0 U2172 ( .I(n2149), .Z(n2148) );
  BUFFD0 U2173 ( .I(n2150), .Z(n2149) );
  BUFFD0 U2174 ( .I(n2151), .Z(n2150) );
  BUFFD0 U2175 ( .I(n2152), .Z(n2151) );
  BUFFD0 U2176 ( .I(n2153), .Z(n2152) );
  BUFFD0 U2177 ( .I(n2154), .Z(n2153) );
  BUFFD0 U2178 ( .I(n2155), .Z(n2154) );
  BUFFD0 U2179 ( .I(n2156), .Z(n2155) );
  BUFFD0 U2180 ( .I(n2157), .Z(n2156) );
  BUFFD0 U2181 ( .I(n2158), .Z(n2157) );
  BUFFD0 U2182 ( .I(n2159), .Z(n2158) );
  BUFFD0 U2183 ( .I(n2160), .Z(n2159) );
  BUFFD0 U2184 ( .I(n2161), .Z(n2160) );
  BUFFD0 U2185 ( .I(n2162), .Z(n2161) );
  BUFFD0 U2186 ( .I(n2163), .Z(n2162) );
  BUFFD0 U2187 ( .I(n2164), .Z(n2163) );
  BUFFD0 U2188 ( .I(n2165), .Z(n2164) );
  BUFFD0 U2189 ( .I(n2166), .Z(n2165) );
  BUFFD0 U2190 ( .I(n2167), .Z(n2166) );
  BUFFD0 U2191 ( .I(n2168), .Z(n2167) );
  BUFFD0 U2192 ( .I(n2169), .Z(n2168) );
  BUFFD0 U2193 ( .I(n2170), .Z(n2169) );
  BUFFD0 U2194 ( .I(n2171), .Z(n2170) );
  BUFFD0 U2195 ( .I(n2172), .Z(n2171) );
  BUFFD0 U2196 ( .I(n2173), .Z(n2172) );
  BUFFD0 U2197 ( .I(n2174), .Z(n2173) );
  BUFFD0 U2198 ( .I(n2175), .Z(n2174) );
  BUFFD0 U2199 ( .I(n2176), .Z(n2175) );
  BUFFD0 U2200 ( .I(n2177), .Z(n2176) );
  BUFFD0 U2201 ( .I(n2178), .Z(n2177) );
  BUFFD0 U2202 ( .I(n2179), .Z(n2178) );
  BUFFD0 U2203 ( .I(n2180), .Z(n2179) );
  BUFFD0 U2204 ( .I(n2181), .Z(n2180) );
  BUFFD0 U2205 ( .I(n2182), .Z(n2181) );
  BUFFD0 U2206 ( .I(n2183), .Z(n2182) );
  BUFFD0 U2207 ( .I(n2184), .Z(n2183) );
  BUFFD0 U2208 ( .I(n2185), .Z(n2184) );
  BUFFD0 U2209 ( .I(n2130), .Z(n2185) );
  BUFFD0 U2210 ( .I(n2190), .Z(n2186) );
  BUFFD0 U2211 ( .I(N76), .Z(n2187) );
  BUFFD0 U2212 ( .I(n2187), .Z(n2188) );
  BUFFD0 U2213 ( .I(n2188), .Z(n2189) );
  BUFFD0 U2214 ( .I(n2191), .Z(n2190) );
  BUFFD0 U2215 ( .I(n2192), .Z(n2191) );
  BUFFD0 U2216 ( .I(n2193), .Z(n2192) );
  BUFFD0 U2217 ( .I(n2194), .Z(n2193) );
  BUFFD0 U2218 ( .I(n2195), .Z(n2194) );
  BUFFD0 U2219 ( .I(n2196), .Z(n2195) );
  BUFFD0 U2220 ( .I(n2197), .Z(n2196) );
  BUFFD0 U2221 ( .I(n2198), .Z(n2197) );
  BUFFD0 U2222 ( .I(n2199), .Z(n2198) );
  BUFFD0 U2223 ( .I(n2200), .Z(n2199) );
  BUFFD0 U2224 ( .I(n2201), .Z(n2200) );
  BUFFD0 U2225 ( .I(n2202), .Z(n2201) );
  BUFFD0 U2226 ( .I(n2203), .Z(n2202) );
  BUFFD0 U2227 ( .I(n2204), .Z(n2203) );
  BUFFD0 U2228 ( .I(n2205), .Z(n2204) );
  BUFFD0 U2229 ( .I(n2206), .Z(n2205) );
  BUFFD0 U2230 ( .I(n2207), .Z(n2206) );
  BUFFD0 U2231 ( .I(n2208), .Z(n2207) );
  BUFFD0 U2232 ( .I(n2209), .Z(n2208) );
  BUFFD0 U2233 ( .I(n2210), .Z(n2209) );
  BUFFD0 U2234 ( .I(n2211), .Z(n2210) );
  BUFFD0 U2235 ( .I(n2212), .Z(n2211) );
  BUFFD0 U2236 ( .I(n2213), .Z(n2212) );
  BUFFD0 U2237 ( .I(n2214), .Z(n2213) );
  BUFFD0 U2238 ( .I(n2215), .Z(n2214) );
  BUFFD0 U2239 ( .I(n2216), .Z(n2215) );
  BUFFD0 U2240 ( .I(n2217), .Z(n2216) );
  BUFFD0 U2241 ( .I(n2218), .Z(n2217) );
  BUFFD0 U2242 ( .I(n2219), .Z(n2218) );
  BUFFD0 U2243 ( .I(n2220), .Z(n2219) );
  BUFFD0 U2244 ( .I(n2221), .Z(n2220) );
  BUFFD0 U2245 ( .I(n2222), .Z(n2221) );
  BUFFD0 U2246 ( .I(n2223), .Z(n2222) );
  BUFFD0 U2247 ( .I(n2224), .Z(n2223) );
  BUFFD0 U2248 ( .I(n2225), .Z(n2224) );
  BUFFD0 U2249 ( .I(n2226), .Z(n2225) );
  BUFFD0 U2250 ( .I(n2227), .Z(n2226) );
  BUFFD0 U2251 ( .I(n2228), .Z(n2227) );
  BUFFD0 U2252 ( .I(n2229), .Z(n2228) );
  BUFFD0 U2253 ( .I(n2230), .Z(n2229) );
  BUFFD0 U2254 ( .I(n2231), .Z(n2230) );
  BUFFD0 U2255 ( .I(n2232), .Z(n2231) );
  BUFFD0 U2256 ( .I(n2233), .Z(n2232) );
  BUFFD0 U2257 ( .I(n2234), .Z(n2233) );
  BUFFD0 U2258 ( .I(n2235), .Z(n2234) );
  BUFFD0 U2259 ( .I(n2236), .Z(n2235) );
  BUFFD0 U2260 ( .I(n2237), .Z(n2236) );
  BUFFD0 U2261 ( .I(n2238), .Z(n2237) );
  BUFFD0 U2262 ( .I(n2239), .Z(n2238) );
  BUFFD0 U2263 ( .I(n2240), .Z(n2239) );
  BUFFD0 U2264 ( .I(n2241), .Z(n2240) );
  BUFFD0 U2265 ( .I(n2242), .Z(n2241) );
  BUFFD0 U2266 ( .I(n2243), .Z(n2242) );
  BUFFD0 U2267 ( .I(n2244), .Z(n2243) );
  BUFFD0 U2268 ( .I(n2684), .Z(n2244) );
  BUFFD0 U2269 ( .I(n2249), .Z(n2245) );
  BUFFD0 U2270 ( .I(N77), .Z(n2246) );
  BUFFD0 U2271 ( .I(n2246), .Z(n2247) );
  BUFFD0 U2272 ( .I(n2247), .Z(n2248) );
  BUFFD0 U2273 ( .I(n2250), .Z(n2249) );
  BUFFD0 U2274 ( .I(n2251), .Z(n2250) );
  BUFFD0 U2275 ( .I(n2252), .Z(n2251) );
  BUFFD0 U2276 ( .I(n2253), .Z(n2252) );
  BUFFD0 U2277 ( .I(n2254), .Z(n2253) );
  BUFFD0 U2278 ( .I(n2255), .Z(n2254) );
  BUFFD0 U2279 ( .I(n2256), .Z(n2255) );
  BUFFD0 U2280 ( .I(n2257), .Z(n2256) );
  BUFFD0 U2281 ( .I(n2258), .Z(n2257) );
  BUFFD0 U2282 ( .I(n2259), .Z(n2258) );
  BUFFD0 U2283 ( .I(n2260), .Z(n2259) );
  BUFFD0 U2284 ( .I(n2261), .Z(n2260) );
  BUFFD0 U2285 ( .I(n2262), .Z(n2261) );
  BUFFD0 U2286 ( .I(n2263), .Z(n2262) );
  BUFFD0 U2287 ( .I(n2264), .Z(n2263) );
  BUFFD0 U2288 ( .I(n2265), .Z(n2264) );
  BUFFD0 U2289 ( .I(n2266), .Z(n2265) );
  BUFFD0 U2290 ( .I(n2267), .Z(n2266) );
  BUFFD0 U2291 ( .I(n2268), .Z(n2267) );
  BUFFD0 U2292 ( .I(n2269), .Z(n2268) );
  BUFFD0 U2293 ( .I(n2270), .Z(n2269) );
  BUFFD0 U2294 ( .I(n2271), .Z(n2270) );
  BUFFD0 U2295 ( .I(n2272), .Z(n2271) );
  BUFFD0 U2296 ( .I(n2273), .Z(n2272) );
  BUFFD0 U2297 ( .I(n2274), .Z(n2273) );
  BUFFD0 U2298 ( .I(n2275), .Z(n2274) );
  BUFFD0 U2299 ( .I(n2276), .Z(n2275) );
  BUFFD0 U2300 ( .I(n2277), .Z(n2276) );
  BUFFD0 U2301 ( .I(n2278), .Z(n2277) );
  BUFFD0 U2302 ( .I(n2279), .Z(n2278) );
  BUFFD0 U2303 ( .I(n2280), .Z(n2279) );
  BUFFD0 U2304 ( .I(n2281), .Z(n2280) );
  BUFFD0 U2305 ( .I(n2282), .Z(n2281) );
  BUFFD0 U2306 ( .I(n2283), .Z(n2282) );
  BUFFD0 U2307 ( .I(n2284), .Z(n2283) );
  BUFFD0 U2308 ( .I(n2285), .Z(n2284) );
  BUFFD0 U2309 ( .I(n2286), .Z(n2285) );
  BUFFD0 U2310 ( .I(n2287), .Z(n2286) );
  BUFFD0 U2311 ( .I(n2288), .Z(n2287) );
  BUFFD0 U2312 ( .I(n2289), .Z(n2288) );
  BUFFD0 U2313 ( .I(n2290), .Z(n2289) );
  BUFFD0 U2314 ( .I(n2291), .Z(n2290) );
  BUFFD0 U2315 ( .I(n2292), .Z(n2291) );
  BUFFD0 U2316 ( .I(n2293), .Z(n2292) );
  BUFFD0 U2317 ( .I(n2294), .Z(n2293) );
  BUFFD0 U2318 ( .I(n2295), .Z(n2294) );
  BUFFD0 U2319 ( .I(n2296), .Z(n2295) );
  BUFFD0 U2320 ( .I(n2297), .Z(n2296) );
  BUFFD0 U2321 ( .I(n2298), .Z(n2297) );
  BUFFD0 U2322 ( .I(n2299), .Z(n2298) );
  BUFFD0 U2323 ( .I(n2300), .Z(n2299) );
  BUFFD0 U2324 ( .I(n2301), .Z(n2300) );
  BUFFD0 U2325 ( .I(n2302), .Z(n2301) );
  BUFFD0 U2326 ( .I(n2303), .Z(n2302) );
  BUFFD0 U2327 ( .I(n2677), .Z(n2303) );
  BUFFD0 U2328 ( .I(n2308), .Z(n2304) );
  BUFFD0 U2329 ( .I(N78), .Z(n2305) );
  BUFFD0 U2330 ( .I(n2305), .Z(n2306) );
  BUFFD0 U2331 ( .I(n2306), .Z(n2307) );
  BUFFD0 U2332 ( .I(n2309), .Z(n2308) );
  BUFFD0 U2333 ( .I(n2310), .Z(n2309) );
  BUFFD0 U2334 ( .I(n2311), .Z(n2310) );
  BUFFD0 U2335 ( .I(n2312), .Z(n2311) );
  BUFFD0 U2336 ( .I(n2313), .Z(n2312) );
  BUFFD0 U2337 ( .I(n2314), .Z(n2313) );
  BUFFD0 U2338 ( .I(n2315), .Z(n2314) );
  BUFFD0 U2339 ( .I(n2316), .Z(n2315) );
  BUFFD0 U2340 ( .I(n2317), .Z(n2316) );
  BUFFD0 U2341 ( .I(n2318), .Z(n2317) );
  BUFFD0 U2342 ( .I(n2319), .Z(n2318) );
  BUFFD0 U2343 ( .I(n2320), .Z(n2319) );
  BUFFD0 U2344 ( .I(n2321), .Z(n2320) );
  BUFFD0 U2345 ( .I(n2322), .Z(n2321) );
  BUFFD0 U2346 ( .I(n2323), .Z(n2322) );
  BUFFD0 U2347 ( .I(n2324), .Z(n2323) );
  BUFFD0 U2348 ( .I(n2325), .Z(n2324) );
  BUFFD0 U2349 ( .I(n2326), .Z(n2325) );
  BUFFD0 U2350 ( .I(n2327), .Z(n2326) );
  BUFFD0 U2351 ( .I(n2328), .Z(n2327) );
  BUFFD0 U2352 ( .I(n2329), .Z(n2328) );
  BUFFD0 U2353 ( .I(n2330), .Z(n2329) );
  BUFFD0 U2354 ( .I(n2331), .Z(n2330) );
  BUFFD0 U2355 ( .I(n2332), .Z(n2331) );
  BUFFD0 U2356 ( .I(n2333), .Z(n2332) );
  BUFFD0 U2357 ( .I(n2334), .Z(n2333) );
  BUFFD0 U2358 ( .I(n2335), .Z(n2334) );
  BUFFD0 U2359 ( .I(n2336), .Z(n2335) );
  BUFFD0 U2360 ( .I(n2337), .Z(n2336) );
  BUFFD0 U2361 ( .I(n2338), .Z(n2337) );
  BUFFD0 U2362 ( .I(n2339), .Z(n2338) );
  BUFFD0 U2363 ( .I(n2340), .Z(n2339) );
  BUFFD0 U2364 ( .I(n2341), .Z(n2340) );
  BUFFD0 U2365 ( .I(n2342), .Z(n2341) );
  BUFFD0 U2366 ( .I(n2343), .Z(n2342) );
  BUFFD0 U2367 ( .I(n2344), .Z(n2343) );
  BUFFD0 U2368 ( .I(n2345), .Z(n2344) );
  BUFFD0 U2369 ( .I(n2346), .Z(n2345) );
  BUFFD0 U2370 ( .I(n2347), .Z(n2346) );
  BUFFD0 U2371 ( .I(n2348), .Z(n2347) );
  BUFFD0 U2372 ( .I(n2349), .Z(n2348) );
  BUFFD0 U2373 ( .I(n2350), .Z(n2349) );
  BUFFD0 U2374 ( .I(n2351), .Z(n2350) );
  BUFFD0 U2375 ( .I(n2352), .Z(n2351) );
  BUFFD0 U2376 ( .I(n2353), .Z(n2352) );
  BUFFD0 U2377 ( .I(n2354), .Z(n2353) );
  BUFFD0 U2378 ( .I(n2355), .Z(n2354) );
  BUFFD0 U2379 ( .I(n2356), .Z(n2355) );
  BUFFD0 U2380 ( .I(n2357), .Z(n2356) );
  BUFFD0 U2381 ( .I(n2358), .Z(n2357) );
  BUFFD0 U2382 ( .I(n2359), .Z(n2358) );
  BUFFD0 U2383 ( .I(n2707), .Z(n2359) );
  BUFFD0 U2384 ( .I(n2364), .Z(n2360) );
  BUFFD0 U2385 ( .I(n2675), .Z(n2361) );
  BUFFD0 U2386 ( .I(n2361), .Z(n2362) );
  BUFFD0 U2387 ( .I(n2362), .Z(n2363) );
  BUFFD0 U2388 ( .I(n2365), .Z(n2364) );
  BUFFD0 U2389 ( .I(n2366), .Z(n2365) );
  BUFFD0 U2390 ( .I(n2367), .Z(n2366) );
  BUFFD0 U2391 ( .I(n2368), .Z(n2367) );
  BUFFD0 U2392 ( .I(n2369), .Z(n2368) );
  BUFFD0 U2393 ( .I(n2370), .Z(n2369) );
  BUFFD0 U2394 ( .I(n2371), .Z(n2370) );
  BUFFD0 U2395 ( .I(n2372), .Z(n2371) );
  BUFFD0 U2396 ( .I(n2373), .Z(n2372) );
  BUFFD0 U2397 ( .I(n2374), .Z(n2373) );
  BUFFD0 U2398 ( .I(n2375), .Z(n2374) );
  BUFFD0 U2399 ( .I(n2376), .Z(n2375) );
  BUFFD0 U2400 ( .I(n2377), .Z(n2376) );
  BUFFD0 U2401 ( .I(n2378), .Z(n2377) );
  BUFFD0 U2402 ( .I(n2379), .Z(n2378) );
  BUFFD0 U2403 ( .I(n2380), .Z(n2379) );
  BUFFD0 U2404 ( .I(n2381), .Z(n2380) );
  BUFFD0 U2405 ( .I(n2382), .Z(n2381) );
  BUFFD0 U2406 ( .I(n2383), .Z(n2382) );
  BUFFD0 U2407 ( .I(n2384), .Z(n2383) );
  BUFFD0 U2408 ( .I(n2385), .Z(n2384) );
  BUFFD0 U2409 ( .I(n2386), .Z(n2385) );
  BUFFD0 U2410 ( .I(n2387), .Z(n2386) );
  BUFFD0 U2411 ( .I(n2388), .Z(n2387) );
  BUFFD0 U2412 ( .I(n2389), .Z(n2388) );
  BUFFD0 U2413 ( .I(n2390), .Z(n2389) );
  BUFFD0 U2414 ( .I(n2391), .Z(n2390) );
  BUFFD0 U2415 ( .I(n2392), .Z(n2391) );
  BUFFD0 U2416 ( .I(n2393), .Z(n2392) );
  BUFFD0 U2417 ( .I(n2394), .Z(n2393) );
  BUFFD0 U2418 ( .I(n2395), .Z(n2394) );
  BUFFD0 U2419 ( .I(n2396), .Z(n2395) );
  BUFFD0 U2420 ( .I(n2397), .Z(n2396) );
  BUFFD0 U2421 ( .I(n2398), .Z(n2397) );
  BUFFD0 U2422 ( .I(n2399), .Z(n2398) );
  BUFFD0 U2423 ( .I(n2400), .Z(n2399) );
  BUFFD0 U2424 ( .I(n2401), .Z(n2400) );
  BUFFD0 U2425 ( .I(n2402), .Z(n2401) );
  BUFFD0 U2426 ( .I(n2403), .Z(n2402) );
  BUFFD0 U2427 ( .I(n2404), .Z(n2403) );
  BUFFD0 U2428 ( .I(n2405), .Z(n2404) );
  BUFFD0 U2429 ( .I(n2406), .Z(n2405) );
  BUFFD0 U2430 ( .I(n2407), .Z(n2406) );
  BUFFD0 U2431 ( .I(n2408), .Z(n2407) );
  BUFFD0 U2432 ( .I(n2409), .Z(n2408) );
  BUFFD0 U2433 ( .I(n2410), .Z(n2409) );
  BUFFD0 U2434 ( .I(n2411), .Z(n2410) );
  BUFFD0 U2435 ( .I(n2412), .Z(n2411) );
  BUFFD0 U2436 ( .I(n2413), .Z(n2412) );
  BUFFD0 U2437 ( .I(n2414), .Z(n2413) );
  BUFFD0 U2438 ( .I(n2415), .Z(n2414) );
  BUFFD0 U2439 ( .I(n2416), .Z(n2415) );
  BUFFD0 U2440 ( .I(n2417), .Z(n2416) );
  BUFFD0 U2441 ( .I(n2418), .Z(n2417) );
  BUFFD0 U2442 ( .I(n2363), .Z(n2418) );
  BUFFD0 U2443 ( .I(n2423), .Z(n2419) );
  BUFFD0 U2444 ( .I(n2673), .Z(n2420) );
  BUFFD0 U2445 ( .I(n2420), .Z(n2421) );
  BUFFD0 U2446 ( .I(n2421), .Z(n2422) );
  BUFFD0 U2447 ( .I(n2424), .Z(n2423) );
  BUFFD0 U2448 ( .I(n2425), .Z(n2424) );
  BUFFD0 U2449 ( .I(n2426), .Z(n2425) );
  BUFFD0 U2450 ( .I(n2427), .Z(n2426) );
  BUFFD0 U2451 ( .I(n2428), .Z(n2427) );
  BUFFD0 U2452 ( .I(n2429), .Z(n2428) );
  BUFFD0 U2453 ( .I(n2430), .Z(n2429) );
  BUFFD0 U2454 ( .I(n2431), .Z(n2430) );
  BUFFD0 U2455 ( .I(n2432), .Z(n2431) );
  BUFFD0 U2456 ( .I(n2433), .Z(n2432) );
  BUFFD0 U2457 ( .I(n2434), .Z(n2433) );
  BUFFD0 U2458 ( .I(n2435), .Z(n2434) );
  BUFFD0 U2459 ( .I(n2436), .Z(n2435) );
  BUFFD0 U2460 ( .I(n2437), .Z(n2436) );
  BUFFD0 U2461 ( .I(n2438), .Z(n2437) );
  BUFFD0 U2462 ( .I(n2439), .Z(n2438) );
  BUFFD0 U2463 ( .I(n2440), .Z(n2439) );
  BUFFD0 U2464 ( .I(n2441), .Z(n2440) );
  BUFFD0 U2465 ( .I(n2442), .Z(n2441) );
  BUFFD0 U2466 ( .I(n2443), .Z(n2442) );
  BUFFD0 U2467 ( .I(n2444), .Z(n2443) );
  BUFFD0 U2468 ( .I(n2445), .Z(n2444) );
  BUFFD0 U2469 ( .I(n2446), .Z(n2445) );
  BUFFD0 U2470 ( .I(n2447), .Z(n2446) );
  BUFFD0 U2471 ( .I(n2448), .Z(n2447) );
  BUFFD0 U2472 ( .I(n2449), .Z(n2448) );
  BUFFD0 U2473 ( .I(n2450), .Z(n2449) );
  BUFFD0 U2474 ( .I(n2451), .Z(n2450) );
  BUFFD0 U2475 ( .I(n2452), .Z(n2451) );
  BUFFD0 U2476 ( .I(n2453), .Z(n2452) );
  BUFFD0 U2477 ( .I(n2454), .Z(n2453) );
  BUFFD0 U2478 ( .I(n2455), .Z(n2454) );
  BUFFD0 U2479 ( .I(n2456), .Z(n2455) );
  BUFFD0 U2480 ( .I(n2457), .Z(n2456) );
  BUFFD0 U2481 ( .I(n2458), .Z(n2457) );
  BUFFD0 U2482 ( .I(n2459), .Z(n2458) );
  BUFFD0 U2483 ( .I(n2460), .Z(n2459) );
  BUFFD0 U2484 ( .I(n2461), .Z(n2460) );
  BUFFD0 U2485 ( .I(n2462), .Z(n2461) );
  BUFFD0 U2486 ( .I(n2463), .Z(n2462) );
  BUFFD0 U2487 ( .I(n2464), .Z(n2463) );
  BUFFD0 U2488 ( .I(n2465), .Z(n2464) );
  BUFFD0 U2489 ( .I(n2466), .Z(n2465) );
  BUFFD0 U2490 ( .I(n2467), .Z(n2466) );
  BUFFD0 U2491 ( .I(n2468), .Z(n2467) );
  BUFFD0 U2492 ( .I(n2469), .Z(n2468) );
  BUFFD0 U2493 ( .I(n2470), .Z(n2469) );
  BUFFD0 U2494 ( .I(n2471), .Z(n2470) );
  BUFFD0 U2495 ( .I(n2472), .Z(n2471) );
  BUFFD0 U2496 ( .I(n2473), .Z(n2472) );
  BUFFD0 U2497 ( .I(n2474), .Z(n2473) );
  BUFFD0 U2498 ( .I(n2475), .Z(n2474) );
  BUFFD0 U2499 ( .I(n2476), .Z(n2475) );
  BUFFD0 U2500 ( .I(n2477), .Z(n2476) );
  BUFFD0 U2501 ( .I(n2422), .Z(n2477) );
  BUFFD0 U2502 ( .I(n2482), .Z(n2478) );
  BUFFD0 U2503 ( .I(N81), .Z(n2479) );
  BUFFD0 U2504 ( .I(n2479), .Z(n2480) );
  BUFFD0 U2505 ( .I(n2480), .Z(n2481) );
  BUFFD0 U2506 ( .I(n2483), .Z(n2482) );
  BUFFD0 U2507 ( .I(n2484), .Z(n2483) );
  BUFFD0 U2508 ( .I(n2485), .Z(n2484) );
  BUFFD0 U2509 ( .I(n2486), .Z(n2485) );
  BUFFD0 U2510 ( .I(n2487), .Z(n2486) );
  BUFFD0 U2511 ( .I(n2488), .Z(n2487) );
  BUFFD0 U2512 ( .I(n2489), .Z(n2488) );
  BUFFD0 U2513 ( .I(n2490), .Z(n2489) );
  BUFFD0 U2514 ( .I(n2491), .Z(n2490) );
  BUFFD0 U2515 ( .I(n2492), .Z(n2491) );
  BUFFD0 U2516 ( .I(n2493), .Z(n2492) );
  BUFFD0 U2517 ( .I(n2494), .Z(n2493) );
  BUFFD0 U2518 ( .I(n2495), .Z(n2494) );
  BUFFD0 U2519 ( .I(n2496), .Z(n2495) );
  BUFFD0 U2520 ( .I(n2497), .Z(n2496) );
  BUFFD0 U2521 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2522 ( .I(n2499), .Z(n2498) );
  BUFFD0 U2523 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2524 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2525 ( .I(n2502), .Z(n2501) );
  BUFFD0 U2526 ( .I(n2503), .Z(n2502) );
  BUFFD0 U2527 ( .I(n2504), .Z(n2503) );
  BUFFD0 U2528 ( .I(n2505), .Z(n2504) );
  BUFFD0 U2529 ( .I(n2506), .Z(n2505) );
  BUFFD0 U2530 ( .I(n2507), .Z(n2506) );
  BUFFD0 U2531 ( .I(n2508), .Z(n2507) );
  BUFFD0 U2532 ( .I(n2509), .Z(n2508) );
  BUFFD0 U2533 ( .I(n2510), .Z(n2509) );
  BUFFD0 U2534 ( .I(n2511), .Z(n2510) );
  BUFFD0 U2535 ( .I(n2512), .Z(n2511) );
  BUFFD0 U2536 ( .I(n2513), .Z(n2512) );
  BUFFD0 U2537 ( .I(n2514), .Z(n2513) );
  BUFFD0 U2538 ( .I(n2515), .Z(n2514) );
  BUFFD0 U2539 ( .I(n2516), .Z(n2515) );
  BUFFD0 U2540 ( .I(n2517), .Z(n2516) );
  BUFFD0 U2541 ( .I(n2518), .Z(n2517) );
  BUFFD0 U2542 ( .I(n2519), .Z(n2518) );
  BUFFD0 U2543 ( .I(n2520), .Z(n2519) );
  BUFFD0 U2544 ( .I(n2521), .Z(n2520) );
  BUFFD0 U2545 ( .I(n2522), .Z(n2521) );
  BUFFD0 U2546 ( .I(n2523), .Z(n2522) );
  BUFFD0 U2547 ( .I(n2524), .Z(n2523) );
  BUFFD0 U2548 ( .I(n2525), .Z(n2524) );
  BUFFD0 U2549 ( .I(n2526), .Z(n2525) );
  BUFFD0 U2550 ( .I(n2527), .Z(n2526) );
  BUFFD0 U2551 ( .I(n2528), .Z(n2527) );
  BUFFD0 U2552 ( .I(n2529), .Z(n2528) );
  BUFFD0 U2553 ( .I(n2530), .Z(n2529) );
  BUFFD0 U2554 ( .I(n2531), .Z(n2530) );
  BUFFD0 U2555 ( .I(n2532), .Z(n2531) );
  BUFFD0 U2556 ( .I(n2533), .Z(n2532) );
  BUFFD0 U2557 ( .I(n2534), .Z(n2533) );
  BUFFD0 U2558 ( .I(n2535), .Z(n2534) );
  BUFFD0 U2559 ( .I(n2536), .Z(n2535) );
  BUFFD0 U2560 ( .I(n2676), .Z(n2536) );
  BUFFD0 U2561 ( .I(N75), .Z(n2537) );
  BUFFD0 U2562 ( .I(N68), .Z(n2538) );
  BUFFD0 U2563 ( .I(N74), .Z(n2539) );
  BUFFD0 U2564 ( .I(N82), .Z(n2540) );
  BUFFD0 U2565 ( .I(n2540), .Z(n2541) );
  BUFFD0 U2566 ( .I(n2543), .Z(n2542) );
  BUFFD0 U2567 ( .I(n2544), .Z(n2543) );
  BUFFD0 U2568 ( .I(n2545), .Z(n2544) );
  BUFFD0 U2569 ( .I(n2546), .Z(n2545) );
  BUFFD0 U2570 ( .I(n2547), .Z(n2546) );
  BUFFD0 U2571 ( .I(n2548), .Z(n2547) );
  BUFFD0 U2572 ( .I(n2549), .Z(n2548) );
  BUFFD0 U2573 ( .I(n2550), .Z(n2549) );
  BUFFD0 U2574 ( .I(n2551), .Z(n2550) );
  BUFFD0 U2575 ( .I(n2552), .Z(n2551) );
  BUFFD0 U2576 ( .I(n2553), .Z(n2552) );
  BUFFD0 U2577 ( .I(n2554), .Z(n2553) );
  BUFFD0 U2578 ( .I(n2555), .Z(n2554) );
  BUFFD0 U2579 ( .I(n2556), .Z(n2555) );
  BUFFD0 U2580 ( .I(n2557), .Z(n2556) );
  BUFFD0 U2581 ( .I(n2558), .Z(n2557) );
  BUFFD0 U2582 ( .I(n2559), .Z(n2558) );
  BUFFD0 U2583 ( .I(n2560), .Z(n2559) );
  BUFFD0 U2584 ( .I(n2561), .Z(n2560) );
  BUFFD0 U2585 ( .I(n2562), .Z(n2561) );
  BUFFD0 U2586 ( .I(n2563), .Z(n2562) );
  BUFFD0 U2587 ( .I(n2564), .Z(n2563) );
  BUFFD0 U2588 ( .I(n2565), .Z(n2564) );
  BUFFD0 U2589 ( .I(n2566), .Z(n2565) );
  BUFFD0 U2590 ( .I(n2567), .Z(n2566) );
  BUFFD0 U2591 ( .I(n2568), .Z(n2567) );
  BUFFD0 U2592 ( .I(n2569), .Z(n2568) );
  BUFFD0 U2593 ( .I(n2570), .Z(n2569) );
  BUFFD0 U2594 ( .I(n2571), .Z(n2570) );
  BUFFD0 U2595 ( .I(n2572), .Z(n2571) );
  BUFFD0 U2596 ( .I(n2573), .Z(n2572) );
  BUFFD0 U2597 ( .I(n2574), .Z(n2573) );
  BUFFD0 U2598 ( .I(n2575), .Z(n2574) );
  BUFFD0 U2599 ( .I(n2576), .Z(n2575) );
  BUFFD0 U2600 ( .I(n2577), .Z(n2576) );
  BUFFD0 U2601 ( .I(n2578), .Z(n2577) );
  BUFFD0 U2602 ( .I(n2579), .Z(n2578) );
  BUFFD0 U2603 ( .I(n2580), .Z(n2579) );
  BUFFD0 U2604 ( .I(n2581), .Z(n2580) );
  BUFFD0 U2605 ( .I(n2582), .Z(n2581) );
  BUFFD0 U2606 ( .I(n2583), .Z(n2582) );
  BUFFD0 U2607 ( .I(n2584), .Z(n2583) );
  BUFFD0 U2608 ( .I(n2585), .Z(n2584) );
  BUFFD0 U2609 ( .I(n2586), .Z(n2585) );
  BUFFD0 U2610 ( .I(n2587), .Z(n2586) );
  BUFFD0 U2611 ( .I(n2588), .Z(n2587) );
  BUFFD0 U2612 ( .I(n2589), .Z(n2588) );
  BUFFD0 U2613 ( .I(n2590), .Z(n2589) );
  BUFFD0 U2614 ( .I(n2591), .Z(n2590) );
  BUFFD0 U2615 ( .I(n2592), .Z(n2591) );
  BUFFD0 U2616 ( .I(n2662), .Z(n2592) );
  BUFFD0 U2617 ( .I(n1319), .Z(n2593) );
  BUFFD0 U2618 ( .I(n2617), .Z(n2594) );
  BUFFD0 U2619 ( .I(n2189), .Z(n2595) );
  BUFFD0 U2620 ( .I(N80), .Z(n2596) );
  BUFFD0 U2621 ( .I(N79), .Z(n2597) );
  BUFFD0 U2622 ( .I(n1644), .Z(n2598) );
  BUFFD0 U2623 ( .I(n2481), .Z(n2599) );
  BUFFD0 U2624 ( .I(n1385), .Z(n2600) );
  BUFFD0 U2625 ( .I(n1253), .Z(n2601) );
  BUFFD0 U2626 ( .I(n2623), .Z(n2602) );
  BUFFD0 U2627 ( .I(N65), .Z(n2603) );
  BUFFD0 U2628 ( .I(n1451), .Z(n2604) );
  BUFFD0 U2629 ( .I(n2248), .Z(n2605) );
  BUFFD0 U2630 ( .I(n1955), .Z(n2606) );
  BUFFD0 U2631 ( .I(N73), .Z(n2607) );
  BUFFD0 U2632 ( .I(n1640), .Z(n2608) );
  BUFFD0 U2633 ( .I(N69), .Z(n2609) );
  BUFFD0 U2634 ( .I(n2307), .Z(n2610) );
  BUFFD0 U2635 ( .I(n1890), .Z(n2611) );
  BUFFD0 U2636 ( .I(n1122), .Z(n2612) );
  BUFFD0 U2637 ( .I(n2537), .Z(n2613) );
  BUFFD0 U2638 ( .I(n2538), .Z(n2614) );
  BUFFD0 U2639 ( .I(n1894), .Z(n2615) );
  BUFFD0 U2640 ( .I(n2539), .Z(n2616) );
  BUFFD0 U2641 ( .I(n1187), .Z(n2617) );
  BUFFD0 U2642 ( .I(n2595), .Z(n2618) );
  BUFFD0 U2643 ( .I(n2596), .Z(n2619) );
  BUFFD0 U2644 ( .I(n2597), .Z(n2620) );
  BUFFD0 U2645 ( .I(n2598), .Z(n2621) );
  BUFFD0 U2646 ( .I(n2599), .Z(n2622) );
  BUFFD0 U2647 ( .I(n2641), .Z(n2623) );
  BUFFD0 U2648 ( .I(n2642), .Z(n2624) );
  BUFFD0 U2649 ( .I(n2605), .Z(n2625) );
  BUFFD0 U2650 ( .I(n2606), .Z(n2626) );
  BUFFD0 U2651 ( .I(n2607), .Z(n2627) );
  BUFFD0 U2652 ( .I(n2646), .Z(n2628) );
  BUFFD0 U2653 ( .I(n2647), .Z(n2629) );
  BUFFD0 U2654 ( .I(n2610), .Z(n2630) );
  BUFFD0 U2655 ( .I(n2649), .Z(n2631) );
  BUFFD0 U2656 ( .I(n2613), .Z(n2632) );
  BUFFD0 U2657 ( .I(n2651), .Z(n2633) );
  BUFFD0 U2658 ( .I(n2615), .Z(n2634) );
  BUFFD0 U2659 ( .I(n2616), .Z(n2635) );
  BUFFD0 U2660 ( .I(n2618), .Z(n2636) );
  BUFFD0 U2661 ( .I(n2619), .Z(n2637) );
  BUFFD0 U2662 ( .I(n2620), .Z(n2638) );
  BUFFD0 U2663 ( .I(n2657), .Z(n2639) );
  BUFFD0 U2664 ( .I(n2622), .Z(n2640) );
  BUFFD0 U2665 ( .I(N64), .Z(n2641) );
  BUFFD0 U2666 ( .I(n2659), .Z(n2642) );
  BUFFD0 U2667 ( .I(n2625), .Z(n2643) );
  BUFFD0 U2668 ( .I(n2626), .Z(n2644) );
  BUFFD0 U2669 ( .I(n2627), .Z(n2645) );
  BUFFD0 U2670 ( .I(n2664), .Z(n2646) );
  BUFFD0 U2671 ( .I(n2665), .Z(n2647) );
  BUFFD0 U2672 ( .I(n2630), .Z(n2648) );
  BUFFD0 U2673 ( .I(n2667), .Z(n2649) );
  BUFFD0 U2674 ( .I(n2632), .Z(n2650) );
  BUFFD0 U2675 ( .I(n2668), .Z(n2651) );
  BUFFD0 U2676 ( .I(n2634), .Z(n2652) );
  BUFFD0 U2677 ( .I(n2635), .Z(n2653) );
  BUFFD0 U2678 ( .I(n2636), .Z(n2654) );
  BUFFD0 U2679 ( .I(n2637), .Z(n2655) );
  BUFFD0 U2680 ( .I(n2638), .Z(n2656) );
  BUFFD0 U2681 ( .I(n2674), .Z(n2657) );
  BUFFD0 U2682 ( .I(n2640), .Z(n2658) );
  BUFFD0 U2683 ( .I(n2603), .Z(n2659) );
  BUFFD0 U2684 ( .I(n2643), .Z(n2660) );
  BUFFD0 U2685 ( .I(n2644), .Z(n2661) );
  BUFFD0 U2686 ( .I(n2541), .Z(n2662) );
  BUFFD0 U2687 ( .I(n2645), .Z(n2663) );
  BUFFD0 U2688 ( .I(n2608), .Z(n2664) );
  BUFFD0 U2689 ( .I(n2609), .Z(n2665) );
  BUFFD0 U2690 ( .I(n2648), .Z(n2666) );
  BUFFD0 U2691 ( .I(n2611), .Z(n2667) );
  BUFFD0 U2692 ( .I(n2614), .Z(n2668) );
  BUFFD0 U2693 ( .I(n2650), .Z(n2669) );
  BUFFD0 U2694 ( .I(n2682), .Z(n2670) );
  BUFFD0 U2695 ( .I(n2683), .Z(n2671) );
  BUFFD0 U2696 ( .I(n2654), .Z(n2672) );
  BUFFD0 U2697 ( .I(n2685), .Z(n2673) );
  BUFFD0 U2698 ( .I(n2621), .Z(n2674) );
  BUFFD0 U2699 ( .I(n2686), .Z(n2675) );
  BUFFD0 U2700 ( .I(n2687), .Z(n2676) );
  BUFFD0 U2701 ( .I(n2688), .Z(n2677) );
  BUFFD0 U2702 ( .I(n2661), .Z(n2678) );
  BUFFD0 U2703 ( .I(n2663), .Z(n2679) );
  BUFFD0 U2704 ( .I(n2666), .Z(n2680) );
  BUFFD0 U2705 ( .I(n2693), .Z(n2681) );
  BUFFD0 U2706 ( .I(n2692), .Z(n2682) );
  BUFFD0 U2707 ( .I(n2694), .Z(n2683) );
  BUFFD0 U2708 ( .I(n2697), .Z(n2684) );
  BUFFD0 U2709 ( .I(n2698), .Z(n2687) );
  BUFFD0 U2710 ( .I(n2699), .Z(n2688) );
  BUFFD0 U2711 ( .I(n2678), .Z(n2689) );
  BUFFD0 U2712 ( .I(n2679), .Z(n2690) );
  BUFFD0 U2713 ( .I(n2680), .Z(n2691) );
  BUFFD0 U2714 ( .I(n2653), .Z(n2692) );
  BUFFD0 U2715 ( .I(n2703), .Z(n2693) );
  BUFFD0 U2716 ( .I(n2652), .Z(n2694) );
  BUFFD0 U2717 ( .I(n2655), .Z(n2695) );
  BUFFD0 U2718 ( .I(n2656), .Z(n2696) );
  BUFFD0 U2719 ( .I(n2704), .Z(n2697) );
  BUFFD0 U2720 ( .I(n2658), .Z(n2698) );
  BUFFD0 U2721 ( .I(n2660), .Z(n2699) );
  BUFFD0 U2722 ( .I(n2705), .Z(n2700) );
  BUFFD0 U2723 ( .I(n2690), .Z(n2701) );
  BUFFD0 U2724 ( .I(n2691), .Z(n2702) );
  BUFFD0 U2725 ( .I(n2669), .Z(n2703) );
  BUFFD0 U2726 ( .I(n2672), .Z(n2704) );
  BUFFD0 U2727 ( .I(n2708), .Z(n2705) );
  BUFFD0 U2728 ( .I(n2709), .Z(n2706) );
  BUFFD0 U2729 ( .I(n2710), .Z(n2707) );
  BUFFD0 U2730 ( .I(n2689), .Z(n2708) );
  BUFFD0 U2731 ( .I(n2711), .Z(n2709) );
  BUFFD0 U2732 ( .I(n2712), .Z(n2710) );
  BUFFD0 U2733 ( .I(n2701), .Z(n2711) );
  BUFFD0 U2734 ( .I(n2702), .Z(n2712) );
  BUFFD0 U2735 ( .I(n3057), .Z(n2713) );
  BUFFD0 U2736 ( .I(n2715), .Z(n2714) );
  BUFFD0 U2737 ( .I(n2716), .Z(n2715) );
  BUFFD0 U2738 ( .I(n2717), .Z(n2716) );
  BUFFD0 U2739 ( .I(n2718), .Z(n2717) );
  BUFFD0 U2740 ( .I(n2719), .Z(n2718) );
  BUFFD0 U2741 ( .I(n2720), .Z(n2719) );
  BUFFD0 U2742 ( .I(n2721), .Z(n2720) );
  BUFFD0 U2743 ( .I(n2722), .Z(n2721) );
  BUFFD0 U2744 ( .I(n2723), .Z(n2722) );
  BUFFD0 U2745 ( .I(n2724), .Z(n2723) );
  BUFFD0 U2746 ( .I(n2725), .Z(n2724) );
  BUFFD0 U2747 ( .I(n2726), .Z(n2725) );
  BUFFD0 U2748 ( .I(n2727), .Z(n2726) );
  BUFFD0 U2749 ( .I(n2728), .Z(n2727) );
  BUFFD0 U2750 ( .I(n2729), .Z(n2728) );
  BUFFD0 U2751 ( .I(n2730), .Z(n2729) );
  BUFFD0 U2752 ( .I(n2731), .Z(n2730) );
  BUFFD0 U2753 ( .I(n2732), .Z(n2731) );
  BUFFD0 U2754 ( .I(n2733), .Z(n2732) );
  BUFFD0 U2755 ( .I(n2734), .Z(n2733) );
  BUFFD0 U2756 ( .I(n2735), .Z(n2734) );
  BUFFD0 U2757 ( .I(n2736), .Z(n2735) );
  BUFFD0 U2758 ( .I(n2737), .Z(n2736) );
  BUFFD0 U2759 ( .I(n2738), .Z(n2737) );
  BUFFD0 U2760 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2761 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2762 ( .I(n2741), .Z(n2740) );
  BUFFD0 U2763 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2764 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2765 ( .I(n2744), .Z(n2743) );
  BUFFD0 U2766 ( .I(n2745), .Z(n2744) );
  BUFFD0 U2767 ( .I(n2746), .Z(n2745) );
  BUFFD0 U2768 ( .I(n2747), .Z(n2746) );
  BUFFD0 U2769 ( .I(n2748), .Z(n2747) );
  BUFFD0 U2770 ( .I(n2749), .Z(n2748) );
  BUFFD0 U2771 ( .I(n2750), .Z(n2749) );
  BUFFD0 U2772 ( .I(n2751), .Z(n2750) );
  BUFFD0 U2773 ( .I(n2752), .Z(n2751) );
  BUFFD0 U2774 ( .I(n2753), .Z(n2752) );
  BUFFD0 U2775 ( .I(n2754), .Z(n2753) );
  BUFFD0 U2776 ( .I(n2755), .Z(n2754) );
  BUFFD0 U2777 ( .I(n2756), .Z(n2755) );
  BUFFD0 U2778 ( .I(n2757), .Z(n2756) );
  BUFFD0 U2779 ( .I(n2758), .Z(n2757) );
  BUFFD0 U2780 ( .I(n2759), .Z(n2758) );
  BUFFD0 U2781 ( .I(n2760), .Z(n2759) );
  BUFFD0 U2782 ( .I(n2761), .Z(n2760) );
  BUFFD0 U2783 ( .I(n2762), .Z(n2761) );
  BUFFD0 U2784 ( .I(n2763), .Z(n2762) );
  BUFFD0 U2785 ( .I(n2764), .Z(n2763) );
  BUFFD0 U2786 ( .I(n2765), .Z(n2764) );
  BUFFD0 U2787 ( .I(n2766), .Z(n2765) );
  BUFFD0 U2788 ( .I(n2767), .Z(n2766) );
  BUFFD0 U2789 ( .I(Read), .Z(n2767) );
  CKAN2D0 U2790 ( .A1(Dreadyr), .A2(ChipEna), .Z(Dready) );
  BUFFD1 U2791 ( .I(n3103), .Z(n3067) );
  BUFFD1 U2792 ( .I(n3105), .Z(n3068) );
  BUFFD1 U2793 ( .I(n3105), .Z(n3069) );
  BUFFD1 U2794 ( .I(n3104), .Z(n3070) );
  BUFFD1 U2795 ( .I(n3104), .Z(n3071) );
  BUFFD1 U2796 ( .I(n3103), .Z(n3072) );
  BUFFD1 U2797 ( .I(n3103), .Z(n3073) );
  BUFFD1 U2798 ( .I(n3101), .Z(n3074) );
  BUFFD1 U2799 ( .I(n3101), .Z(n3075) );
  BUFFD1 U2800 ( .I(n3104), .Z(n3076) );
  BUFFD1 U2801 ( .I(n3105), .Z(n3077) );
  BUFFD1 U2802 ( .I(n3100), .Z(n3078) );
  BUFFD1 U2803 ( .I(n3100), .Z(n3079) );
  BUFFD1 U2804 ( .I(n3110), .Z(n3080) );
  BUFFD1 U2805 ( .I(n3099), .Z(n3081) );
  BUFFD1 U2806 ( .I(n3098), .Z(n3082) );
  BUFFD1 U2807 ( .I(n3098), .Z(n3083) );
  BUFFD1 U2808 ( .I(n3097), .Z(n3084) );
  BUFFD1 U2809 ( .I(n3097), .Z(n3085) );
  BUFFD1 U2810 ( .I(n3096), .Z(n3086) );
  BUFFD1 U2811 ( .I(n3096), .Z(n3087) );
  BUFFD1 U2812 ( .I(n3097), .Z(n3088) );
  BUFFD1 U2813 ( .I(n3096), .Z(n3089) );
  BUFFD1 U2814 ( .I(n3095), .Z(n3090) );
  BUFFD1 U2815 ( .I(n3095), .Z(n3091) );
  BUFFD1 U2816 ( .I(n3095), .Z(n3092) );
  BUFFD1 U2817 ( .I(n3094), .Z(n3093) );
  BUFFD1 U2818 ( .I(n3094), .Z(n3062) );
  BUFFD1 U2819 ( .I(n3098), .Z(n3063) );
  BUFFD1 U2820 ( .I(n3103), .Z(n3064) );
  BUFFD1 U2821 ( .I(n3100), .Z(n3065) );
  BUFFD1 U2822 ( .I(n3094), .Z(n3066) );
  BUFFD1 U2823 ( .I(n3107), .Z(n3105) );
  BUFFD1 U2824 ( .I(n3107), .Z(n3104) );
  BUFFD1 U2825 ( .I(n3108), .Z(n3103) );
  BUFFD1 U2826 ( .I(n3113), .Z(n3102) );
  BUFFD1 U2827 ( .I(n3108), .Z(n3101) );
  BUFFD1 U2828 ( .I(n3095), .Z(n3100) );
  BUFFD1 U2829 ( .I(n3095), .Z(n3099) );
  BUFFD1 U2830 ( .I(n3106), .Z(n3098) );
  BUFFD1 U2831 ( .I(n3109), .Z(n3097) );
  BUFFD1 U2832 ( .I(n3109), .Z(n3096) );
  BUFFD1 U2833 ( .I(n3111), .Z(n3095) );
  BUFFD1 U2834 ( .I(n3110), .Z(n3094) );
  BUFFD1 U2835 ( .I(n3113), .Z(n3107) );
  BUFFD1 U2836 ( .I(n3113), .Z(n3108) );
  BUFFD1 U2837 ( .I(n3112), .Z(n3109) );
  BUFFD1 U2838 ( .I(n3111), .Z(n3110) );
  BUFFD1 U2839 ( .I(n3115), .Z(n3113) );
  BUFFD1 U2840 ( .I(n3115), .Z(n3112) );
  BUFFD1 U2841 ( .I(n3115), .Z(n3111) );
  BUFFD1 U2842 ( .I(n3114), .Z(n3106) );
  BUFFD1 U2843 ( .I(n3115), .Z(n3114) );
  INVD1 U2844 ( .I(Reset), .ZN(n3115) );
  BUFFD1 U2845 ( .I(n3045), .Z(n3024) );
  BUFFD1 U2846 ( .I(n3047), .Z(n3023) );
  BUFFD1 U2847 ( .I(n3025), .Z(n3022) );
  BUFFD1 U2848 ( .I(n3025), .Z(n3021) );
  BUFFD1 U2849 ( .I(n3026), .Z(n3020) );
  BUFFD1 U2850 ( .I(n3026), .Z(n3019) );
  BUFFD1 U2851 ( .I(n3027), .Z(n3018) );
  BUFFD1 U2852 ( .I(n3027), .Z(n3017) );
  BUFFD1 U2853 ( .I(n3028), .Z(n3016) );
  BUFFD1 U2854 ( .I(n3028), .Z(n3015) );
  BUFFD1 U2855 ( .I(n3029), .Z(n3014) );
  BUFFD1 U2856 ( .I(n3029), .Z(n3013) );
  BUFFD1 U2857 ( .I(n3030), .Z(n3012) );
  BUFFD1 U2858 ( .I(n3030), .Z(n3011) );
  BUFFD1 U2859 ( .I(n3031), .Z(n3010) );
  BUFFD1 U2860 ( .I(n3031), .Z(n3009) );
  BUFFD1 U2861 ( .I(n3032), .Z(n3008) );
  BUFFD1 U2862 ( .I(n3032), .Z(n3007) );
  BUFFD1 U2863 ( .I(n3033), .Z(n3006) );
  BUFFD1 U2864 ( .I(n3033), .Z(n3005) );
  BUFFD1 U2865 ( .I(n3034), .Z(n3004) );
  BUFFD1 U2866 ( .I(n3034), .Z(n3003) );
  BUFFD1 U2867 ( .I(n3035), .Z(n3002) );
  BUFFD1 U2868 ( .I(n3041), .Z(n3001) );
  BUFFD1 U2869 ( .I(n3036), .Z(n3000) );
  BUFFD1 U2870 ( .I(n3036), .Z(n2999) );
  BUFFD1 U2871 ( .I(n3037), .Z(n2998) );
  BUFFD1 U2872 ( .I(n3037), .Z(n2997) );
  BUFFD1 U2873 ( .I(n3038), .Z(n2996) );
  BUFFD1 U2874 ( .I(n3038), .Z(n2995) );
  BUFFD1 U2875 ( .I(n3039), .Z(n2994) );
  BUFFD1 U2876 ( .I(n3039), .Z(n2993) );
  BUFFD1 U2877 ( .I(n3040), .Z(n2992) );
  BUFFD1 U2878 ( .I(n3040), .Z(n2991) );
  BUFFD1 U2879 ( .I(n3041), .Z(n2990) );
  BUFFD1 U2880 ( .I(n3041), .Z(n2989) );
  BUFFD1 U2881 ( .I(n3042), .Z(n2988) );
  BUFFD1 U2882 ( .I(n3042), .Z(n2987) );
  BUFFD1 U2883 ( .I(n3043), .Z(n2986) );
  BUFFD1 U2884 ( .I(n3043), .Z(n2985) );
  BUFFD1 U2885 ( .I(n3044), .Z(n2984) );
  BUFFD1 U2886 ( .I(n3044), .Z(n2983) );
  INVD1 U2887 ( .I(n185), .ZN(n2976) );
  INVD1 U2888 ( .I(n185), .ZN(n2975) );
  INVD1 U2889 ( .I(n193), .ZN(n2959) );
  BUFFD1 U2890 ( .I(n3045), .Z(n2982) );
  BUFFD1 U2891 ( .I(n3046), .Z(n3045) );
  BUFFD1 U2892 ( .I(n3052), .Z(n3025) );
  BUFFD1 U2893 ( .I(n3052), .Z(n3026) );
  BUFFD1 U2894 ( .I(n3052), .Z(n3027) );
  BUFFD1 U2895 ( .I(n3051), .Z(n3028) );
  BUFFD1 U2896 ( .I(n3051), .Z(n3029) );
  BUFFD1 U2897 ( .I(n3051), .Z(n3030) );
  BUFFD1 U2898 ( .I(n3050), .Z(n3031) );
  BUFFD1 U2899 ( .I(n3050), .Z(n3032) );
  BUFFD1 U2900 ( .I(n3050), .Z(n3033) );
  BUFFD1 U2901 ( .I(n3049), .Z(n3034) );
  BUFFD1 U2902 ( .I(n3049), .Z(n3035) );
  BUFFD1 U2903 ( .I(n3031), .Z(n3036) );
  BUFFD1 U2904 ( .I(n3048), .Z(n3037) );
  BUFFD1 U2905 ( .I(n3026), .Z(n3038) );
  BUFFD1 U2906 ( .I(n3025), .Z(n3039) );
  BUFFD1 U2907 ( .I(n3047), .Z(n3040) );
  BUFFD1 U2908 ( .I(n3047), .Z(n3041) );
  BUFFD1 U2909 ( .I(n3047), .Z(n3042) );
  BUFFD1 U2910 ( .I(n3046), .Z(n3043) );
  BUFFD1 U2911 ( .I(n3046), .Z(n3044) );
  INVD1 U2912 ( .I(n196), .ZN(n2974) );
  INVD1 U2913 ( .I(n194), .ZN(n2972) );
  INVD1 U2914 ( .I(n194), .ZN(n2971) );
  INVD1 U2915 ( .I(n191), .ZN(n2970) );
  INVD1 U2916 ( .I(n191), .ZN(n2969) );
  INVD1 U2917 ( .I(n192), .ZN(n2968) );
  INVD1 U2918 ( .I(n192), .ZN(n2967) );
  INVD1 U2919 ( .I(n195), .ZN(n2966) );
  INVD1 U2920 ( .I(n195), .ZN(n2965) );
  INVD1 U2921 ( .I(n198), .ZN(n2964) );
  INVD1 U2922 ( .I(n198), .ZN(n2963) );
  INVD1 U2923 ( .I(n2961), .ZN(n2962) );
  INVD1 U2924 ( .I(n190), .ZN(n2957) );
  INVD1 U2925 ( .I(n190), .ZN(n2956) );
  INVD1 U2926 ( .I(n188), .ZN(n2955) );
  INVD1 U2927 ( .I(n188), .ZN(n2954) );
  INVD1 U2928 ( .I(n186), .ZN(n2953) );
  INVD1 U2929 ( .I(n186), .ZN(n2952) );
  INVD1 U2930 ( .I(n187), .ZN(n2951) );
  INVD1 U2931 ( .I(n187), .ZN(n2950) );
  INVD1 U2932 ( .I(n189), .ZN(n2949) );
  INVD1 U2933 ( .I(n189), .ZN(n2948) );
  INVD1 U2934 ( .I(n197), .ZN(n2947) );
  INVD1 U2935 ( .I(n197), .ZN(n2946) );
  INVD1 U2936 ( .I(n2945), .ZN(n2944) );
  BUFFD1 U2937 ( .I(n3048), .Z(n3052) );
  BUFFD1 U2938 ( .I(n2980), .Z(n3051) );
  BUFFD1 U2939 ( .I(n2980), .Z(n3050) );
  BUFFD1 U2940 ( .I(n2979), .Z(n3049) );
  BUFFD1 U2941 ( .I(n2978), .Z(n3048) );
  BUFFD1 U2942 ( .I(n2977), .Z(n3047) );
  BUFFD1 U2943 ( .I(n2977), .Z(n3046) );
  BUFFD1 U2944 ( .I(N44), .Z(n2909) );
  BUFFD1 U2945 ( .I(N44), .Z(n2910) );
  BUFFD1 U2946 ( .I(N44), .Z(n2911) );
  BUFFD1 U2947 ( .I(n2908), .Z(n2912) );
  BUFFD1 U2948 ( .I(n2908), .Z(n2913) );
  BUFFD1 U2949 ( .I(N45), .Z(n2903) );
  BUFFD1 U2950 ( .I(n3060), .Z(n2904) );
  BUFFD1 U2951 ( .I(N45), .Z(n2905) );
  BUFFD1 U2952 ( .I(n2902), .Z(n2906) );
  BUFFD1 U2953 ( .I(n2902), .Z(n2907) );
  INVD1 U2954 ( .I(N628), .ZN(n2945) );
  INVD1 U2955 ( .I(n193), .ZN(n2958) );
  INVD1 U2956 ( .I(n3058), .ZN(n3056) );
  INVD1 U2957 ( .I(n3058), .ZN(n3055) );
  INVD1 U2958 ( .I(n3058), .ZN(n3057) );
  BUFFD1 U2959 ( .I(ClockW), .Z(n2980) );
  BUFFD1 U2960 ( .I(n3046), .Z(n2979) );
  BUFFD1 U2961 ( .I(n2981), .Z(n2978) );
  BUFFD1 U2962 ( .I(n2981), .Z(n2977) );
  INVD1 U2963 ( .I(n3054), .ZN(n3053) );
  XOR3D1 U2964 ( .A1(n3148), .A2(n425), .A3(n3147), .Z(n3149) );
  XOR3D1 U2965 ( .A1(n2628), .A2(n2624), .A3(n3134), .Z(n3136) );
  XOR3D1 U2966 ( .A1(n3131), .A2(N57), .A3(n3130), .Z(n3132) );
  XOR3D1 U2967 ( .A1(n2684), .A2(n2681), .A3(n3137), .Z(n3138) );
  INVD1 U2968 ( .I(n2900), .ZN(n2901) );
  BUFFD1 U2969 ( .I(n3059), .Z(n2908) );
  BUFFD1 U2970 ( .I(n3060), .Z(n2902) );
  ND2D1 U2971 ( .A1(n3117), .A2(n3122), .ZN(n3120) );
  ND2D1 U2972 ( .A1(n3119), .A2(n3118), .ZN(n3124) );
  ND2D1 U2973 ( .A1(n3123), .A2(n3122), .ZN(n3127) );
  INVD1 U2974 ( .I(N364), .ZN(n2961) );
  INVD1 U2975 ( .I(n196), .ZN(n2973) );
  INVD1 U2976 ( .I(n2714), .ZN(n3058) );
  INVD1 U2977 ( .I(ClockR), .ZN(n3054) );
  BUFFD1 U2978 ( .I(ClockW), .Z(n2981) );
  MUX4D0 U2979 ( .I0(n2775), .I1(n2773), .I2(n2774), .I3(n2772), .S0(N47), 
        .S1(N46), .Z(N80) );
  MUX4D0 U2980 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(N44), .S1(N45), .Z(n2774)
         );
  MUX4D0 U2981 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n2912), .S1(n2902), .Z(
        n2773) );
  MUX4D0 U2982 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n3059), .S1(n2904), .Z(
        n2775) );
  MUX4D0 U2983 ( .I0(n2779), .I1(n2777), .I2(n2778), .I3(n2776), .S0(N47), 
        .S1(N46), .Z(N79) );
  MUX4D0 U2984 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(N44), .S1(N45), .Z(n2778)
         );
  MUX4D0 U2985 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(N44), .S1(n3060), .Z(
        n2777) );
  MUX4D0 U2986 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(N44), .S1(N45), .Z(n2779)
         );
  MUX4D0 U2987 ( .I0(n2799), .I1(n2797), .I2(n2798), .I3(n2796), .S0(N47), 
        .S1(N46), .Z(N74) );
  MUX4D0 U2988 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n2911), .S1(N45), .Z(n2798) );
  MUX4D0 U2989 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n2911), .S1(N45), .Z(
        n2797) );
  MUX4D0 U2990 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(N44), .S1(n2906), .Z(n2799) );
  MUX4D0 U2991 ( .I0(n2819), .I1(n2817), .I2(n2818), .I3(n2816), .S0(n2901), 
        .S1(n3061), .Z(N69) );
  MUX4D0 U2992 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n2908), .S1(n2907), .Z(
        n2818) );
  MUX4D0 U2993 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n2908), .S1(n2905), 
        .Z(n2817) );
  MUX4D0 U2994 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(N44), .S1(n2902), .Z(
        n2819) );
  MUX4D0 U2995 ( .I0(n2823), .I1(n2821), .I2(n2822), .I3(n2820), .S0(N47), 
        .S1(n3061), .Z(N68) );
  MUX4D0 U2996 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n2909), .S1(n2904), .Z(
        n2822) );
  MUX4D0 U2997 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n2910), .S1(n2904), 
        .Z(n2821) );
  MUX4D0 U2998 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n2912), .S1(n2907), .Z(
        n2823) );
  MUX4D0 U2999 ( .I0(n2847), .I1(n2845), .I2(n2846), .I3(n2844), .S0(N47), 
        .S1(n3061), .Z(N62) );
  MUX4D0 U3000 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n2909), .S1(n2903), .Z(
        n2846) );
  MUX4D0 U3001 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n2909), .S1(n2903), 
        .Z(n2845) );
  MUX4D0 U3002 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n2909), .S1(n2903), .Z(
        n2847) );
  MUX4D0 U3003 ( .I0(n2851), .I1(n2849), .I2(n2850), .I3(n2848), .S0(n2901), 
        .S1(N46), .Z(N61) );
  MUX4D0 U3004 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n2909), .S1(n2903), .Z(
        n2850) );
  MUX4D0 U3005 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n2909), .S1(n2903), 
        .Z(n2849) );
  MUX4D0 U3006 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n2909), .S1(n2903), .Z(
        n2851) );
  MUX4D0 U3007 ( .I0(n2875), .I1(n2873), .I2(n2874), .I3(n2872), .S0(n2901), 
        .S1(n3061), .Z(N55) );
  MUX4D0 U3008 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n2911), .S1(n2905), .Z(
        n2874) );
  MUX4D0 U3009 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n2911), .S1(n2905), 
        .Z(n2873) );
  MUX4D0 U3010 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n2911), .S1(n2905), .Z(
        n2875) );
  MUX4D0 U3011 ( .I0(n2879), .I1(n2877), .I2(n2878), .I3(n2876), .S0(n2901), 
        .S1(n3061), .Z(N54) );
  MUX4D0 U3012 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n2912), .S1(n2906), .Z(
        n2878) );
  MUX4D0 U3013 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n2912), .S1(n2906), 
        .Z(n2877) );
  MUX4D0 U3014 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n2912), .S1(n2906), .Z(
        n2879) );
  MUX4D0 U3015 ( .I0(n2891), .I1(n2889), .I2(n2890), .I3(n2888), .S0(n2901), 
        .S1(n3061), .Z(N51) );
  MUX4D0 U3016 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n2913), .S1(n2907), .Z(
        n2890) );
  MUX4D0 U3017 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n2913), .S1(n2907), 
        .Z(n2889) );
  MUX4D0 U3018 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n2913), .S1(n2907), .Z(
        n2891) );
  MUX4D0 U3019 ( .I0(n2895), .I1(n2893), .I2(n2894), .I3(n2892), .S0(n2901), 
        .S1(n3061), .Z(N50) );
  MUX4D0 U3020 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n2913), .S1(n2907), .Z(
        n2894) );
  MUX4D0 U3021 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n2913), .S1(n2907), 
        .Z(n2893) );
  MUX4D0 U3022 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n2913), .S1(n2907), .Z(
        n2895) );
  MUX4D0 U3023 ( .I0(n2795), .I1(n2793), .I2(n2794), .I3(n2792), .S0(N47), 
        .S1(N46), .Z(N75) );
  MUX4D0 U3024 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n2912), .S1(n2902), .Z(
        n2794) );
  MUX4D0 U3025 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n2913), .S1(n2906), .Z(
        n2793) );
  MUX4D0 U3026 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(N44), .S1(n2902), .Z(n2795) );
  MUX4D0 U3027 ( .I0(n2835), .I1(n2833), .I2(n2834), .I3(n2832), .S0(n2901), 
        .S1(n3061), .Z(N65) );
  MUX4D0 U3028 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(N44), .S1(n3060), .Z(
        n2834) );
  MUX4D0 U3029 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(N44), .S1(n2907), .Z(
        n2833) );
  MUX4D0 U3030 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n2913), .S1(n3060), .Z(
        n2835) );
  MUX4D0 U3031 ( .I0(n2863), .I1(n2861), .I2(n2862), .I3(n2860), .S0(n2901), 
        .S1(n3061), .Z(N58) );
  MUX4D0 U3032 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n2910), .S1(n2904), .Z(
        n2862) );
  MUX4D0 U3033 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n2910), .S1(n2904), 
        .Z(n2861) );
  MUX4D0 U3034 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n2910), .S1(n2904), .Z(
        n2863) );
  MUX4D0 U3035 ( .I0(n2867), .I1(n2865), .I2(n2866), .I3(n2864), .S0(n2901), 
        .S1(n3061), .Z(N57) );
  MUX4D0 U3036 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n2911), .S1(n2905), .Z(
        n2866) );
  MUX4D0 U3037 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n2911), .S1(n2905), 
        .Z(n2865) );
  MUX4D0 U3038 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n2911), .S1(n2905), .Z(
        n2867) );
  MUX4D0 U3039 ( .I0(n2771), .I1(n2769), .I2(n2770), .I3(n2768), .S0(n2901), 
        .S1(n3061), .Z(N81) );
  MUX4D0 U3040 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n2908), .S1(n2902), .Z(
        n2770) );
  MUX4D0 U3041 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n3059), .S1(n3060), .Z(
        n2769) );
  MUX4D0 U3042 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n3059), .S1(n3060), .Z(
        n2771) );
  MUX4D0 U3043 ( .I0(n2787), .I1(n2785), .I2(n2786), .I3(n2784), .S0(N47), 
        .S1(N46), .Z(N77) );
  MUX4D0 U3044 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n2908), .S1(n3060), .Z(
        n2786) );
  MUX4D0 U3045 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n3059), .S1(n2905), .Z(
        n2785) );
  MUX4D0 U3046 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n2913), .S1(n2905), .Z(
        n2787) );
  MUX4D0 U3047 ( .I0(n2811), .I1(n2809), .I2(n2810), .I3(n2808), .S0(N47), 
        .S1(N46), .Z(N71) );
  MUX4D0 U3048 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n2910), .S1(n2904), .Z(
        n2810) );
  MUX4D0 U3049 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n2909), .S1(n2903), 
        .Z(n2809) );
  MUX4D0 U3050 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n2910), .S1(n2904), .Z(
        n2811) );
  MUX4D0 U3051 ( .I0(n2815), .I1(n2813), .I2(n2814), .I3(n2812), .S0(N47), 
        .S1(N46), .Z(N70) );
  MUX4D0 U3052 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n2909), .S1(n2903), .Z(
        n2814) );
  MUX4D0 U3053 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n2910), .S1(n2903), 
        .Z(n2813) );
  MUX4D0 U3054 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n2909), .S1(n2903), .Z(
        n2815) );
  MUX4D0 U3055 ( .I0(n2827), .I1(n2825), .I2(n2826), .I3(n2824), .S0(N47), 
        .S1(N46), .Z(N67) );
  MUX4D0 U3056 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n2913), .S1(n2907), .Z(
        n2826) );
  MUX4D0 U3057 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n2913), .S1(n2903), 
        .Z(n2825) );
  MUX4D0 U3058 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n2910), .S1(n2907), .Z(
        n2827) );
  MUX4D0 U3059 ( .I0(n2843), .I1(n2841), .I2(n2842), .I3(n2840), .S0(N47), 
        .S1(n3061), .Z(N63) );
  MUX4D0 U3060 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n2909), .S1(n2903), .Z(
        n2842) );
  MUX4D0 U3061 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n2909), .S1(n2903), 
        .Z(n2841) );
  MUX4D0 U3062 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n2909), .S1(n2903), .Z(
        n2843) );
  MUX4D0 U3063 ( .I0(n2855), .I1(n2853), .I2(n2854), .I3(n2852), .S0(n2901), 
        .S1(n3061), .Z(N60) );
  MUX4D0 U3064 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n2910), .S1(n2904), .Z(
        n2854) );
  MUX4D0 U3065 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n2910), .S1(n2904), 
        .Z(n2853) );
  MUX4D0 U3066 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n2910), .S1(n2904), .Z(
        n2855) );
  MUX4D0 U3067 ( .I0(n2871), .I1(n2869), .I2(n2870), .I3(n2868), .S0(n2901), 
        .S1(n3061), .Z(N56) );
  MUX4D0 U3068 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n2911), .S1(n2905), .Z(
        n2870) );
  MUX4D0 U3069 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n2911), .S1(n2905), 
        .Z(n2869) );
  MUX4D0 U3070 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n2911), .S1(n2905), .Z(
        n2871) );
  MUX4D0 U3071 ( .I0(n2883), .I1(n2881), .I2(n2882), .I3(n2880), .S0(n2901), 
        .S1(n3061), .Z(N53) );
  MUX4D0 U3072 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n2912), .S1(n2906), .Z(
        n2882) );
  MUX4D0 U3073 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n2912), .S1(n2906), 
        .Z(n2881) );
  MUX4D0 U3074 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n2912), .S1(n2906), .Z(
        n2883) );
  MUX4D0 U3075 ( .I0(n2887), .I1(n2885), .I2(n2886), .I3(n2884), .S0(n2901), 
        .S1(n3061), .Z(N52) );
  MUX4D0 U3076 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n2912), .S1(n2906), .Z(
        n2886) );
  MUX4D0 U3077 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n2912), .S1(n2906), 
        .Z(n2885) );
  MUX4D0 U3078 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n2912), .S1(n2906), .Z(
        n2887) );
  MUX4D0 U3079 ( .I0(n2791), .I1(n2789), .I2(n2790), .I3(n2788), .S0(N47), 
        .S1(n3061), .Z(N76) );
  MUX4D0 U3080 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n2911), .S1(n2905), .Z(
        n2790) );
  MUX4D0 U3081 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n3059), .S1(n3060), .Z(
        n2789) );
  MUX4D0 U3082 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n2911), .S1(n2905), .Z(
        n2791) );
  MUX4D0 U3083 ( .I0(n2807), .I1(n2805), .I2(n2806), .I3(n2804), .S0(n2901), 
        .S1(n3061), .Z(N72) );
  MUX4D0 U3084 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(N44), .S1(N45), .Z(n2806)
         );
  MUX4D0 U3085 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n2909), .S1(n3060), .Z(
        n2805) );
  MUX4D0 U3086 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n2912), .S1(N45), .Z(n2807) );
  MUX4D0 U3087 ( .I0(n2831), .I1(n2829), .I2(n2830), .I3(n2828), .S0(N47), 
        .S1(N46), .Z(N66) );
  MUX4D0 U3088 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n3059), .S1(n3060), .Z(
        n2830) );
  MUX4D0 U3089 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n2908), .S1(n3060), 
        .Z(n2829) );
  MUX4D0 U3090 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(N44), .S1(n3060), .Z(
        n2831) );
  MUX4D0 U3091 ( .I0(n2839), .I1(n2837), .I2(n2838), .I3(n2836), .S0(N47), 
        .S1(N46), .Z(N64) );
  MUX4D0 U3092 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n2908), .S1(n3060), .Z(
        n2838) );
  MUX4D0 U3093 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n2909), .S1(n2904), 
        .Z(n2837) );
  MUX4D0 U3094 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n2908), .S1(n3060), .Z(
        n2839) );
  MUX4D0 U3095 ( .I0(n2859), .I1(n2857), .I2(n2858), .I3(n2856), .S0(n2901), 
        .S1(n3061), .Z(N59) );
  MUX4D0 U3096 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n2910), .S1(n2904), .Z(
        n2858) );
  MUX4D0 U3097 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n2910), .S1(n2904), 
        .Z(n2857) );
  MUX4D0 U3098 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n2910), .S1(n2904), .Z(
        n2859) );
  MUX4D0 U3099 ( .I0(n2899), .I1(n2897), .I2(n2898), .I3(n2896), .S0(n2901), 
        .S1(n3061), .Z(N49) );
  MUX4D0 U3100 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n2913), .S1(n2907), .Z(
        n2898) );
  MUX4D0 U3101 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n2913), .S1(n2907), 
        .Z(n2897) );
  MUX4D0 U3102 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n2913), .S1(n2907), .Z(
        n2899) );
  MUX4D0 U3103 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n2913), .S1(n2907), 
        .Z(n2896) );
  MUX4D0 U3104 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n3059), .S1(n2906), .Z(
        n2768) );
  MUX4D0 U3105 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(N44), .S1(N45), .Z(n2772) );
  MUX4D0 U3106 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(N44), .S1(N45), .Z(n2776) );
  MUX4D0 U3107 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n2908), .S1(n2907), .Z(
        n2784) );
  MUX4D0 U3108 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n3059), .S1(n2902), .Z(
        n2788) );
  MUX4D0 U3109 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n2908), .S1(n2904), .Z(
        n2792) );
  MUX4D0 U3110 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n2912), .S1(n3060), .Z(
        n2796) );
  MUX4D0 U3111 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n2908), .S1(N45), .Z(
        n2804) );
  MUX4D0 U3112 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n2909), .S1(n2903), 
        .Z(n2808) );
  MUX4D0 U3113 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n2910), .S1(n2903), 
        .Z(n2812) );
  MUX4D0 U3114 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n2908), .S1(n3060), 
        .Z(n2816) );
  MUX4D0 U3115 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n2913), .S1(n3060), 
        .Z(n2820) );
  MUX4D0 U3116 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n2913), .S1(n2903), 
        .Z(n2824) );
  MUX4D0 U3117 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n3059), .S1(n3060), 
        .Z(n2828) );
  MUX4D0 U3118 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n2908), .S1(N45), .Z(
        n2832) );
  MUX4D0 U3119 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n2908), .S1(n3060), 
        .Z(n2836) );
  MUX4D0 U3120 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n2909), .S1(n2903), 
        .Z(n2840) );
  MUX4D0 U3121 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n2909), .S1(n2903), 
        .Z(n2844) );
  MUX4D0 U3122 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n2909), .S1(n2903), 
        .Z(n2848) );
  MUX4D0 U3123 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n2910), .S1(n2904), 
        .Z(n2852) );
  MUX4D0 U3124 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n2910), .S1(n2904), 
        .Z(n2856) );
  MUX4D0 U3125 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n2910), .S1(n2904), 
        .Z(n2860) );
  MUX4D0 U3126 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n2911), .S1(n2905), 
        .Z(n2864) );
  MUX4D0 U3127 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n2911), .S1(n2905), 
        .Z(n2868) );
  MUX4D0 U3128 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n2911), .S1(n2905), 
        .Z(n2872) );
  MUX4D0 U3129 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n2912), .S1(n2906), 
        .Z(n2876) );
  MUX4D0 U3130 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n2912), .S1(n2906), 
        .Z(n2880) );
  MUX4D0 U3131 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n2912), .S1(n2906), 
        .Z(n2884) );
  MUX4D0 U3132 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n2913), .S1(n2907), 
        .Z(n2888) );
  MUX4D0 U3133 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n2913), .S1(n2907), 
        .Z(n2892) );
  BUFFD1 U3134 ( .I(N46), .Z(n3061) );
  BUFFD1 U3135 ( .I(N45), .Z(n3060) );
  MUX4D0 U3136 ( .I0(n2803), .I1(n2801), .I2(n2802), .I3(n2800), .S0(N47), 
        .S1(N46), .Z(N73) );
  MUX4D0 U3137 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n2911), .S1(n2904), .Z(
        n2802) );
  MUX4D0 U3138 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n2911), .S1(n2902), .Z(
        n2801) );
  MUX4D0 U3139 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n2908), .S1(n2905), .Z(
        n2803) );
  MUX4D0 U3140 ( .I0(n2783), .I1(n2781), .I2(n2782), .I3(n2780), .S0(N47), 
        .S1(N46), .Z(N78) );
  MUX4D0 U3141 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n2910), .S1(n2902), .Z(
        n2782) );
  MUX4D0 U3142 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n2908), .S1(n2902), .Z(
        n2781) );
  MUX4D0 U3143 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n2908), .S1(n2905), .Z(
        n2783) );
  MUX4D0 U3144 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n2911), .S1(n2905), .Z(
        n2780) );
  MUX4D0 U3145 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n2908), .S1(n2902), .Z(
        n2800) );
  ND2D1 U3146 ( .A1(AddrW[1]), .A2(n3118), .ZN(n3125) );
  ND2D1 U3147 ( .A1(AddrW[2]), .A2(AddrW[1]), .ZN(n3128) );
  ND2D1 U3148 ( .A1(n3117), .A2(AddrW[0]), .ZN(n3121) );
  ND2D1 U3149 ( .A1(AddrW[2]), .A2(n3119), .ZN(n3126) );
  ND2D1 U3150 ( .A1(AddrW[0]), .A2(n3123), .ZN(n3129) );
  INR2D1 U3151 ( .A1(Write), .B1(AddrW[3]), .ZN(n3117) );
  INVD1 U3152 ( .I(AddrW[1]), .ZN(n3119) );
  INVD1 U3153 ( .I(AddrW[0]), .ZN(n3122) );
  INVD1 U3154 ( .I(AddrW[2]), .ZN(n3118) );
  AN2D1 U3155 ( .A1(Write), .A2(AddrW[3]), .Z(n3123) );
  INR2D1 U3156 ( .A1(ClkW), .B1(N9), .ZN(ClockW) );
  INR2D1 U3157 ( .A1(ClkR), .B1(N9), .ZN(ClockR) );
  INVD0 U3158 ( .I(ChipEna), .ZN(N9) );
endmodule


module ClockComparator_1 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n1,
         n2, n3, n4, n6, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n89, n90, n91, n92, n93;

  AO211D1 U8 ( .A1(n92), .A2(n91), .B(N8), .C(N5), .Z(n90) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n93), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n93), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n89), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n89), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(n1), .CP(ClockIn), .CDN(n93), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(n13), .CP(ClockIn), .CDN(n93), .QN(n92) );
  DFSND1 ZeroCounters_reg ( .D(n23), .CP(ClockIn), .SDN(n89), .QN(n93) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(n6), .Z(n4) );
  BUFFD0 U7 ( .I(n10), .Z(n6) );
  BUFFD0 U9 ( .I(n11), .Z(n10) );
  BUFFD0 U10 ( .I(n12), .Z(n11) );
  BUFFD0 U11 ( .I(n85), .Z(n12) );
  BUFFD0 U12 ( .I(n14), .Z(n13) );
  BUFFD0 U13 ( .I(n15), .Z(n14) );
  BUFFD0 U14 ( .I(n16), .Z(n15) );
  BUFFD0 U15 ( .I(n17), .Z(n16) );
  BUFFD0 U16 ( .I(n18), .Z(n17) );
  BUFFD0 U17 ( .I(n19), .Z(n18) );
  BUFFD0 U18 ( .I(n20), .Z(n19) );
  BUFFD0 U19 ( .I(n82), .Z(n20) );
  BUFFD0 U20 ( .I(N5), .Z(n21) );
  BUFFD0 U21 ( .I(N6), .Z(n22) );
  BUFFD0 U22 ( .I(n28), .Z(n23) );
  BUFFD0 U23 ( .I(n21), .Z(n24) );
  BUFFD0 U24 ( .I(n22), .Z(n25) );
  BUFFD0 U25 ( .I(n24), .Z(n26) );
  BUFFD0 U26 ( .I(n25), .Z(n27) );
  BUFFD0 U27 ( .I(n31), .Z(n28) );
  BUFFD0 U28 ( .I(n26), .Z(n29) );
  BUFFD0 U29 ( .I(n27), .Z(n30) );
  BUFFD0 U30 ( .I(n34), .Z(n31) );
  BUFFD0 U31 ( .I(n29), .Z(n32) );
  BUFFD0 U32 ( .I(n30), .Z(n33) );
  BUFFD0 U33 ( .I(n37), .Z(n34) );
  BUFFD0 U34 ( .I(n32), .Z(n35) );
  BUFFD0 U35 ( .I(n33), .Z(n36) );
  BUFFD0 U36 ( .I(n40), .Z(n37) );
  BUFFD0 U37 ( .I(n35), .Z(n38) );
  BUFFD0 U38 ( .I(n36), .Z(n39) );
  BUFFD0 U39 ( .I(N9), .Z(n40) );
  BUFFD0 U40 ( .I(n38), .Z(n41) );
  BUFFD0 U41 ( .I(n39), .Z(n42) );
  BUFFD0 U42 ( .I(n41), .Z(n43) );
  BUFFD0 U43 ( .I(n42), .Z(n44) );
  BUFFD0 U44 ( .I(n43), .Z(n45) );
  BUFFD0 U45 ( .I(n44), .Z(n46) );
  BUFFD0 U46 ( .I(n45), .Z(n47) );
  BUFFD0 U47 ( .I(n46), .Z(n48) );
  BUFFD0 U48 ( .I(n47), .Z(n49) );
  BUFFD0 U49 ( .I(n48), .Z(n50) );
  BUFFD0 U50 ( .I(n49), .Z(n51) );
  BUFFD0 U51 ( .I(n50), .Z(n52) );
  BUFFD0 U52 ( .I(n51), .Z(n53) );
  BUFFD0 U53 ( .I(n52), .Z(n54) );
  BUFFD0 U54 ( .I(n53), .Z(n55) );
  BUFFD0 U55 ( .I(n54), .Z(n56) );
  BUFFD0 U56 ( .I(n55), .Z(n57) );
  BUFFD0 U57 ( .I(n56), .Z(n58) );
  BUFFD0 U58 ( .I(n57), .Z(n59) );
  BUFFD0 U59 ( .I(n58), .Z(n60) );
  BUFFD0 U60 ( .I(n59), .Z(n61) );
  BUFFD0 U61 ( .I(n60), .Z(n62) );
  BUFFD0 U62 ( .I(n61), .Z(n63) );
  BUFFD0 U63 ( .I(n62), .Z(n64) );
  BUFFD0 U64 ( .I(n63), .Z(n65) );
  BUFFD0 U65 ( .I(n64), .Z(n66) );
  BUFFD0 U66 ( .I(n65), .Z(n67) );
  BUFFD0 U67 ( .I(n66), .Z(n68) );
  BUFFD0 U68 ( .I(n67), .Z(n69) );
  BUFFD0 U69 ( .I(n68), .Z(n70) );
  BUFFD0 U70 ( .I(n69), .Z(n71) );
  BUFFD0 U71 ( .I(n70), .Z(n72) );
  BUFFD0 U72 ( .I(n71), .Z(n73) );
  BUFFD0 U73 ( .I(n72), .Z(n74) );
  BUFFD0 U74 ( .I(n73), .Z(n75) );
  BUFFD0 U75 ( .I(n74), .Z(n76) );
  BUFFD0 U76 ( .I(n75), .Z(n77) );
  BUFFD0 U77 ( .I(n76), .Z(n78) );
  BUFFD0 U78 ( .I(n77), .Z(n79) );
  BUFFD0 U79 ( .I(n78), .Z(n80) );
  BUFFD0 U80 ( .I(n79), .Z(n81) );
  CKBXD0 U81 ( .I(n80), .Z(n82) );
  BUFFD0 U82 ( .I(n81), .Z(n83) );
  BUFFD0 U83 ( .I(\ClockInN[0] ), .Z(n84) );
  XNR2D0 U84 ( .A1(n84), .A2(n92), .ZN(N6) );
  CKBD0 U85 ( .CLK(n83), .C(n85) );
  INVD1 U86 ( .I(Reset), .ZN(n89) );
  NR2D1 U87 ( .A1(n82), .A2(n85), .ZN(N9) );
  OAI21D1 U88 ( .A1(n91), .A2(n92), .B(n90), .ZN(N20) );
  NR2D1 U89 ( .A1(N19), .A2(N7), .ZN(n91) );
  XNR2D1 U90 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module ClockComparator_2 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n1,
         n2, n3, n4, n6, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n152, n153, n154, n155, n156;

  AO211D1 U8 ( .A1(n155), .A2(n154), .B(N8), .C(N5), .Z(n153) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n156), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n156), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n152), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n152), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(n1), .CP(ClockIn), .CDN(n156), .Q(
        \ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(n27), .CP(ClockIn), .CDN(n156), .QN(n155) );
  DFSND1 ZeroCounters_reg ( .D(n49), .CP(ClockIn), .SDN(n152), .QN(n156) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(n6), .Z(n4) );
  BUFFD0 U7 ( .I(n10), .Z(n6) );
  BUFFD0 U9 ( .I(n11), .Z(n10) );
  BUFFD0 U10 ( .I(n12), .Z(n11) );
  BUFFD0 U11 ( .I(n13), .Z(n12) );
  BUFFD0 U12 ( .I(n14), .Z(n13) );
  BUFFD0 U13 ( .I(n15), .Z(n14) );
  BUFFD0 U14 ( .I(n16), .Z(n15) );
  BUFFD0 U15 ( .I(n17), .Z(n16) );
  BUFFD0 U16 ( .I(n18), .Z(n17) );
  BUFFD0 U17 ( .I(n19), .Z(n18) );
  BUFFD0 U18 ( .I(n20), .Z(n19) );
  BUFFD0 U19 ( .I(n21), .Z(n20) );
  BUFFD0 U20 ( .I(n22), .Z(n21) );
  BUFFD0 U21 ( .I(n23), .Z(n22) );
  BUFFD0 U22 ( .I(n24), .Z(n23) );
  BUFFD0 U23 ( .I(n25), .Z(n24) );
  BUFFD0 U24 ( .I(n148), .Z(n25) );
  BUFFD0 U25 ( .I(N5), .Z(n26) );
  BUFFD0 U26 ( .I(n28), .Z(n27) );
  BUFFD0 U27 ( .I(n29), .Z(n28) );
  BUFFD0 U28 ( .I(n30), .Z(n29) );
  BUFFD0 U29 ( .I(n31), .Z(n30) );
  BUFFD0 U30 ( .I(n32), .Z(n31) );
  BUFFD0 U31 ( .I(n33), .Z(n32) );
  BUFFD0 U32 ( .I(n34), .Z(n33) );
  BUFFD0 U33 ( .I(n35), .Z(n34) );
  BUFFD0 U34 ( .I(n36), .Z(n35) );
  BUFFD0 U35 ( .I(n37), .Z(n36) );
  BUFFD0 U36 ( .I(n38), .Z(n37) );
  BUFFD0 U37 ( .I(n39), .Z(n38) );
  BUFFD0 U38 ( .I(n40), .Z(n39) );
  BUFFD0 U39 ( .I(n41), .Z(n40) );
  BUFFD0 U40 ( .I(n42), .Z(n41) );
  BUFFD0 U41 ( .I(n43), .Z(n42) );
  BUFFD0 U42 ( .I(n44), .Z(n43) );
  BUFFD0 U43 ( .I(n45), .Z(n44) );
  BUFFD0 U44 ( .I(n46), .Z(n45) );
  BUFFD0 U45 ( .I(n47), .Z(n46) );
  BUFFD0 U46 ( .I(n145), .Z(n47) );
  BUFFD0 U47 ( .I(N6), .Z(n48) );
  BUFFD0 U48 ( .I(n52), .Z(n49) );
  BUFFD0 U49 ( .I(n26), .Z(n50) );
  BUFFD0 U50 ( .I(n48), .Z(n51) );
  BUFFD0 U51 ( .I(n53), .Z(n52) );
  BUFFD0 U52 ( .I(n58), .Z(n53) );
  BUFFD0 U53 ( .I(n50), .Z(n54) );
  BUFFD0 U54 ( .I(n51), .Z(n55) );
  BUFFD0 U55 ( .I(n54), .Z(n56) );
  BUFFD0 U56 ( .I(n55), .Z(n57) );
  BUFFD0 U57 ( .I(n61), .Z(n58) );
  BUFFD0 U58 ( .I(n56), .Z(n59) );
  BUFFD0 U59 ( .I(n57), .Z(n60) );
  BUFFD0 U60 ( .I(n62), .Z(n61) );
  BUFFD0 U61 ( .I(n67), .Z(n62) );
  BUFFD0 U62 ( .I(n59), .Z(n63) );
  BUFFD0 U63 ( .I(n60), .Z(n64) );
  BUFFD0 U64 ( .I(n63), .Z(n65) );
  BUFFD0 U65 ( .I(n64), .Z(n66) );
  BUFFD0 U66 ( .I(n70), .Z(n67) );
  BUFFD0 U67 ( .I(n65), .Z(n68) );
  BUFFD0 U68 ( .I(n66), .Z(n69) );
  BUFFD0 U69 ( .I(n71), .Z(n70) );
  BUFFD0 U70 ( .I(n76), .Z(n71) );
  BUFFD0 U71 ( .I(n68), .Z(n72) );
  BUFFD0 U72 ( .I(n69), .Z(n73) );
  BUFFD0 U73 ( .I(n72), .Z(n74) );
  BUFFD0 U74 ( .I(n73), .Z(n75) );
  BUFFD0 U75 ( .I(n79), .Z(n76) );
  BUFFD0 U76 ( .I(n74), .Z(n77) );
  BUFFD0 U77 ( .I(n75), .Z(n78) );
  BUFFD0 U78 ( .I(n80), .Z(n79) );
  BUFFD0 U79 ( .I(n85), .Z(n80) );
  BUFFD0 U80 ( .I(n77), .Z(n81) );
  BUFFD0 U81 ( .I(n78), .Z(n82) );
  BUFFD0 U82 ( .I(n81), .Z(n83) );
  BUFFD0 U83 ( .I(n82), .Z(n84) );
  BUFFD0 U84 ( .I(n86), .Z(n85) );
  BUFFD0 U85 ( .I(n87), .Z(n86) );
  BUFFD0 U86 ( .I(n88), .Z(n87) );
  BUFFD0 U87 ( .I(n89), .Z(n88) );
  BUFFD0 U88 ( .I(n90), .Z(n89) );
  BUFFD0 U89 ( .I(n91), .Z(n90) );
  BUFFD0 U90 ( .I(N9), .Z(n91) );
  BUFFD0 U91 ( .I(n83), .Z(n92) );
  BUFFD0 U92 ( .I(n84), .Z(n93) );
  BUFFD0 U93 ( .I(n92), .Z(n94) );
  BUFFD0 U94 ( .I(n93), .Z(n95) );
  BUFFD0 U95 ( .I(n94), .Z(n96) );
  BUFFD0 U96 ( .I(n95), .Z(n97) );
  BUFFD0 U97 ( .I(n96), .Z(n98) );
  BUFFD0 U98 ( .I(n97), .Z(n99) );
  BUFFD0 U99 ( .I(n98), .Z(n100) );
  BUFFD0 U100 ( .I(n99), .Z(n101) );
  BUFFD0 U101 ( .I(n100), .Z(n102) );
  BUFFD0 U102 ( .I(n101), .Z(n103) );
  BUFFD0 U103 ( .I(n102), .Z(n104) );
  BUFFD0 U104 ( .I(n103), .Z(n105) );
  BUFFD0 U105 ( .I(n104), .Z(n106) );
  BUFFD0 U106 ( .I(n105), .Z(n107) );
  BUFFD0 U107 ( .I(n106), .Z(n108) );
  BUFFD0 U108 ( .I(n107), .Z(n109) );
  BUFFD0 U109 ( .I(n108), .Z(n110) );
  BUFFD0 U110 ( .I(n109), .Z(n111) );
  BUFFD0 U111 ( .I(n110), .Z(n112) );
  BUFFD0 U112 ( .I(n111), .Z(n113) );
  BUFFD0 U113 ( .I(n112), .Z(n114) );
  BUFFD0 U114 ( .I(n113), .Z(n115) );
  BUFFD0 U115 ( .I(n114), .Z(n116) );
  BUFFD0 U116 ( .I(n115), .Z(n117) );
  BUFFD0 U117 ( .I(n116), .Z(n118) );
  BUFFD0 U118 ( .I(n117), .Z(n119) );
  BUFFD0 U119 ( .I(n118), .Z(n120) );
  BUFFD0 U120 ( .I(n119), .Z(n121) );
  BUFFD0 U121 ( .I(n120), .Z(n122) );
  BUFFD0 U122 ( .I(n121), .Z(n123) );
  BUFFD0 U123 ( .I(n122), .Z(n124) );
  BUFFD0 U124 ( .I(n123), .Z(n125) );
  BUFFD0 U125 ( .I(n124), .Z(n126) );
  BUFFD0 U126 ( .I(n125), .Z(n127) );
  BUFFD0 U127 ( .I(n126), .Z(n128) );
  BUFFD0 U128 ( .I(n127), .Z(n129) );
  BUFFD0 U129 ( .I(n128), .Z(n130) );
  BUFFD0 U130 ( .I(n129), .Z(n131) );
  BUFFD0 U131 ( .I(n130), .Z(n132) );
  BUFFD0 U132 ( .I(n131), .Z(n133) );
  BUFFD0 U133 ( .I(n132), .Z(n134) );
  BUFFD0 U134 ( .I(n133), .Z(n135) );
  BUFFD0 U135 ( .I(n134), .Z(n136) );
  BUFFD0 U136 ( .I(n135), .Z(n137) );
  BUFFD0 U137 ( .I(n136), .Z(n138) );
  BUFFD0 U138 ( .I(n137), .Z(n139) );
  BUFFD0 U139 ( .I(n138), .Z(n140) );
  BUFFD0 U140 ( .I(n139), .Z(n141) );
  BUFFD0 U141 ( .I(n140), .Z(n142) );
  BUFFD0 U142 ( .I(n141), .Z(n143) );
  BUFFD0 U143 ( .I(n142), .Z(n144) );
  CKBD0 U144 ( .CLK(n143), .C(n145) );
  BUFFD0 U145 ( .I(n144), .Z(n146) );
  BUFFD0 U146 ( .I(\ClockInN[0] ), .Z(n147) );
  XNR2D0 U147 ( .A1(n147), .A2(n155), .ZN(N6) );
  CKBD0 U148 ( .CLK(n146), .C(n148) );
  INVD1 U149 ( .I(Reset), .ZN(n152) );
  NR2D1 U150 ( .A1(n145), .A2(n148), .ZN(N9) );
  OAI21D1 U151 ( .A1(n154), .A2(n155), .B(n153), .ZN(N20) );
  NR2D1 U152 ( .A1(N19), .A2(N7), .ZN(n154) );
  XNR2D1 U153 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module ClockComparator_3 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n1,
         n2, n3, n4, n6, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n89, n90, n91, n92, n93;

  AO211D1 U8 ( .A1(n92), .A2(n91), .B(N8), .C(N5), .Z(n90) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n93), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n93), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n89), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n89), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(n1), .CP(ClockIn), .CDN(n93), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(n13), .CP(ClockIn), .CDN(n93), .QN(n92) );
  DFSND1 ZeroCounters_reg ( .D(n25), .CP(ClockIn), .SDN(n89), .QN(n93) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(n6), .Z(n4) );
  BUFFD0 U7 ( .I(n10), .Z(n6) );
  BUFFD0 U9 ( .I(n11), .Z(n10) );
  BUFFD0 U10 ( .I(n12), .Z(n11) );
  BUFFD0 U11 ( .I(n85), .Z(n12) );
  BUFFD0 U12 ( .I(n14), .Z(n13) );
  BUFFD0 U13 ( .I(n15), .Z(n14) );
  BUFFD0 U14 ( .I(n16), .Z(n15) );
  BUFFD0 U15 ( .I(n17), .Z(n16) );
  BUFFD0 U16 ( .I(n18), .Z(n17) );
  BUFFD0 U17 ( .I(n19), .Z(n18) );
  BUFFD0 U18 ( .I(n20), .Z(n19) );
  BUFFD0 U19 ( .I(n82), .Z(n20) );
  BUFFD0 U20 ( .I(N5), .Z(n21) );
  BUFFD0 U21 ( .I(N6), .Z(n22) );
  BUFFD0 U22 ( .I(n21), .Z(n23) );
  BUFFD0 U23 ( .I(n22), .Z(n24) );
  BUFFD0 U24 ( .I(n28), .Z(n25) );
  BUFFD0 U25 ( .I(n23), .Z(n26) );
  BUFFD0 U26 ( .I(n24), .Z(n27) );
  BUFFD0 U27 ( .I(n31), .Z(n28) );
  BUFFD0 U28 ( .I(n26), .Z(n29) );
  BUFFD0 U29 ( .I(n27), .Z(n30) );
  BUFFD0 U30 ( .I(n32), .Z(n31) );
  BUFFD0 U31 ( .I(n33), .Z(n32) );
  BUFFD0 U32 ( .I(n34), .Z(n33) );
  BUFFD0 U33 ( .I(N9), .Z(n34) );
  BUFFD0 U34 ( .I(n29), .Z(n35) );
  BUFFD0 U35 ( .I(n30), .Z(n36) );
  BUFFD0 U36 ( .I(n35), .Z(n37) );
  BUFFD0 U37 ( .I(n36), .Z(n38) );
  BUFFD0 U38 ( .I(n37), .Z(n39) );
  BUFFD0 U39 ( .I(n38), .Z(n40) );
  BUFFD0 U40 ( .I(n39), .Z(n41) );
  BUFFD0 U41 ( .I(n40), .Z(n42) );
  BUFFD0 U42 ( .I(n41), .Z(n43) );
  BUFFD0 U43 ( .I(n42), .Z(n44) );
  BUFFD0 U44 ( .I(n43), .Z(n45) );
  BUFFD0 U45 ( .I(n44), .Z(n46) );
  BUFFD0 U46 ( .I(n45), .Z(n47) );
  BUFFD0 U47 ( .I(n46), .Z(n48) );
  BUFFD0 U48 ( .I(n47), .Z(n49) );
  BUFFD0 U49 ( .I(n48), .Z(n50) );
  BUFFD0 U50 ( .I(n49), .Z(n51) );
  BUFFD0 U51 ( .I(n50), .Z(n52) );
  BUFFD0 U52 ( .I(n51), .Z(n53) );
  BUFFD0 U53 ( .I(n52), .Z(n54) );
  BUFFD0 U54 ( .I(n53), .Z(n55) );
  BUFFD0 U55 ( .I(n54), .Z(n56) );
  BUFFD0 U56 ( .I(n55), .Z(n57) );
  BUFFD0 U57 ( .I(n56), .Z(n58) );
  BUFFD0 U58 ( .I(n57), .Z(n59) );
  BUFFD0 U59 ( .I(n58), .Z(n60) );
  BUFFD0 U60 ( .I(n59), .Z(n61) );
  BUFFD0 U61 ( .I(n60), .Z(n62) );
  BUFFD0 U62 ( .I(n61), .Z(n63) );
  BUFFD0 U63 ( .I(n62), .Z(n64) );
  BUFFD0 U64 ( .I(n63), .Z(n65) );
  BUFFD0 U65 ( .I(n64), .Z(n66) );
  BUFFD0 U66 ( .I(n65), .Z(n67) );
  BUFFD0 U67 ( .I(n66), .Z(n68) );
  BUFFD0 U68 ( .I(n67), .Z(n69) );
  BUFFD0 U69 ( .I(n68), .Z(n70) );
  BUFFD0 U70 ( .I(n69), .Z(n71) );
  BUFFD0 U71 ( .I(n70), .Z(n72) );
  BUFFD0 U72 ( .I(n71), .Z(n73) );
  BUFFD0 U73 ( .I(n72), .Z(n74) );
  BUFFD0 U74 ( .I(n73), .Z(n75) );
  BUFFD0 U75 ( .I(n74), .Z(n76) );
  BUFFD0 U76 ( .I(n75), .Z(n77) );
  BUFFD0 U77 ( .I(n76), .Z(n78) );
  BUFFD0 U78 ( .I(n77), .Z(n79) );
  BUFFD0 U79 ( .I(n78), .Z(n80) );
  BUFFD0 U80 ( .I(n79), .Z(n81) );
  CKBXD0 U81 ( .I(n80), .Z(n82) );
  BUFFD0 U82 ( .I(n81), .Z(n83) );
  BUFFD0 U83 ( .I(\ClockInN[0] ), .Z(n84) );
  XNR2D0 U84 ( .A1(n84), .A2(n92), .ZN(N6) );
  CKBD0 U85 ( .CLK(n83), .C(n85) );
  INVD1 U86 ( .I(Reset), .ZN(n89) );
  NR2D1 U87 ( .A1(n82), .A2(n85), .ZN(N9) );
  OAI21D1 U88 ( .A1(n91), .A2(n92), .B(n90), .ZN(N20) );
  NR2D1 U89 ( .A1(N19), .A2(N7), .ZN(n91) );
  XNR2D1 U90 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module VFO_1 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_1_DW01_dec_0 \Sampler/sub_193  ( .A({n210, n209, DivideFactor[3:2], n72, 
        n107}), .SUM({N40, N39, N38, N37, N36, N35}) );
  VFO_1_DW01_inc_0 \Sampler/add_190  ( .A({n210, n209, DivideFactor[3:2], n72, 
        n107}), .SUM({N32, N31, N30, N29, N28, N27}) );
  VFO_1_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n240), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n240), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n240), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n240), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n240), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n240), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n267), .CP(FastClock), .CDN(n240), .Q(ClockOut)
         );
  DFSND1 \DivideFactor_reg[4]  ( .D(n3), .CP(Sample), .SDN(n240), .Q(
        DivideFactor[4]), .QN(n251) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n40), .CP(Sample), .SDN(n240), .Q(
        DivideFactor[1]), .QN(n263) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n74), .CP(Sample), .SDN(n240), .Q(
        DivideFactor[0]), .QN(n261) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(n108), .E(n1), .CP(Sample), .CDN(n240), 
        .Q(DivideFactor[3]), .QN(n256) );
  EDFCND1 \DivideFactor_reg[2]  ( .D(n142), .E(n1), .CP(Sample), .CDN(n240), 
        .Q(DivideFactor[2]) );
  EDFCND1 \DivideFactor_reg[5]  ( .D(n176), .E(n1), .CP(Sample), .CDN(n240), 
        .Q(DivideFactor[5]), .QN(n246) );
  BUFFD0 U3 ( .I(n237), .Z(n1) );
  MUX2D0 U4 ( .I0(n238), .I1(n250), .S(AdjustFreq[0]), .Z(n2) );
  BUFFD0 U5 ( .I(n5), .Z(n3) );
  BUFFD0 U6 ( .I(n265), .Z(n4) );
  BUFFD0 U7 ( .I(n6), .Z(n5) );
  BUFFD0 U8 ( .I(n7), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(n10), .Z(n9) );
  BUFFD0 U12 ( .I(n11), .Z(n10) );
  BUFFD0 U13 ( .I(n12), .Z(n11) );
  BUFFD0 U14 ( .I(n13), .Z(n12) );
  BUFFD0 U15 ( .I(n14), .Z(n13) );
  BUFFD0 U16 ( .I(n15), .Z(n14) );
  CKBXD0 U17 ( .I(DivideFactor[4]), .Z(n209) );
  BUFFD0 U18 ( .I(n16), .Z(n15) );
  BUFFD0 U19 ( .I(n20), .Z(n16) );
  BUFFD0 U20 ( .I(n22), .Z(n20) );
  BUFFD0 U21 ( .I(n23), .Z(n22) );
  BUFFD0 U22 ( .I(n24), .Z(n23) );
  BUFFD0 U23 ( .I(n25), .Z(n24) );
  BUFFD0 U24 ( .I(n26), .Z(n25) );
  BUFFD0 U25 ( .I(n27), .Z(n26) );
  BUFFD0 U26 ( .I(n28), .Z(n27) );
  BUFFD0 U27 ( .I(n29), .Z(n28) );
  BUFFD0 U28 ( .I(n30), .Z(n29) );
  BUFFD0 U29 ( .I(n31), .Z(n30) );
  BUFFD0 U30 ( .I(n32), .Z(n31) );
  BUFFD0 U31 ( .I(n33), .Z(n32) );
  BUFFD0 U32 ( .I(n34), .Z(n33) );
  BUFFD0 U33 ( .I(n35), .Z(n34) );
  BUFFD0 U34 ( .I(n36), .Z(n35) );
  BUFFD0 U35 ( .I(n37), .Z(n36) );
  BUFFD0 U36 ( .I(n38), .Z(n37) );
  BUFFD0 U37 ( .I(n39), .Z(n38) );
  BUFFD0 U38 ( .I(n4), .Z(n39) );
  BUFFD0 U39 ( .I(n42), .Z(n40) );
  BUFFD0 U40 ( .I(n266), .Z(n41) );
  BUFFD0 U41 ( .I(n43), .Z(n42) );
  BUFFD0 U42 ( .I(n44), .Z(n43) );
  BUFFD0 U43 ( .I(n45), .Z(n44) );
  BUFFD0 U44 ( .I(n46), .Z(n45) );
  BUFFD0 U45 ( .I(n47), .Z(n46) );
  BUFFD0 U46 ( .I(n48), .Z(n47) );
  BUFFD0 U47 ( .I(n49), .Z(n48) );
  BUFFD0 U48 ( .I(n50), .Z(n49) );
  BUFFD0 U49 ( .I(n51), .Z(n50) );
  BUFFD0 U50 ( .I(n52), .Z(n51) );
  BUFFD0 U51 ( .I(n53), .Z(n52) );
  BUFFD0 U52 ( .I(n54), .Z(n53) );
  BUFFD0 U53 ( .I(n55), .Z(n54) );
  BUFFD0 U54 ( .I(n56), .Z(n55) );
  BUFFD0 U55 ( .I(n57), .Z(n56) );
  BUFFD0 U56 ( .I(n58), .Z(n57) );
  BUFFD0 U57 ( .I(n59), .Z(n58) );
  BUFFD0 U58 ( .I(n60), .Z(n59) );
  BUFFD0 U59 ( .I(n61), .Z(n60) );
  BUFFD0 U60 ( .I(n62), .Z(n61) );
  BUFFD0 U61 ( .I(n63), .Z(n62) );
  BUFFD0 U62 ( .I(n64), .Z(n63) );
  BUFFD0 U63 ( .I(n65), .Z(n64) );
  BUFFD0 U64 ( .I(n66), .Z(n65) );
  BUFFD0 U65 ( .I(n67), .Z(n66) );
  BUFFD0 U66 ( .I(n68), .Z(n67) );
  BUFFD0 U67 ( .I(n69), .Z(n68) );
  BUFFD0 U68 ( .I(n70), .Z(n69) );
  BUFFD0 U69 ( .I(n71), .Z(n70) );
  BUFFD0 U70 ( .I(n41), .Z(n71) );
  BUFFD0 U71 ( .I(n73), .Z(n72) );
  BUFFD0 U72 ( .I(DivideFactor[1]), .Z(n73) );
  BUFFD0 U73 ( .I(n76), .Z(n74) );
  BUFFD0 U74 ( .I(n264), .Z(n75) );
  BUFFD0 U75 ( .I(n77), .Z(n76) );
  BUFFD0 U76 ( .I(n78), .Z(n77) );
  BUFFD0 U77 ( .I(n79), .Z(n78) );
  BUFFD0 U78 ( .I(n80), .Z(n79) );
  BUFFD0 U79 ( .I(n81), .Z(n80) );
  BUFFD0 U80 ( .I(n82), .Z(n81) );
  BUFFD0 U81 ( .I(n83), .Z(n82) );
  BUFFD0 U82 ( .I(n84), .Z(n83) );
  BUFFD0 U83 ( .I(n85), .Z(n84) );
  BUFFD0 U84 ( .I(n86), .Z(n85) );
  BUFFD0 U85 ( .I(n87), .Z(n86) );
  BUFFD0 U86 ( .I(n88), .Z(n87) );
  BUFFD0 U87 ( .I(n89), .Z(n88) );
  BUFFD0 U88 ( .I(n90), .Z(n89) );
  BUFFD0 U89 ( .I(n91), .Z(n90) );
  BUFFD0 U90 ( .I(n92), .Z(n91) );
  BUFFD0 U91 ( .I(n93), .Z(n92) );
  BUFFD0 U92 ( .I(n94), .Z(n93) );
  BUFFD0 U93 ( .I(n95), .Z(n94) );
  BUFFD0 U94 ( .I(n96), .Z(n95) );
  BUFFD0 U95 ( .I(n97), .Z(n96) );
  BUFFD0 U96 ( .I(n98), .Z(n97) );
  BUFFD0 U97 ( .I(n99), .Z(n98) );
  BUFFD0 U98 ( .I(n100), .Z(n99) );
  BUFFD0 U99 ( .I(n101), .Z(n100) );
  BUFFD0 U100 ( .I(n102), .Z(n101) );
  BUFFD0 U101 ( .I(n103), .Z(n102) );
  BUFFD0 U102 ( .I(n104), .Z(n103) );
  BUFFD0 U103 ( .I(n105), .Z(n104) );
  BUFFD0 U104 ( .I(n75), .Z(n105) );
  BUFFD0 U105 ( .I(DivideFactor[0]), .Z(n106) );
  CKBXD0 U106 ( .I(n106), .Z(n107) );
  BUFFD0 U107 ( .I(n110), .Z(n108) );
  BUFFD0 U108 ( .I(N51), .Z(n109) );
  BUFFD0 U109 ( .I(n111), .Z(n110) );
  BUFFD0 U110 ( .I(n112), .Z(n111) );
  BUFFD0 U111 ( .I(n113), .Z(n112) );
  BUFFD0 U112 ( .I(n114), .Z(n113) );
  BUFFD0 U113 ( .I(n115), .Z(n114) );
  BUFFD0 U114 ( .I(n116), .Z(n115) );
  BUFFD0 U115 ( .I(n117), .Z(n116) );
  BUFFD0 U116 ( .I(n118), .Z(n117) );
  BUFFD0 U117 ( .I(n119), .Z(n118) );
  BUFFD0 U118 ( .I(n120), .Z(n119) );
  BUFFD0 U119 ( .I(n121), .Z(n120) );
  BUFFD0 U120 ( .I(n122), .Z(n121) );
  BUFFD0 U121 ( .I(n123), .Z(n122) );
  BUFFD0 U122 ( .I(n124), .Z(n123) );
  BUFFD0 U123 ( .I(n125), .Z(n124) );
  BUFFD0 U124 ( .I(n126), .Z(n125) );
  BUFFD0 U125 ( .I(n127), .Z(n126) );
  BUFFD0 U126 ( .I(n128), .Z(n127) );
  BUFFD0 U127 ( .I(n129), .Z(n128) );
  BUFFD0 U128 ( .I(n130), .Z(n129) );
  BUFFD0 U129 ( .I(n131), .Z(n130) );
  BUFFD0 U130 ( .I(n132), .Z(n131) );
  BUFFD0 U131 ( .I(n133), .Z(n132) );
  BUFFD0 U132 ( .I(n134), .Z(n133) );
  BUFFD0 U133 ( .I(n135), .Z(n134) );
  BUFFD0 U134 ( .I(n136), .Z(n135) );
  BUFFD0 U135 ( .I(n137), .Z(n136) );
  BUFFD0 U136 ( .I(n138), .Z(n137) );
  BUFFD0 U137 ( .I(n139), .Z(n138) );
  BUFFD0 U138 ( .I(n140), .Z(n139) );
  BUFFD0 U139 ( .I(n141), .Z(n140) );
  BUFFD0 U140 ( .I(n109), .Z(n141) );
  BUFFD0 U141 ( .I(n144), .Z(n142) );
  BUFFD0 U142 ( .I(N49), .Z(n143) );
  BUFFD0 U143 ( .I(n145), .Z(n144) );
  BUFFD0 U144 ( .I(n146), .Z(n145) );
  BUFFD0 U145 ( .I(n147), .Z(n146) );
  BUFFD0 U146 ( .I(n148), .Z(n147) );
  BUFFD0 U147 ( .I(n149), .Z(n148) );
  BUFFD0 U148 ( .I(n150), .Z(n149) );
  BUFFD0 U149 ( .I(n151), .Z(n150) );
  BUFFD0 U150 ( .I(n152), .Z(n151) );
  BUFFD0 U151 ( .I(n153), .Z(n152) );
  BUFFD0 U152 ( .I(n154), .Z(n153) );
  BUFFD0 U153 ( .I(n155), .Z(n154) );
  BUFFD0 U154 ( .I(n156), .Z(n155) );
  BUFFD0 U155 ( .I(n157), .Z(n156) );
  BUFFD0 U156 ( .I(n158), .Z(n157) );
  BUFFD0 U157 ( .I(n159), .Z(n158) );
  BUFFD0 U158 ( .I(n160), .Z(n159) );
  BUFFD0 U159 ( .I(n161), .Z(n160) );
  BUFFD0 U160 ( .I(n162), .Z(n161) );
  BUFFD0 U161 ( .I(n163), .Z(n162) );
  BUFFD0 U162 ( .I(n164), .Z(n163) );
  BUFFD0 U163 ( .I(n165), .Z(n164) );
  BUFFD0 U164 ( .I(n166), .Z(n165) );
  BUFFD0 U165 ( .I(n167), .Z(n166) );
  BUFFD0 U166 ( .I(n168), .Z(n167) );
  BUFFD0 U167 ( .I(n169), .Z(n168) );
  BUFFD0 U168 ( .I(n170), .Z(n169) );
  BUFFD0 U169 ( .I(n171), .Z(n170) );
  BUFFD0 U170 ( .I(n172), .Z(n171) );
  BUFFD0 U171 ( .I(n173), .Z(n172) );
  BUFFD0 U172 ( .I(n174), .Z(n173) );
  BUFFD0 U173 ( .I(n175), .Z(n174) );
  BUFFD0 U174 ( .I(n143), .Z(n175) );
  BUFFD0 U175 ( .I(n178), .Z(n176) );
  BUFFD0 U176 ( .I(N55), .Z(n177) );
  BUFFD0 U177 ( .I(n179), .Z(n178) );
  BUFFD0 U178 ( .I(n180), .Z(n179) );
  BUFFD0 U179 ( .I(n181), .Z(n180) );
  BUFFD0 U180 ( .I(n182), .Z(n181) );
  BUFFD0 U181 ( .I(n183), .Z(n182) );
  BUFFD0 U182 ( .I(n184), .Z(n183) );
  BUFFD0 U183 ( .I(n185), .Z(n184) );
  BUFFD0 U184 ( .I(n186), .Z(n185) );
  BUFFD0 U185 ( .I(n187), .Z(n186) );
  BUFFD0 U186 ( .I(n188), .Z(n187) );
  BUFFD0 U187 ( .I(n189), .Z(n188) );
  BUFFD0 U188 ( .I(n190), .Z(n189) );
  BUFFD0 U189 ( .I(n191), .Z(n190) );
  BUFFD0 U190 ( .I(n192), .Z(n191) );
  BUFFD0 U191 ( .I(n193), .Z(n192) );
  BUFFD0 U192 ( .I(n194), .Z(n193) );
  BUFFD0 U193 ( .I(n195), .Z(n194) );
  BUFFD0 U194 ( .I(n196), .Z(n195) );
  BUFFD0 U195 ( .I(n197), .Z(n196) );
  BUFFD0 U196 ( .I(n198), .Z(n197) );
  BUFFD0 U197 ( .I(n199), .Z(n198) );
  BUFFD0 U198 ( .I(n200), .Z(n199) );
  BUFFD0 U199 ( .I(n201), .Z(n200) );
  BUFFD0 U200 ( .I(n202), .Z(n201) );
  BUFFD0 U201 ( .I(n203), .Z(n202) );
  BUFFD0 U202 ( .I(n204), .Z(n203) );
  BUFFD0 U203 ( .I(n205), .Z(n204) );
  BUFFD0 U204 ( .I(n206), .Z(n205) );
  BUFFD0 U205 ( .I(n207), .Z(n206) );
  BUFFD0 U206 ( .I(n177), .Z(n207) );
  BUFFD0 U207 ( .I(DivideFactor[5]), .Z(n208) );
  CKBD0 U208 ( .CLK(n208), .C(n210) );
  CKNXD0 U209 ( .I(n2), .ZN(n211) );
  CKBD0 U210 ( .CLK(n211), .C(n212) );
  CKBD0 U211 ( .CLK(n212), .C(n213) );
  CKBD0 U212 ( .CLK(n213), .C(n214) );
  CKBD0 U213 ( .CLK(n214), .C(n215) );
  CKBD0 U214 ( .CLK(n215), .C(n216) );
  CKBD0 U215 ( .CLK(n216), .C(n217) );
  CKBD0 U216 ( .CLK(n217), .C(n218) );
  CKBD0 U217 ( .CLK(n218), .C(n219) );
  CKBD0 U218 ( .CLK(n219), .C(n220) );
  CKBD0 U219 ( .CLK(n220), .C(n221) );
  BUFFD0 U220 ( .I(n221), .Z(n222) );
  CKBD0 U221 ( .CLK(n222), .C(n223) );
  CKBD0 U222 ( .CLK(n223), .C(n224) );
  CKBD0 U223 ( .CLK(n224), .C(n225) );
  CKBD0 U224 ( .CLK(n225), .C(n226) );
  CKBD0 U225 ( .CLK(n226), .C(n227) );
  CKBD0 U226 ( .CLK(n227), .C(n228) );
  CKBD0 U227 ( .CLK(n228), .C(n229) );
  CKBD0 U228 ( .CLK(n229), .C(n230) );
  CKBD0 U229 ( .CLK(n230), .C(n231) );
  BUFFD0 U230 ( .I(n231), .Z(n232) );
  CKBD0 U231 ( .CLK(n232), .C(n233) );
  BUFFD0 U232 ( .I(n233), .Z(n234) );
  CKBD0 U233 ( .CLK(n234), .C(n235) );
  BUFFD0 U234 ( .I(n235), .Z(n236) );
  CKBXD0 U235 ( .I(n236), .Z(n237) );
  BUFFD0 U236 ( .I(n249), .Z(n238) );
  INVD1 U237 ( .I(Reset), .ZN(n240) );
  AO222D0 U238 ( .A1(N27), .A2(n241), .B1(N35), .B2(n242), .C1(n107), .C2(n2), 
        .Z(n264) );
  AO222D0 U239 ( .A1(N31), .A2(n241), .B1(N39), .B2(n242), .C1(n209), .C2(n2), 
        .Z(n265) );
  AO222D0 U240 ( .A1(N28), .A2(n241), .B1(N36), .B2(n242), .C1(n72), .C2(n2), 
        .Z(n266) );
  AN2D0 U241 ( .A1(n243), .A2(n244), .Z(n242) );
  AN3D0 U242 ( .A1(n245), .A2(n246), .A3(n247), .Z(n241) );
  CKXOR2D0 U243 ( .A1(ClockOut), .A2(n248), .Z(n267) );
  AO22D0 U244 ( .A1(N32), .A2(n247), .B1(N40), .B2(n243), .Z(N55) );
  CKND2D0 U245 ( .A1(AdjustFreq[1]), .A2(n244), .ZN(n250) );
  ND3D0 U246 ( .A1(n251), .A2(n246), .A3(n252), .ZN(n244) );
  ND4D0 U247 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(n72), .A4(n107), 
        .ZN(n252) );
  IND3D0 U248 ( .A1(AdjustFreq[1]), .B1(n246), .B2(n245), .ZN(n249) );
  CKND2D0 U249 ( .A1(n209), .A2(DivideFactor[3]), .ZN(n245) );
  AO22D0 U250 ( .A1(N30), .A2(n247), .B1(N38), .B2(n243), .Z(N51) );
  AO22D0 U251 ( .A1(N29), .A2(n247), .B1(N37), .B2(n243), .Z(N49) );
  AN2D0 U252 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n243) );
  NR2D0 U253 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n247) );
  INR2D0 U254 ( .A1(N14), .B1(n248), .ZN(N21) );
  INR2D0 U255 ( .A1(N13), .B1(n248), .ZN(N20) );
  INR2D0 U256 ( .A1(N12), .B1(n248), .ZN(N19) );
  INR2D0 U257 ( .A1(N11), .B1(n248), .ZN(N18) );
  INR2D0 U258 ( .A1(N10), .B1(n248), .ZN(N17) );
  INR2D0 U259 ( .A1(N9), .B1(n248), .ZN(N16) );
  OA21D0 U260 ( .A1(FastDivvy[5]), .A2(n246), .B(n253), .Z(n248) );
  IOA22D0 U261 ( .B1(n254), .B2(n255), .A1(n246), .A2(FastDivvy[5]), .ZN(n253)
         );
  AOI221D0 U262 ( .A1(FastDivvy[4]), .A2(n251), .B1(FastDivvy[3]), .B2(n256), 
        .C(n257), .ZN(n255) );
  AOI221D0 U263 ( .A1(DivideFactor[3]), .A2(n258), .B1(DivideFactor[2]), .B2(
        n259), .C(n260), .ZN(n257) );
  IAO21D0 U264 ( .A1(n259), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n260)
         );
  OAI32D0 U265 ( .A1(n261), .A2(FastDivvy[0]), .A3(n262), .B1(FastDivvy[1]), 
        .B2(n263), .ZN(n259) );
  AN2D0 U266 ( .A1(FastDivvy[1]), .A2(n263), .Z(n262) );
  CKND0 U267 ( .CLK(FastDivvy[3]), .CN(n258) );
  NR2D0 U268 ( .A1(FastDivvy[4]), .A2(n251), .ZN(n254) );
  CKND0 U269 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U270 ( .A1(WireD[5]), .A2(n240), .ZN(WireD[0]) );
endmodule


module VFO_2 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_2_DW01_dec_0 \Sampler/sub_193  ( .A({n64, n182, DivideFactor[3], n123, 
        n240, n300}), .SUM({N40, N39, N38, N37, N36, N35}) );
  VFO_2_DW01_inc_0 \Sampler/add_190  ( .A({n64, n182, DivideFactor[3], n123, 
        n240, n300}), .SUM({N32, N31, N30, N29, N28, N27}) );
  VFO_2_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n416), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n444), .CP(FastClock), .CDN(n416), .Q(ClockOut)
         );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(n2), .E(n361), .CP(Sample), .CDN(n416), 
        .Q(DivideFactor[5]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(n65), .E(n361), .CP(Sample), .CDN(n416), 
        .Q(DivideFactor[2]) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n124), .CP(Sample), .SDN(n416), .Q(
        DivideFactor[4]), .QN(n428) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n183), .CP(Sample), .SDN(n416), .Q(
        DivideFactor[1]), .QN(n440) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n242), .CP(Sample), .SDN(n416), .Q(
        DivideFactor[0]), .QN(n438) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(n301), .E(n361), .CP(Sample), .CDN(n416), 
        .Q(DivideFactor[3]), .QN(n433) );
  INVD4 U3 ( .I(n1), .ZN(N54) );
  MUX2D0 U4 ( .I0(n415), .I1(n427), .S(AdjustFreq[0]), .Z(n1) );
  BUFFD0 U5 ( .I(n5), .Z(n2) );
  BUFFD0 U6 ( .I(N55), .Z(n3) );
  BUFFD0 U7 ( .I(n3), .Z(n4) );
  BUFFD0 U8 ( .I(n6), .Z(n5) );
  BUFFD0 U9 ( .I(n7), .Z(n6) );
  BUFFD0 U10 ( .I(n8), .Z(n7) );
  BUFFD0 U11 ( .I(n9), .Z(n8) );
  BUFFD0 U12 ( .I(n10), .Z(n9) );
  BUFFD0 U13 ( .I(n11), .Z(n10) );
  BUFFD0 U14 ( .I(n12), .Z(n11) );
  BUFFD0 U15 ( .I(n13), .Z(n12) );
  BUFFD0 U16 ( .I(n14), .Z(n13) );
  BUFFD0 U17 ( .I(n15), .Z(n14) );
  BUFFD0 U18 ( .I(n16), .Z(n15) );
  BUFFD0 U19 ( .I(n20), .Z(n16) );
  BUFFD0 U20 ( .I(n22), .Z(n20) );
  BUFFD0 U21 ( .I(n23), .Z(n22) );
  BUFFD0 U22 ( .I(n24), .Z(n23) );
  BUFFD0 U23 ( .I(n25), .Z(n24) );
  BUFFD0 U24 ( .I(n26), .Z(n25) );
  BUFFD0 U25 ( .I(n27), .Z(n26) );
  BUFFD0 U26 ( .I(n28), .Z(n27) );
  BUFFD0 U27 ( .I(n29), .Z(n28) );
  BUFFD0 U28 ( .I(n30), .Z(n29) );
  BUFFD0 U29 ( .I(n31), .Z(n30) );
  BUFFD0 U30 ( .I(n32), .Z(n31) );
  BUFFD0 U31 ( .I(n33), .Z(n32) );
  BUFFD0 U32 ( .I(n34), .Z(n33) );
  BUFFD0 U33 ( .I(n35), .Z(n34) );
  BUFFD0 U34 ( .I(n36), .Z(n35) );
  BUFFD0 U35 ( .I(n37), .Z(n36) );
  BUFFD0 U36 ( .I(n38), .Z(n37) );
  BUFFD0 U37 ( .I(n39), .Z(n38) );
  BUFFD0 U38 ( .I(n40), .Z(n39) );
  BUFFD0 U39 ( .I(n41), .Z(n40) );
  BUFFD0 U40 ( .I(n42), .Z(n41) );
  BUFFD0 U41 ( .I(n43), .Z(n42) );
  BUFFD0 U42 ( .I(n44), .Z(n43) );
  BUFFD0 U43 ( .I(n45), .Z(n44) );
  BUFFD0 U44 ( .I(n46), .Z(n45) );
  BUFFD0 U45 ( .I(n47), .Z(n46) );
  BUFFD0 U46 ( .I(n48), .Z(n47) );
  BUFFD0 U47 ( .I(n49), .Z(n48) );
  BUFFD0 U48 ( .I(n50), .Z(n49) );
  BUFFD0 U49 ( .I(n51), .Z(n50) );
  BUFFD0 U50 ( .I(n52), .Z(n51) );
  BUFFD0 U51 ( .I(n53), .Z(n52) );
  BUFFD0 U52 ( .I(n54), .Z(n53) );
  BUFFD0 U53 ( .I(n55), .Z(n54) );
  BUFFD0 U54 ( .I(n56), .Z(n55) );
  BUFFD0 U55 ( .I(n57), .Z(n56) );
  BUFFD0 U56 ( .I(n58), .Z(n57) );
  BUFFD0 U57 ( .I(n59), .Z(n58) );
  BUFFD0 U58 ( .I(n60), .Z(n59) );
  BUFFD0 U59 ( .I(n61), .Z(n60) );
  BUFFD0 U60 ( .I(n62), .Z(n61) );
  BUFFD0 U61 ( .I(n4), .Z(n62) );
  BUFFD0 U62 ( .I(DivideFactor[5]), .Z(n63) );
  CKBD0 U63 ( .CLK(n63), .C(n64) );
  BUFFD0 U64 ( .I(n69), .Z(n65) );
  BUFFD0 U65 ( .I(N49), .Z(n66) );
  BUFFD0 U66 ( .I(n66), .Z(n67) );
  BUFFD0 U67 ( .I(n67), .Z(n68) );
  BUFFD0 U68 ( .I(n70), .Z(n69) );
  BUFFD0 U69 ( .I(n71), .Z(n70) );
  BUFFD0 U70 ( .I(n72), .Z(n71) );
  BUFFD0 U71 ( .I(n73), .Z(n72) );
  BUFFD0 U72 ( .I(n74), .Z(n73) );
  BUFFD0 U73 ( .I(n75), .Z(n74) );
  BUFFD0 U74 ( .I(n76), .Z(n75) );
  BUFFD0 U75 ( .I(n77), .Z(n76) );
  BUFFD0 U76 ( .I(n78), .Z(n77) );
  BUFFD0 U77 ( .I(n79), .Z(n78) );
  BUFFD0 U78 ( .I(n80), .Z(n79) );
  BUFFD0 U79 ( .I(n81), .Z(n80) );
  BUFFD0 U80 ( .I(n82), .Z(n81) );
  BUFFD0 U81 ( .I(n83), .Z(n82) );
  BUFFD0 U82 ( .I(n84), .Z(n83) );
  BUFFD0 U83 ( .I(n85), .Z(n84) );
  BUFFD0 U84 ( .I(n86), .Z(n85) );
  BUFFD0 U85 ( .I(n87), .Z(n86) );
  BUFFD0 U86 ( .I(n88), .Z(n87) );
  BUFFD0 U87 ( .I(n89), .Z(n88) );
  BUFFD0 U88 ( .I(n90), .Z(n89) );
  BUFFD0 U89 ( .I(n91), .Z(n90) );
  BUFFD0 U90 ( .I(n92), .Z(n91) );
  BUFFD0 U91 ( .I(n93), .Z(n92) );
  BUFFD0 U92 ( .I(n94), .Z(n93) );
  BUFFD0 U93 ( .I(n95), .Z(n94) );
  BUFFD0 U94 ( .I(n96), .Z(n95) );
  BUFFD0 U95 ( .I(n97), .Z(n96) );
  BUFFD0 U96 ( .I(n98), .Z(n97) );
  BUFFD0 U97 ( .I(n99), .Z(n98) );
  BUFFD0 U98 ( .I(n100), .Z(n99) );
  BUFFD0 U99 ( .I(n101), .Z(n100) );
  BUFFD0 U100 ( .I(n102), .Z(n101) );
  BUFFD0 U101 ( .I(n103), .Z(n102) );
  BUFFD0 U102 ( .I(n104), .Z(n103) );
  BUFFD0 U103 ( .I(n105), .Z(n104) );
  BUFFD0 U104 ( .I(n106), .Z(n105) );
  BUFFD0 U105 ( .I(n107), .Z(n106) );
  BUFFD0 U106 ( .I(n108), .Z(n107) );
  BUFFD0 U107 ( .I(n109), .Z(n108) );
  BUFFD0 U108 ( .I(n110), .Z(n109) );
  BUFFD0 U109 ( .I(n111), .Z(n110) );
  BUFFD0 U110 ( .I(n112), .Z(n111) );
  BUFFD0 U111 ( .I(n113), .Z(n112) );
  BUFFD0 U112 ( .I(n114), .Z(n113) );
  BUFFD0 U113 ( .I(n115), .Z(n114) );
  BUFFD0 U114 ( .I(n116), .Z(n115) );
  BUFFD0 U115 ( .I(n117), .Z(n116) );
  BUFFD0 U116 ( .I(n118), .Z(n117) );
  BUFFD0 U117 ( .I(n119), .Z(n118) );
  BUFFD0 U118 ( .I(n120), .Z(n119) );
  BUFFD0 U119 ( .I(n121), .Z(n120) );
  BUFFD0 U120 ( .I(n68), .Z(n121) );
  BUFFD0 U121 ( .I(DivideFactor[2]), .Z(n122) );
  CKBD0 U122 ( .CLK(n122), .C(n123) );
  BUFFD0 U123 ( .I(n127), .Z(n124) );
  BUFFD0 U124 ( .I(n442), .Z(n125) );
  BUFFD0 U125 ( .I(n125), .Z(n126) );
  BUFFD0 U126 ( .I(n128), .Z(n127) );
  BUFFD0 U127 ( .I(n129), .Z(n128) );
  BUFFD0 U128 ( .I(n130), .Z(n129) );
  BUFFD0 U129 ( .I(n131), .Z(n130) );
  BUFFD0 U130 ( .I(n132), .Z(n131) );
  BUFFD0 U131 ( .I(n133), .Z(n132) );
  BUFFD0 U132 ( .I(n134), .Z(n133) );
  BUFFD0 U133 ( .I(n135), .Z(n134) );
  BUFFD0 U134 ( .I(n136), .Z(n135) );
  BUFFD0 U135 ( .I(n137), .Z(n136) );
  BUFFD0 U136 ( .I(n138), .Z(n137) );
  BUFFD0 U137 ( .I(n139), .Z(n138) );
  BUFFD0 U138 ( .I(n140), .Z(n139) );
  BUFFD0 U139 ( .I(n141), .Z(n140) );
  BUFFD0 U140 ( .I(n142), .Z(n141) );
  BUFFD0 U141 ( .I(n143), .Z(n142) );
  BUFFD0 U142 ( .I(n144), .Z(n143) );
  BUFFD0 U143 ( .I(n145), .Z(n144) );
  BUFFD0 U144 ( .I(n146), .Z(n145) );
  BUFFD0 U145 ( .I(n147), .Z(n146) );
  BUFFD0 U146 ( .I(n148), .Z(n147) );
  BUFFD0 U147 ( .I(n149), .Z(n148) );
  BUFFD0 U148 ( .I(n150), .Z(n149) );
  BUFFD0 U149 ( .I(n151), .Z(n150) );
  BUFFD0 U150 ( .I(n152), .Z(n151) );
  BUFFD0 U151 ( .I(n153), .Z(n152) );
  BUFFD0 U152 ( .I(n154), .Z(n153) );
  BUFFD0 U153 ( .I(n155), .Z(n154) );
  BUFFD0 U154 ( .I(n156), .Z(n155) );
  BUFFD0 U155 ( .I(n157), .Z(n156) );
  BUFFD0 U156 ( .I(n158), .Z(n157) );
  BUFFD0 U157 ( .I(n159), .Z(n158) );
  BUFFD0 U158 ( .I(n160), .Z(n159) );
  BUFFD0 U159 ( .I(n161), .Z(n160) );
  CKBXD0 U160 ( .I(DivideFactor[4]), .Z(n182) );
  BUFFD0 U161 ( .I(n162), .Z(n161) );
  BUFFD0 U162 ( .I(n163), .Z(n162) );
  BUFFD0 U163 ( .I(n164), .Z(n163) );
  BUFFD0 U164 ( .I(n165), .Z(n164) );
  BUFFD0 U165 ( .I(n166), .Z(n165) );
  BUFFD0 U166 ( .I(n167), .Z(n166) );
  BUFFD0 U167 ( .I(n168), .Z(n167) );
  BUFFD0 U168 ( .I(n169), .Z(n168) );
  BUFFD0 U169 ( .I(n170), .Z(n169) );
  BUFFD0 U170 ( .I(n171), .Z(n170) );
  BUFFD0 U171 ( .I(n172), .Z(n171) );
  BUFFD0 U172 ( .I(n173), .Z(n172) );
  BUFFD0 U173 ( .I(n174), .Z(n173) );
  BUFFD0 U174 ( .I(n175), .Z(n174) );
  BUFFD0 U175 ( .I(n176), .Z(n175) );
  BUFFD0 U176 ( .I(n177), .Z(n176) );
  BUFFD0 U177 ( .I(n178), .Z(n177) );
  BUFFD0 U178 ( .I(n179), .Z(n178) );
  BUFFD0 U179 ( .I(n180), .Z(n179) );
  BUFFD0 U180 ( .I(n181), .Z(n180) );
  BUFFD0 U181 ( .I(n126), .Z(n181) );
  BUFFD0 U182 ( .I(n186), .Z(n183) );
  BUFFD0 U183 ( .I(n443), .Z(n184) );
  BUFFD0 U184 ( .I(n184), .Z(n185) );
  BUFFD0 U185 ( .I(n187), .Z(n186) );
  BUFFD0 U186 ( .I(n188), .Z(n187) );
  BUFFD0 U187 ( .I(n189), .Z(n188) );
  BUFFD0 U188 ( .I(n190), .Z(n189) );
  BUFFD0 U189 ( .I(n191), .Z(n190) );
  BUFFD0 U190 ( .I(n192), .Z(n191) );
  BUFFD0 U191 ( .I(n193), .Z(n192) );
  BUFFD0 U192 ( .I(n194), .Z(n193) );
  BUFFD0 U193 ( .I(n195), .Z(n194) );
  BUFFD0 U194 ( .I(n196), .Z(n195) );
  BUFFD0 U195 ( .I(n197), .Z(n196) );
  BUFFD0 U196 ( .I(n198), .Z(n197) );
  BUFFD0 U197 ( .I(n199), .Z(n198) );
  BUFFD0 U198 ( .I(n200), .Z(n199) );
  BUFFD0 U199 ( .I(n201), .Z(n200) );
  BUFFD0 U200 ( .I(n202), .Z(n201) );
  BUFFD0 U201 ( .I(n203), .Z(n202) );
  BUFFD0 U202 ( .I(n204), .Z(n203) );
  BUFFD0 U203 ( .I(n205), .Z(n204) );
  BUFFD0 U204 ( .I(n206), .Z(n205) );
  BUFFD0 U205 ( .I(n207), .Z(n206) );
  BUFFD0 U206 ( .I(n208), .Z(n207) );
  BUFFD0 U207 ( .I(n209), .Z(n208) );
  BUFFD0 U208 ( .I(n210), .Z(n209) );
  BUFFD0 U209 ( .I(n211), .Z(n210) );
  BUFFD0 U210 ( .I(n212), .Z(n211) );
  BUFFD0 U211 ( .I(n213), .Z(n212) );
  BUFFD0 U212 ( .I(n214), .Z(n213) );
  BUFFD0 U213 ( .I(n215), .Z(n214) );
  BUFFD0 U214 ( .I(n216), .Z(n215) );
  BUFFD0 U215 ( .I(n217), .Z(n216) );
  BUFFD0 U216 ( .I(n218), .Z(n217) );
  BUFFD0 U217 ( .I(n219), .Z(n218) );
  BUFFD0 U218 ( .I(n220), .Z(n219) );
  BUFFD0 U219 ( .I(n221), .Z(n220) );
  BUFFD0 U220 ( .I(n222), .Z(n221) );
  BUFFD0 U221 ( .I(n223), .Z(n222) );
  BUFFD0 U222 ( .I(n224), .Z(n223) );
  BUFFD0 U223 ( .I(n225), .Z(n224) );
  BUFFD0 U224 ( .I(n226), .Z(n225) );
  BUFFD0 U225 ( .I(n227), .Z(n226) );
  BUFFD0 U226 ( .I(n228), .Z(n227) );
  BUFFD0 U227 ( .I(n229), .Z(n228) );
  BUFFD0 U228 ( .I(n230), .Z(n229) );
  BUFFD0 U229 ( .I(n231), .Z(n230) );
  BUFFD0 U230 ( .I(n232), .Z(n231) );
  BUFFD0 U231 ( .I(n233), .Z(n232) );
  BUFFD0 U232 ( .I(n234), .Z(n233) );
  BUFFD0 U233 ( .I(n235), .Z(n234) );
  BUFFD0 U234 ( .I(n236), .Z(n235) );
  BUFFD0 U235 ( .I(n237), .Z(n236) );
  BUFFD0 U236 ( .I(n238), .Z(n237) );
  BUFFD0 U237 ( .I(n239), .Z(n238) );
  BUFFD0 U238 ( .I(n185), .Z(n239) );
  BUFFD0 U239 ( .I(n241), .Z(n240) );
  BUFFD0 U240 ( .I(DivideFactor[1]), .Z(n241) );
  BUFFD0 U241 ( .I(n245), .Z(n242) );
  BUFFD0 U242 ( .I(n441), .Z(n243) );
  BUFFD0 U243 ( .I(n243), .Z(n244) );
  BUFFD0 U244 ( .I(n246), .Z(n245) );
  BUFFD0 U245 ( .I(n247), .Z(n246) );
  BUFFD0 U246 ( .I(n248), .Z(n247) );
  BUFFD0 U247 ( .I(n249), .Z(n248) );
  BUFFD0 U248 ( .I(n250), .Z(n249) );
  BUFFD0 U249 ( .I(n251), .Z(n250) );
  BUFFD0 U250 ( .I(n252), .Z(n251) );
  BUFFD0 U251 ( .I(n253), .Z(n252) );
  BUFFD0 U252 ( .I(n254), .Z(n253) );
  BUFFD0 U253 ( .I(n255), .Z(n254) );
  BUFFD0 U254 ( .I(n256), .Z(n255) );
  BUFFD0 U255 ( .I(n257), .Z(n256) );
  BUFFD0 U256 ( .I(n258), .Z(n257) );
  BUFFD0 U257 ( .I(n259), .Z(n258) );
  BUFFD0 U258 ( .I(n260), .Z(n259) );
  BUFFD0 U259 ( .I(n261), .Z(n260) );
  BUFFD0 U260 ( .I(n262), .Z(n261) );
  BUFFD0 U261 ( .I(n263), .Z(n262) );
  BUFFD0 U262 ( .I(n264), .Z(n263) );
  BUFFD0 U263 ( .I(n265), .Z(n264) );
  BUFFD0 U264 ( .I(n266), .Z(n265) );
  BUFFD0 U265 ( .I(n267), .Z(n266) );
  BUFFD0 U266 ( .I(n268), .Z(n267) );
  BUFFD0 U267 ( .I(n269), .Z(n268) );
  BUFFD0 U268 ( .I(n270), .Z(n269) );
  BUFFD0 U269 ( .I(n271), .Z(n270) );
  BUFFD0 U270 ( .I(n272), .Z(n271) );
  BUFFD0 U271 ( .I(n273), .Z(n272) );
  BUFFD0 U272 ( .I(n274), .Z(n273) );
  BUFFD0 U273 ( .I(n275), .Z(n274) );
  BUFFD0 U274 ( .I(n276), .Z(n275) );
  BUFFD0 U275 ( .I(n277), .Z(n276) );
  BUFFD0 U276 ( .I(n278), .Z(n277) );
  BUFFD0 U277 ( .I(n279), .Z(n278) );
  BUFFD0 U278 ( .I(n280), .Z(n279) );
  BUFFD0 U279 ( .I(n281), .Z(n280) );
  BUFFD0 U280 ( .I(n282), .Z(n281) );
  BUFFD0 U281 ( .I(n283), .Z(n282) );
  BUFFD0 U282 ( .I(n284), .Z(n283) );
  BUFFD0 U283 ( .I(n285), .Z(n284) );
  BUFFD0 U284 ( .I(n286), .Z(n285) );
  BUFFD0 U285 ( .I(n287), .Z(n286) );
  BUFFD0 U286 ( .I(n288), .Z(n287) );
  BUFFD0 U287 ( .I(n289), .Z(n288) );
  BUFFD0 U288 ( .I(n290), .Z(n289) );
  BUFFD0 U289 ( .I(n291), .Z(n290) );
  BUFFD0 U290 ( .I(n292), .Z(n291) );
  BUFFD0 U291 ( .I(n293), .Z(n292) );
  BUFFD0 U292 ( .I(n294), .Z(n293) );
  BUFFD0 U293 ( .I(n295), .Z(n294) );
  BUFFD0 U294 ( .I(n296), .Z(n295) );
  BUFFD0 U295 ( .I(n297), .Z(n296) );
  BUFFD0 U296 ( .I(n298), .Z(n297) );
  BUFFD0 U297 ( .I(n244), .Z(n298) );
  BUFFD0 U298 ( .I(DivideFactor[0]), .Z(n299) );
  CKBXD0 U299 ( .I(n299), .Z(n300) );
  BUFFD0 U300 ( .I(n305), .Z(n301) );
  BUFFD0 U301 ( .I(N51), .Z(n302) );
  BUFFD0 U302 ( .I(n302), .Z(n303) );
  BUFFD0 U303 ( .I(n303), .Z(n304) );
  BUFFD0 U304 ( .I(n306), .Z(n305) );
  BUFFD0 U305 ( .I(n307), .Z(n306) );
  BUFFD0 U306 ( .I(n308), .Z(n307) );
  BUFFD0 U307 ( .I(n309), .Z(n308) );
  BUFFD0 U308 ( .I(n310), .Z(n309) );
  BUFFD0 U309 ( .I(n311), .Z(n310) );
  BUFFD0 U310 ( .I(n312), .Z(n311) );
  BUFFD0 U311 ( .I(n313), .Z(n312) );
  BUFFD0 U312 ( .I(n314), .Z(n313) );
  BUFFD0 U313 ( .I(n315), .Z(n314) );
  BUFFD0 U314 ( .I(n316), .Z(n315) );
  BUFFD0 U315 ( .I(n317), .Z(n316) );
  BUFFD0 U316 ( .I(n318), .Z(n317) );
  BUFFD0 U317 ( .I(n319), .Z(n318) );
  BUFFD0 U318 ( .I(n320), .Z(n319) );
  BUFFD0 U319 ( .I(n321), .Z(n320) );
  BUFFD0 U320 ( .I(n322), .Z(n321) );
  BUFFD0 U321 ( .I(n323), .Z(n322) );
  BUFFD0 U322 ( .I(n324), .Z(n323) );
  BUFFD0 U323 ( .I(n325), .Z(n324) );
  BUFFD0 U324 ( .I(n326), .Z(n325) );
  BUFFD0 U325 ( .I(n327), .Z(n326) );
  BUFFD0 U326 ( .I(n328), .Z(n327) );
  BUFFD0 U327 ( .I(n329), .Z(n328) );
  BUFFD0 U328 ( .I(n330), .Z(n329) );
  BUFFD0 U329 ( .I(n331), .Z(n330) );
  BUFFD0 U330 ( .I(n332), .Z(n331) );
  BUFFD0 U331 ( .I(n333), .Z(n332) );
  BUFFD0 U332 ( .I(n334), .Z(n333) );
  BUFFD0 U333 ( .I(n335), .Z(n334) );
  BUFFD0 U334 ( .I(n336), .Z(n335) );
  BUFFD0 U335 ( .I(n337), .Z(n336) );
  BUFFD0 U336 ( .I(n338), .Z(n337) );
  BUFFD0 U337 ( .I(n339), .Z(n338) );
  BUFFD0 U338 ( .I(n340), .Z(n339) );
  BUFFD0 U339 ( .I(n341), .Z(n340) );
  BUFFD0 U340 ( .I(n342), .Z(n341) );
  BUFFD0 U341 ( .I(n343), .Z(n342) );
  BUFFD0 U342 ( .I(n344), .Z(n343) );
  BUFFD0 U343 ( .I(n345), .Z(n344) );
  BUFFD0 U344 ( .I(n346), .Z(n345) );
  BUFFD0 U345 ( .I(n347), .Z(n346) );
  BUFFD0 U346 ( .I(n348), .Z(n347) );
  BUFFD0 U347 ( .I(n349), .Z(n348) );
  BUFFD0 U348 ( .I(n350), .Z(n349) );
  BUFFD0 U349 ( .I(n351), .Z(n350) );
  BUFFD0 U350 ( .I(n352), .Z(n351) );
  BUFFD0 U351 ( .I(n353), .Z(n352) );
  BUFFD0 U352 ( .I(n354), .Z(n353) );
  BUFFD0 U353 ( .I(n355), .Z(n354) );
  BUFFD0 U354 ( .I(n356), .Z(n355) );
  BUFFD0 U355 ( .I(n357), .Z(n356) );
  BUFFD0 U356 ( .I(n358), .Z(n357) );
  BUFFD0 U357 ( .I(n359), .Z(n358) );
  BUFFD0 U358 ( .I(n304), .Z(n359) );
  BUFFD0 U359 ( .I(n362), .Z(n360) );
  BUFFD0 U360 ( .I(n360), .Z(n361) );
  BUFFD0 U361 ( .I(n363), .Z(n362) );
  BUFFD0 U362 ( .I(n364), .Z(n363) );
  BUFFD0 U363 ( .I(n365), .Z(n364) );
  BUFFD0 U364 ( .I(n366), .Z(n365) );
  BUFFD0 U365 ( .I(n367), .Z(n366) );
  BUFFD0 U366 ( .I(n368), .Z(n367) );
  BUFFD0 U367 ( .I(n369), .Z(n368) );
  BUFFD0 U368 ( .I(n370), .Z(n369) );
  BUFFD0 U369 ( .I(n371), .Z(n370) );
  BUFFD0 U370 ( .I(n372), .Z(n371) );
  BUFFD0 U371 ( .I(n373), .Z(n372) );
  BUFFD0 U372 ( .I(n374), .Z(n373) );
  BUFFD0 U373 ( .I(n375), .Z(n374) );
  BUFFD0 U374 ( .I(n376), .Z(n375) );
  BUFFD0 U375 ( .I(n377), .Z(n376) );
  BUFFD0 U376 ( .I(n378), .Z(n377) );
  BUFFD0 U377 ( .I(n379), .Z(n378) );
  BUFFD0 U378 ( .I(n380), .Z(n379) );
  BUFFD0 U379 ( .I(n381), .Z(n380) );
  BUFFD0 U380 ( .I(n382), .Z(n381) );
  BUFFD0 U381 ( .I(n383), .Z(n382) );
  BUFFD0 U382 ( .I(n384), .Z(n383) );
  BUFFD0 U383 ( .I(n385), .Z(n384) );
  BUFFD0 U384 ( .I(n386), .Z(n385) );
  BUFFD0 U385 ( .I(n387), .Z(n386) );
  BUFFD0 U386 ( .I(n388), .Z(n387) );
  BUFFD0 U387 ( .I(n389), .Z(n388) );
  BUFFD0 U388 ( .I(n390), .Z(n389) );
  BUFFD0 U389 ( .I(n391), .Z(n390) );
  BUFFD0 U390 ( .I(n392), .Z(n391) );
  BUFFD0 U391 ( .I(n393), .Z(n392) );
  BUFFD0 U392 ( .I(n394), .Z(n393) );
  BUFFD0 U393 ( .I(n395), .Z(n394) );
  BUFFD0 U394 ( .I(n396), .Z(n395) );
  BUFFD0 U395 ( .I(n397), .Z(n396) );
  BUFFD0 U396 ( .I(n398), .Z(n397) );
  BUFFD0 U397 ( .I(n399), .Z(n398) );
  BUFFD0 U398 ( .I(n400), .Z(n399) );
  BUFFD0 U399 ( .I(n401), .Z(n400) );
  BUFFD0 U400 ( .I(n402), .Z(n401) );
  BUFFD0 U401 ( .I(n403), .Z(n402) );
  BUFFD0 U402 ( .I(n404), .Z(n403) );
  BUFFD0 U403 ( .I(n405), .Z(n404) );
  BUFFD0 U404 ( .I(n406), .Z(n405) );
  BUFFD0 U405 ( .I(n407), .Z(n406) );
  BUFFD0 U406 ( .I(n408), .Z(n407) );
  BUFFD0 U407 ( .I(n409), .Z(n408) );
  BUFFD0 U408 ( .I(n410), .Z(n409) );
  BUFFD0 U409 ( .I(n411), .Z(n410) );
  BUFFD0 U410 ( .I(n412), .Z(n411) );
  BUFFD0 U411 ( .I(n413), .Z(n412) );
  BUFFD0 U412 ( .I(n414), .Z(n413) );
  BUFFD0 U413 ( .I(N54), .Z(n414) );
  BUFFD0 U414 ( .I(n426), .Z(n415) );
  INVD1 U415 ( .I(Reset), .ZN(n416) );
  AO222D0 U416 ( .A1(N27), .A2(n417), .B1(N35), .B2(n418), .C1(n300), .C2(n419), .Z(n441) );
  AO222D0 U417 ( .A1(N31), .A2(n417), .B1(N39), .B2(n418), .C1(n182), .C2(n419), .Z(n442) );
  AO222D0 U418 ( .A1(N28), .A2(n417), .B1(N36), .B2(n418), .C1(n240), .C2(n419), .Z(n443) );
  CKND0 U419 ( .CLK(n360), .CN(n419) );
  AN2D0 U420 ( .A1(n420), .A2(n421), .Z(n418) );
  AN3D0 U421 ( .A1(n422), .A2(n423), .A3(n424), .Z(n417) );
  CKXOR2D0 U422 ( .A1(ClockOut), .A2(n425), .Z(n444) );
  AO22D0 U423 ( .A1(N32), .A2(n424), .B1(N40), .B2(n420), .Z(N55) );
  CKND2D0 U424 ( .A1(AdjustFreq[1]), .A2(n421), .ZN(n427) );
  ND3D0 U425 ( .A1(n428), .A2(n423), .A3(n429), .ZN(n421) );
  ND4D0 U426 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(n240), .A4(n300), .ZN(n429) );
  IND3D0 U427 ( .A1(AdjustFreq[1]), .B1(n423), .B2(n422), .ZN(n426) );
  CKND2D0 U428 ( .A1(n182), .A2(DivideFactor[3]), .ZN(n422) );
  AO22D0 U429 ( .A1(N30), .A2(n424), .B1(N38), .B2(n420), .Z(N51) );
  AO22D0 U430 ( .A1(N29), .A2(n424), .B1(N37), .B2(n420), .Z(N49) );
  AN2D0 U431 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n420) );
  NR2D0 U432 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n424) );
  INR2D0 U433 ( .A1(N14), .B1(n425), .ZN(N21) );
  INR2D0 U434 ( .A1(N13), .B1(n425), .ZN(N20) );
  INR2D0 U435 ( .A1(N12), .B1(n425), .ZN(N19) );
  INR2D0 U436 ( .A1(N11), .B1(n425), .ZN(N18) );
  INR2D0 U437 ( .A1(N10), .B1(n425), .ZN(N17) );
  INR2D0 U438 ( .A1(N9), .B1(n425), .ZN(N16) );
  OA21D0 U439 ( .A1(FastDivvy[5]), .A2(n423), .B(n430), .Z(n425) );
  IOA22D0 U440 ( .B1(n431), .B2(n432), .A1(n423), .A2(FastDivvy[5]), .ZN(n430)
         );
  AOI221D0 U441 ( .A1(FastDivvy[4]), .A2(n428), .B1(FastDivvy[3]), .B2(n433), 
        .C(n434), .ZN(n432) );
  AOI221D0 U442 ( .A1(DivideFactor[3]), .A2(n435), .B1(DivideFactor[2]), .B2(
        n436), .C(n437), .ZN(n434) );
  IAO21D0 U443 ( .A1(n436), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n437)
         );
  OAI32D0 U444 ( .A1(n438), .A2(FastDivvy[0]), .A3(n439), .B1(FastDivvy[1]), 
        .B2(n440), .ZN(n436) );
  AN2D0 U445 ( .A1(FastDivvy[1]), .A2(n440), .Z(n439) );
  CKND0 U446 ( .CLK(FastDivvy[3]), .CN(n435) );
  NR2D0 U447 ( .A1(FastDivvy[4]), .A2(n428), .ZN(n431) );
  CKND0 U448 ( .CLK(DivideFactor[5]), .CN(n423) );
  CKND0 U449 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U450 ( .A1(WireD[5]), .A2(n416), .ZN(WireD[0]) );
endmodule


module VFO_3 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_3_DW01_dec_0 \Sampler/sub_193  ( .A({n103, n168, n36, n69, n201, n237}), 
        .SUM({N40, N39, N38, N37, N36, N35}) );
  VFO_3_DW01_inc_0 \Sampler/add_190  ( .A({n103, n168, n36, n69, n201, n237}), 
        .SUM({N32, N31, N30, N29, N28, N27}) );
  VFO_3_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n239), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n239), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n239), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n239), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n239), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n239), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n267), .CP(FastClock), .CDN(n239), .Q(ClockOut)
         );
  EDFCND1 \DivideFactor_reg[3]  ( .D(n1), .E(n106), .CP(Sample), .CDN(n239), 
        .Q(DivideFactor[3]), .QN(n256) );
  EDFCND1 \DivideFactor_reg[2]  ( .D(n37), .E(n106), .CP(Sample), .CDN(n239), 
        .Q(DivideFactor[2]) );
  EDFCND1 \DivideFactor_reg[5]  ( .D(n70), .E(n106), .CP(Sample), .CDN(n239), 
        .Q(DivideFactor[5]), .QN(n246) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n135), .CP(Sample), .SDN(n239), .Q(
        DivideFactor[4]), .QN(n251) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n169), .CP(Sample), .SDN(n239), .Q(
        DivideFactor[1]), .QN(n263) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n203), .CP(Sample), .SDN(n239), .Q(
        DivideFactor[0]), .QN(n261) );
  CKBD0 U3 ( .CLK(n136), .C(n135) );
  BUFFD0 U4 ( .I(n3), .Z(n1) );
  BUFFD0 U5 ( .I(N51), .Z(n2) );
  BUFFD0 U6 ( .I(n4), .Z(n3) );
  BUFFD0 U7 ( .I(n5), .Z(n4) );
  BUFFD0 U8 ( .I(n6), .Z(n5) );
  BUFFD0 U9 ( .I(n7), .Z(n6) );
  BUFFD0 U10 ( .I(n8), .Z(n7) );
  BUFFD0 U11 ( .I(n9), .Z(n8) );
  BUFFD0 U12 ( .I(n10), .Z(n9) );
  BUFFD0 U13 ( .I(n11), .Z(n10) );
  BUFFD0 U14 ( .I(n12), .Z(n11) );
  BUFFD0 U15 ( .I(n13), .Z(n12) );
  BUFFD0 U16 ( .I(n14), .Z(n13) );
  BUFFD0 U17 ( .I(n15), .Z(n14) );
  BUFFD0 U18 ( .I(n16), .Z(n15) );
  BUFFD0 U19 ( .I(n20), .Z(n16) );
  BUFFD0 U20 ( .I(n22), .Z(n20) );
  BUFFD0 U21 ( .I(n23), .Z(n22) );
  BUFFD0 U22 ( .I(n24), .Z(n23) );
  BUFFD0 U23 ( .I(n25), .Z(n24) );
  BUFFD0 U24 ( .I(n26), .Z(n25) );
  BUFFD0 U25 ( .I(n27), .Z(n26) );
  BUFFD0 U26 ( .I(n28), .Z(n27) );
  BUFFD0 U27 ( .I(n29), .Z(n28) );
  BUFFD0 U28 ( .I(n30), .Z(n29) );
  BUFFD0 U29 ( .I(n31), .Z(n30) );
  BUFFD0 U30 ( .I(n32), .Z(n31) );
  BUFFD0 U31 ( .I(n33), .Z(n32) );
  BUFFD0 U32 ( .I(n34), .Z(n33) );
  BUFFD0 U33 ( .I(n35), .Z(n34) );
  BUFFD0 U34 ( .I(n2), .Z(n35) );
  BUFFD0 U35 ( .I(n142), .Z(n36) );
  CKBD0 U36 ( .CLK(DivideFactor[3]), .C(n142) );
  BUFFD0 U37 ( .I(n39), .Z(n37) );
  BUFFD0 U38 ( .I(N49), .Z(n38) );
  BUFFD0 U39 ( .I(n40), .Z(n39) );
  BUFFD0 U40 ( .I(n41), .Z(n40) );
  BUFFD0 U41 ( .I(n42), .Z(n41) );
  BUFFD0 U42 ( .I(n43), .Z(n42) );
  BUFFD0 U43 ( .I(n44), .Z(n43) );
  BUFFD0 U44 ( .I(n45), .Z(n44) );
  BUFFD0 U45 ( .I(n46), .Z(n45) );
  BUFFD0 U46 ( .I(n47), .Z(n46) );
  BUFFD0 U47 ( .I(n48), .Z(n47) );
  BUFFD0 U48 ( .I(n49), .Z(n48) );
  BUFFD0 U49 ( .I(n50), .Z(n49) );
  BUFFD0 U50 ( .I(n51), .Z(n50) );
  BUFFD0 U51 ( .I(n52), .Z(n51) );
  BUFFD0 U52 ( .I(n53), .Z(n52) );
  BUFFD0 U53 ( .I(n54), .Z(n53) );
  BUFFD0 U54 ( .I(n55), .Z(n54) );
  BUFFD0 U55 ( .I(n56), .Z(n55) );
  BUFFD0 U56 ( .I(n57), .Z(n56) );
  BUFFD0 U57 ( .I(n58), .Z(n57) );
  BUFFD0 U58 ( .I(n59), .Z(n58) );
  BUFFD0 U59 ( .I(n60), .Z(n59) );
  BUFFD0 U60 ( .I(n61), .Z(n60) );
  BUFFD0 U61 ( .I(n62), .Z(n61) );
  BUFFD0 U62 ( .I(n63), .Z(n62) );
  BUFFD0 U63 ( .I(n64), .Z(n63) );
  BUFFD0 U64 ( .I(n65), .Z(n64) );
  BUFFD0 U65 ( .I(n66), .Z(n65) );
  BUFFD0 U66 ( .I(n67), .Z(n66) );
  BUFFD0 U67 ( .I(n38), .Z(n67) );
  BUFFD0 U68 ( .I(DivideFactor[2]), .Z(n68) );
  CKBD0 U69 ( .CLK(n68), .C(n69) );
  BUFFD0 U70 ( .I(n72), .Z(n70) );
  BUFFD0 U71 ( .I(N55), .Z(n71) );
  BUFFD0 U72 ( .I(n73), .Z(n72) );
  BUFFD0 U73 ( .I(n74), .Z(n73) );
  BUFFD0 U74 ( .I(n75), .Z(n74) );
  BUFFD0 U75 ( .I(n76), .Z(n75) );
  BUFFD0 U76 ( .I(n77), .Z(n76) );
  BUFFD0 U77 ( .I(n78), .Z(n77) );
  BUFFD0 U78 ( .I(n79), .Z(n78) );
  BUFFD0 U79 ( .I(n80), .Z(n79) );
  BUFFD0 U80 ( .I(n81), .Z(n80) );
  BUFFD0 U81 ( .I(n82), .Z(n81) );
  BUFFD0 U82 ( .I(n83), .Z(n82) );
  BUFFD0 U83 ( .I(n84), .Z(n83) );
  BUFFD0 U84 ( .I(n85), .Z(n84) );
  BUFFD0 U85 ( .I(n86), .Z(n85) );
  BUFFD0 U86 ( .I(n87), .Z(n86) );
  BUFFD0 U87 ( .I(n88), .Z(n87) );
  BUFFD0 U88 ( .I(n89), .Z(n88) );
  BUFFD0 U89 ( .I(n90), .Z(n89) );
  BUFFD0 U90 ( .I(n91), .Z(n90) );
  BUFFD0 U91 ( .I(n92), .Z(n91) );
  BUFFD0 U92 ( .I(n93), .Z(n92) );
  BUFFD0 U93 ( .I(n94), .Z(n93) );
  BUFFD0 U94 ( .I(n95), .Z(n94) );
  BUFFD0 U95 ( .I(n96), .Z(n95) );
  BUFFD0 U96 ( .I(n97), .Z(n96) );
  BUFFD0 U97 ( .I(n98), .Z(n97) );
  BUFFD0 U98 ( .I(n99), .Z(n98) );
  BUFFD0 U99 ( .I(n100), .Z(n99) );
  BUFFD0 U100 ( .I(n71), .Z(n100) );
  BUFFD0 U101 ( .I(DivideFactor[5]), .Z(n101) );
  BUFFD0 U102 ( .I(n101), .Z(n102) );
  CKBD0 U103 ( .CLK(n102), .C(n103) );
  ND2D1P5 U104 ( .A1(AdjustFreq[1]), .A2(n244), .ZN(n250) );
  BUFFD0 U105 ( .I(N54), .Z(n104) );
  BUFFD0 U106 ( .I(n104), .Z(n105) );
  BUFFD0 U107 ( .I(n107), .Z(n106) );
  BUFFD0 U108 ( .I(n108), .Z(n107) );
  BUFFD0 U109 ( .I(n109), .Z(n108) );
  BUFFD0 U110 ( .I(n110), .Z(n109) );
  BUFFD0 U111 ( .I(n111), .Z(n110) );
  BUFFD0 U112 ( .I(n112), .Z(n111) );
  BUFFD0 U113 ( .I(n113), .Z(n112) );
  BUFFD0 U114 ( .I(n114), .Z(n113) );
  BUFFD0 U115 ( .I(n115), .Z(n114) );
  BUFFD0 U116 ( .I(n116), .Z(n115) );
  BUFFD0 U117 ( .I(n117), .Z(n116) );
  BUFFD0 U118 ( .I(n118), .Z(n117) );
  BUFFD0 U119 ( .I(n119), .Z(n118) );
  BUFFD0 U120 ( .I(n120), .Z(n119) );
  BUFFD0 U121 ( .I(n121), .Z(n120) );
  BUFFD0 U122 ( .I(n122), .Z(n121) );
  BUFFD0 U123 ( .I(n123), .Z(n122) );
  BUFFD0 U124 ( .I(n124), .Z(n123) );
  BUFFD0 U125 ( .I(n125), .Z(n124) );
  BUFFD0 U126 ( .I(n126), .Z(n125) );
  BUFFD0 U127 ( .I(n127), .Z(n126) );
  BUFFD0 U128 ( .I(n128), .Z(n127) );
  BUFFD0 U129 ( .I(n129), .Z(n128) );
  BUFFD0 U130 ( .I(n130), .Z(n129) );
  BUFFD0 U131 ( .I(n131), .Z(n130) );
  BUFFD0 U132 ( .I(n132), .Z(n131) );
  BUFFD0 U133 ( .I(n133), .Z(n132) );
  BUFFD0 U134 ( .I(n134), .Z(n133) );
  BUFFD0 U135 ( .I(n105), .Z(n134) );
  BUFFD0 U136 ( .I(n137), .Z(n136) );
  BUFFD0 U137 ( .I(n138), .Z(n137) );
  BUFFD0 U138 ( .I(n139), .Z(n138) );
  BUFFD0 U139 ( .I(n140), .Z(n139) );
  BUFFD0 U140 ( .I(n143), .Z(n140) );
  BUFFD0 U141 ( .I(DivideFactor[4]), .Z(n141) );
  BUFFD0 U142 ( .I(n144), .Z(n143) );
  BUFFD0 U143 ( .I(n145), .Z(n144) );
  BUFFD0 U144 ( .I(n146), .Z(n145) );
  BUFFD0 U145 ( .I(n147), .Z(n146) );
  CKBXD0 U146 ( .I(n141), .Z(n168) );
  BUFFD0 U147 ( .I(n148), .Z(n147) );
  BUFFD0 U148 ( .I(n149), .Z(n148) );
  BUFFD0 U149 ( .I(n150), .Z(n149) );
  BUFFD0 U150 ( .I(n151), .Z(n150) );
  BUFFD0 U151 ( .I(n152), .Z(n151) );
  BUFFD0 U152 ( .I(n153), .Z(n152) );
  BUFFD0 U153 ( .I(n154), .Z(n153) );
  BUFFD0 U154 ( .I(n155), .Z(n154) );
  BUFFD0 U155 ( .I(n156), .Z(n155) );
  BUFFD0 U156 ( .I(n157), .Z(n156) );
  BUFFD0 U157 ( .I(n158), .Z(n157) );
  BUFFD0 U158 ( .I(n159), .Z(n158) );
  BUFFD0 U159 ( .I(n160), .Z(n159) );
  BUFFD0 U160 ( .I(n161), .Z(n160) );
  BUFFD0 U161 ( .I(n162), .Z(n161) );
  BUFFD0 U162 ( .I(n163), .Z(n162) );
  BUFFD0 U163 ( .I(n164), .Z(n163) );
  BUFFD0 U164 ( .I(n165), .Z(n164) );
  BUFFD0 U165 ( .I(n166), .Z(n165) );
  BUFFD0 U166 ( .I(n167), .Z(n166) );
  BUFFD0 U167 ( .I(n265), .Z(n167) );
  BUFFD0 U168 ( .I(n170), .Z(n169) );
  BUFFD0 U169 ( .I(n171), .Z(n170) );
  BUFFD0 U170 ( .I(n172), .Z(n171) );
  BUFFD0 U171 ( .I(n173), .Z(n172) );
  BUFFD0 U172 ( .I(n174), .Z(n173) );
  BUFFD0 U173 ( .I(n175), .Z(n174) );
  BUFFD0 U174 ( .I(n176), .Z(n175) );
  BUFFD0 U175 ( .I(n177), .Z(n176) );
  BUFFD0 U176 ( .I(n178), .Z(n177) );
  BUFFD0 U177 ( .I(n179), .Z(n178) );
  BUFFD0 U178 ( .I(n180), .Z(n179) );
  BUFFD0 U179 ( .I(n181), .Z(n180) );
  BUFFD0 U180 ( .I(n182), .Z(n181) );
  BUFFD0 U181 ( .I(n183), .Z(n182) );
  BUFFD0 U182 ( .I(n184), .Z(n183) );
  BUFFD0 U183 ( .I(n185), .Z(n184) );
  BUFFD0 U184 ( .I(n186), .Z(n185) );
  BUFFD0 U185 ( .I(n187), .Z(n186) );
  BUFFD0 U186 ( .I(n188), .Z(n187) );
  BUFFD0 U187 ( .I(n189), .Z(n188) );
  BUFFD0 U188 ( .I(n190), .Z(n189) );
  BUFFD0 U189 ( .I(n191), .Z(n190) );
  BUFFD0 U190 ( .I(n192), .Z(n191) );
  BUFFD0 U191 ( .I(n193), .Z(n192) );
  BUFFD0 U192 ( .I(n194), .Z(n193) );
  BUFFD0 U193 ( .I(n195), .Z(n194) );
  BUFFD0 U194 ( .I(n196), .Z(n195) );
  BUFFD0 U195 ( .I(n197), .Z(n196) );
  BUFFD0 U196 ( .I(n198), .Z(n197) );
  BUFFD0 U197 ( .I(n199), .Z(n198) );
  BUFFD0 U198 ( .I(n200), .Z(n199) );
  BUFFD0 U199 ( .I(n266), .Z(n200) );
  BUFFD0 U200 ( .I(n202), .Z(n201) );
  BUFFD0 U201 ( .I(DivideFactor[1]), .Z(n202) );
  BUFFD0 U202 ( .I(n204), .Z(n203) );
  BUFFD0 U203 ( .I(n205), .Z(n204) );
  BUFFD0 U204 ( .I(n206), .Z(n205) );
  BUFFD0 U205 ( .I(n207), .Z(n206) );
  BUFFD0 U206 ( .I(n208), .Z(n207) );
  BUFFD0 U207 ( .I(n209), .Z(n208) );
  BUFFD0 U208 ( .I(n210), .Z(n209) );
  BUFFD0 U209 ( .I(n211), .Z(n210) );
  BUFFD0 U210 ( .I(n212), .Z(n211) );
  BUFFD0 U211 ( .I(n213), .Z(n212) );
  BUFFD0 U212 ( .I(n214), .Z(n213) );
  BUFFD0 U213 ( .I(n215), .Z(n214) );
  BUFFD0 U214 ( .I(n216), .Z(n215) );
  BUFFD0 U215 ( .I(n217), .Z(n216) );
  BUFFD0 U216 ( .I(n218), .Z(n217) );
  BUFFD0 U217 ( .I(n219), .Z(n218) );
  BUFFD0 U218 ( .I(n220), .Z(n219) );
  BUFFD0 U219 ( .I(n221), .Z(n220) );
  BUFFD0 U220 ( .I(n222), .Z(n221) );
  BUFFD0 U221 ( .I(n224), .Z(n222) );
  CKBD0 U222 ( .CLK(n246), .C(n223) );
  BUFFD0 U223 ( .I(n225), .Z(n224) );
  BUFFD0 U224 ( .I(n226), .Z(n225) );
  BUFFD0 U225 ( .I(n227), .Z(n226) );
  BUFFD0 U226 ( .I(n228), .Z(n227) );
  BUFFD0 U227 ( .I(n229), .Z(n228) );
  BUFFD0 U228 ( .I(n230), .Z(n229) );
  BUFFD0 U229 ( .I(n231), .Z(n230) );
  BUFFD0 U230 ( .I(n232), .Z(n231) );
  BUFFD0 U231 ( .I(n233), .Z(n232) );
  BUFFD0 U232 ( .I(n234), .Z(n233) );
  BUFFD0 U233 ( .I(n235), .Z(n234) );
  BUFFD0 U234 ( .I(n264), .Z(n235) );
  BUFFD0 U235 ( .I(DivideFactor[0]), .Z(n236) );
  CKBXD0 U236 ( .I(n236), .Z(n237) );
  INVD1 U237 ( .I(Reset), .ZN(n239) );
  AO222D0 U238 ( .A1(N27), .A2(n240), .B1(N35), .B2(n241), .C1(n237), .C2(n242), .Z(n264) );
  AO222D0 U239 ( .A1(N31), .A2(n240), .B1(N39), .B2(n241), .C1(n168), .C2(n242), .Z(n265) );
  AO222D0 U240 ( .A1(N28), .A2(n240), .B1(N36), .B2(n241), .C1(n201), .C2(n242), .Z(n266) );
  CKND0 U241 ( .CLK(N54), .CN(n242) );
  AN2D0 U242 ( .A1(n243), .A2(n244), .Z(n241) );
  AN3D0 U243 ( .A1(n245), .A2(n223), .A3(n247), .Z(n240) );
  CKXOR2D0 U244 ( .A1(ClockOut), .A2(n248), .Z(n267) );
  AO22D0 U245 ( .A1(N32), .A2(n247), .B1(N40), .B2(n243), .Z(N55) );
  MUX2ND0 U246 ( .I0(n249), .I1(n250), .S(AdjustFreq[0]), .ZN(N54) );
  ND3D0 U247 ( .A1(n251), .A2(n223), .A3(n252), .ZN(n244) );
  ND4D0 U248 ( .A1(n142), .A2(DivideFactor[2]), .A3(n201), .A4(n237), .ZN(n252) );
  IND3D0 U249 ( .A1(AdjustFreq[1]), .B1(n223), .B2(n245), .ZN(n249) );
  CKND2D0 U250 ( .A1(n168), .A2(n142), .ZN(n245) );
  AO22D0 U251 ( .A1(N30), .A2(n247), .B1(N38), .B2(n243), .Z(N51) );
  AO22D0 U252 ( .A1(N29), .A2(n247), .B1(N37), .B2(n243), .Z(N49) );
  AN2D0 U253 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n243) );
  NR2D0 U254 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n247) );
  INR2D0 U255 ( .A1(N14), .B1(n248), .ZN(N21) );
  INR2D0 U256 ( .A1(N13), .B1(n248), .ZN(N20) );
  INR2D0 U257 ( .A1(N12), .B1(n248), .ZN(N19) );
  INR2D0 U258 ( .A1(N11), .B1(n248), .ZN(N18) );
  INR2D0 U259 ( .A1(N10), .B1(n248), .ZN(N17) );
  INR2D0 U260 ( .A1(N9), .B1(n248), .ZN(N16) );
  OA21D0 U261 ( .A1(FastDivvy[5]), .A2(n246), .B(n253), .Z(n248) );
  IOA22D0 U262 ( .B1(n254), .B2(n255), .A1(n246), .A2(FastDivvy[5]), .ZN(n253)
         );
  AOI221D0 U263 ( .A1(FastDivvy[4]), .A2(n251), .B1(FastDivvy[3]), .B2(n256), 
        .C(n257), .ZN(n255) );
  AOI221D0 U264 ( .A1(DivideFactor[3]), .A2(n258), .B1(DivideFactor[2]), .B2(
        n259), .C(n260), .ZN(n257) );
  IAO21D0 U265 ( .A1(n259), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n260)
         );
  OAI32D0 U266 ( .A1(n261), .A2(FastDivvy[0]), .A3(n262), .B1(FastDivvy[1]), 
        .B2(n263), .ZN(n259) );
  AN2D0 U267 ( .A1(FastDivvy[1]), .A2(n263), .Z(n262) );
  CKND0 U268 ( .CLK(FastDivvy[3]), .CN(n258) );
  NR2D0 U269 ( .A1(FastDivvy[4]), .A2(n251), .ZN(n254) );
  CKND0 U270 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U271 ( .A1(WireD[5]), .A2(n239), .ZN(WireD[0]) );
endmodule


module MultiCounter_1 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [3:0] Ctr;

  MultiCounter_1_DW01_inc_0 add_16 ( .A({CarryOut, n10, n5, n1, n6}), .SUM({N5, 
        N4, N3, N2, N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n11), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n11), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n11), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n11), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n11), .Q(CarryOut) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(Ctr[1]), .Z(n4) );
  BUFFD0 U7 ( .I(Ctr[2]), .Z(n5) );
  BUFFD0 U8 ( .I(n7), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(Ctr[0]), .Z(n9) );
  BUFFD0 U12 ( .I(Ctr[3]), .Z(n10) );
  INVD1 U13 ( .I(Reset), .ZN(n11) );
endmodule


module MultiCounter_2 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [3:0] Ctr;

  MultiCounter_2_DW01_inc_0 add_16 ( .A({CarryOut, n10, n5, n1, n6}), .SUM({N5, 
        N4, N3, N2, N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n11), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n11), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n11), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n11), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n11), .Q(CarryOut) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(Ctr[1]), .Z(n4) );
  BUFFD0 U7 ( .I(Ctr[2]), .Z(n5) );
  BUFFD0 U8 ( .I(n7), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(Ctr[0]), .Z(n9) );
  BUFFD0 U12 ( .I(Ctr[3]), .Z(n10) );
  INVD1 U13 ( .I(Reset), .ZN(n11) );
endmodule


module MultiCounter_3 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [3:0] Ctr;

  MultiCounter_3_DW01_inc_0 add_16 ( .A({CarryOut, n10, n5, n1, n6}), .SUM({N5, 
        N4, N3, N2, N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n11), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n11), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n11), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n11), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n11), .Q(CarryOut) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(Ctr[1]), .Z(n4) );
  BUFFD0 U7 ( .I(Ctr[2]), .Z(n5) );
  BUFFD0 U8 ( .I(n7), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(Ctr[0]), .Z(n9) );
  BUFFD0 U12 ( .I(Ctr[3]), .Z(n10) );
  INVD1 U13 ( .I(Reset), .ZN(n11) );
endmodule


module MultiCounter_1_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n15, n16, n17, n18, n19, \carry[4] , \carry[3] , \carry[2] , n3, n4,
         n5, n7, n8, n9, n12, n13, n14;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(n16) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(n18) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(n17) );
  BUFFD0 U1 ( .I(n18), .Z(SUM[1]) );
  BUFFD0 U2 ( .I(n3), .Z(SUM[2]) );
  BUFFD0 U3 ( .I(n4), .Z(n3) );
  BUFFD0 U4 ( .I(n5), .Z(n4) );
  BUFFD0 U5 ( .I(n17), .Z(n5) );
  BUFFD0 U6 ( .I(n7), .Z(SUM[3]) );
  BUFFD0 U7 ( .I(n8), .Z(n7) );
  BUFFD0 U8 ( .I(n9), .Z(n8) );
  BUFFD0 U9 ( .I(n16), .Z(n9) );
  BUFFD0 U10 ( .I(n19), .Z(SUM[0]) );
  BUFFD0 U11 ( .I(n12), .Z(SUM[4]) );
  BUFFD0 U12 ( .I(n13), .Z(n12) );
  BUFFD0 U13 ( .I(n14), .Z(n13) );
  BUFFD0 U14 ( .I(n15), .Z(n14) );
  XOR2D0 U15 ( .A1(\carry[4] ), .A2(A[4]), .Z(n15) );
  CKND0 U16 ( .CLK(A[0]), .CN(n19) );
endmodule


module VFO_1_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_1_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n2, \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D1 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(n2) );
  BUFFD0 U2 ( .I(n2), .Z(SUM[4]) );
  CKND0 U3 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_2_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n15, n16, n17, n18, n19, \carry[4] , \carry[3] , \carry[2] , n3, n4,
         n5, n7, n8, n9, n12, n13, n14;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(n16) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(n18) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(n17) );
  BUFFD0 U1 ( .I(n18), .Z(SUM[1]) );
  BUFFD0 U2 ( .I(n3), .Z(SUM[2]) );
  BUFFD0 U3 ( .I(n4), .Z(n3) );
  BUFFD0 U4 ( .I(n5), .Z(n4) );
  BUFFD0 U5 ( .I(n17), .Z(n5) );
  BUFFD0 U6 ( .I(n7), .Z(SUM[3]) );
  BUFFD0 U7 ( .I(n8), .Z(n7) );
  BUFFD0 U8 ( .I(n9), .Z(n8) );
  BUFFD0 U9 ( .I(n16), .Z(n9) );
  BUFFD0 U10 ( .I(n19), .Z(SUM[0]) );
  BUFFD0 U11 ( .I(n12), .Z(SUM[4]) );
  BUFFD0 U12 ( .I(n13), .Z(n12) );
  BUFFD0 U13 ( .I(n14), .Z(n13) );
  BUFFD0 U14 ( .I(n15), .Z(n14) );
  XOR2D0 U15 ( .A1(\carry[4] ), .A2(A[4]), .Z(n15) );
  CKND0 U16 ( .CLK(A[0]), .CN(n19) );
endmodule


module VFO_2_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  XOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module SerEncoder_DWid32_1_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n11, n12, n13, n14, n15, n6, n7, n8, n9, n10;

  BUFFD0 U1 ( .I(n11), .Z(SUM[5]) );
  XOR2D0 U2 ( .A1(A[5]), .A2(n6), .Z(n11) );
  BUFFD0 U3 ( .I(n12), .Z(SUM[4]) );
  BUFFD0 U4 ( .I(n13), .Z(SUM[2]) );
  BUFFD0 U5 ( .I(n14), .Z(SUM[1]) );
  BUFFD0 U6 ( .I(n15), .Z(SUM[0]) );
  NR2D0 U7 ( .A1(A[4]), .A2(n7), .ZN(n6) );
  XNR2D0 U8 ( .A1(n7), .A2(A[4]), .ZN(n12) );
  OAI21D0 U9 ( .A1(n8), .A2(n9), .B(n7), .ZN(SUM[3]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n7) );
  CKND0 U11 ( .CLK(A[3]), .CN(n9) );
  AO21D0 U12 ( .A1(n10), .A2(A[2]), .B(n8), .Z(n13) );
  NR2D0 U13 ( .A1(n10), .A2(A[2]), .ZN(n8) );
  IOA21D0 U14 ( .A1(A[0]), .A2(A[1]), .B(n10), .ZN(n14) );
  IND2D0 U15 ( .A1(A[1]), .B1(n15), .ZN(n10) );
  CKND0 U16 ( .CLK(A[0]), .CN(n15) );
endmodule


module MultiCounter_3_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n15, n16, n17, n18, n19, \carry[4] , \carry[3] , \carry[2] , n3, n4,
         n5, n7, n8, n9, n12, n13, n14;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(n16) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(n18) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(n17) );
  BUFFD0 U1 ( .I(n18), .Z(SUM[1]) );
  BUFFD0 U2 ( .I(n3), .Z(SUM[2]) );
  BUFFD0 U3 ( .I(n4), .Z(n3) );
  BUFFD0 U4 ( .I(n5), .Z(n4) );
  BUFFD0 U5 ( .I(n17), .Z(n5) );
  BUFFD0 U6 ( .I(n7), .Z(SUM[3]) );
  BUFFD0 U7 ( .I(n8), .Z(n7) );
  BUFFD0 U8 ( .I(n9), .Z(n8) );
  BUFFD0 U9 ( .I(n16), .Z(n9) );
  BUFFD0 U10 ( .I(n19), .Z(SUM[0]) );
  BUFFD0 U11 ( .I(n12), .Z(SUM[4]) );
  BUFFD0 U12 ( .I(n13), .Z(n12) );
  BUFFD0 U13 ( .I(n14), .Z(n13) );
  BUFFD0 U14 ( .I(n15), .Z(n14) );
  XOR2D0 U15 ( .A1(\carry[4] ), .A2(A[4]), .Z(n15) );
  CKND0 U16 ( .CLK(A[0]), .CN(n19) );
endmodule


module VFO_3_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_0_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n2, \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D1 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(n2) );
  BUFFD0 U2 ( .I(n2), .Z(SUM[4]) );
  CKND0 U3 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_0_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n15, n16, n17, n18, n19, \carry[4] , \carry[3] , \carry[2] , n3, n4,
         n5, n7, n8, n9, n12, n13, n14;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(n16) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(n18) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(n17) );
  BUFFD0 U1 ( .I(n18), .Z(SUM[1]) );
  BUFFD0 U2 ( .I(n3), .Z(SUM[2]) );
  BUFFD0 U3 ( .I(n4), .Z(n3) );
  BUFFD0 U4 ( .I(n5), .Z(n4) );
  BUFFD0 U5 ( .I(n17), .Z(n5) );
  BUFFD0 U6 ( .I(n7), .Z(SUM[3]) );
  BUFFD0 U7 ( .I(n8), .Z(n7) );
  BUFFD0 U8 ( .I(n9), .Z(n8) );
  BUFFD0 U9 ( .I(n16), .Z(n9) );
  BUFFD0 U10 ( .I(n19), .Z(SUM[0]) );
  BUFFD0 U11 ( .I(n12), .Z(SUM[4]) );
  BUFFD0 U12 ( .I(n13), .Z(n12) );
  BUFFD0 U13 ( .I(n14), .Z(n13) );
  BUFFD0 U14 ( .I(n15), .Z(n14) );
  XOR2D0 U15 ( .A1(\carry[4] ), .A2(A[4]), .Z(n15) );
  CKND0 U16 ( .CLK(A[0]), .CN(n19) );
endmodule


module VFO_0_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  XOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module SerEncoder_DWid32_0_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n11, n12, n13, n14, n15, n6, n7, n8, n9, n10;

  BUFFD0 U1 ( .I(n11), .Z(SUM[5]) );
  XOR2D0 U2 ( .A1(A[5]), .A2(n6), .Z(n11) );
  BUFFD0 U3 ( .I(n12), .Z(SUM[4]) );
  BUFFD0 U4 ( .I(n13), .Z(SUM[2]) );
  BUFFD0 U5 ( .I(n14), .Z(SUM[1]) );
  BUFFD0 U6 ( .I(n15), .Z(SUM[0]) );
  NR2D0 U7 ( .A1(A[4]), .A2(n7), .ZN(n6) );
  XNR2D0 U8 ( .A1(n7), .A2(A[4]), .ZN(n12) );
  OAI21D0 U9 ( .A1(n8), .A2(n9), .B(n7), .ZN(SUM[3]) );
  CKND2D0 U10 ( .A1(n8), .A2(n9), .ZN(n7) );
  CKND0 U11 ( .CLK(A[3]), .CN(n9) );
  AO21D0 U12 ( .A1(n10), .A2(A[2]), .B(n8), .Z(n13) );
  NR2D0 U13 ( .A1(n10), .A2(A[2]), .ZN(n8) );
  IOA21D0 U14 ( .A1(A[0]), .A2(A[1]), .B(n10), .ZN(n14) );
  IND2D0 U15 ( .A1(A[1]), .B1(n15), .ZN(n10) );
  CKND0 U16 ( .CLK(A[0]), .CN(n15) );
endmodule

